magic
tech scmos
timestamp 1714320391
<< metal1 >>
rect -1388 4104 -1332 4128
rect -481 4126 -419 4133
rect -1080 4094 -1032 4124
rect -779 4096 -728 4123
rect -483 4093 -419 4126
rect -170 4106 -134 4127
rect -483 4087 -421 4093
rect 117 4090 183 4115
rect 715 4096 772 4125
rect 721 4088 772 4096
rect 1022 4095 1083 4120
rect 1326 4098 1369 4128
rect 1628 4106 1665 4123
rect 1930 4095 1975 4122
rect 2219 4101 2278 4133
rect 2809 4089 2880 4127
rect 3109 4091 3177 4125
rect -1389 3381 -1385 3392
rect -1477 3377 -1385 3381
rect -1177 3365 -1173 3378
rect -1089 3365 -1085 3392
rect -1177 3361 -1085 3365
rect -876 3364 -872 3381
rect -789 3364 -785 3392
rect -576 3371 -572 3379
rect -489 3371 -485 3392
rect -576 3367 -485 3371
rect -276 3370 -272 3379
rect -189 3370 -185 3392
rect -276 3366 -185 3370
rect 24 3371 28 3379
rect 111 3371 115 3392
rect 24 3367 115 3371
rect 623 3369 627 3380
rect 711 3369 715 3392
rect 623 3365 715 3369
rect 923 3366 927 3380
rect 1011 3366 1015 3392
rect 1223 3371 1227 3381
rect 1311 3371 1315 3392
rect 1223 3367 1315 3371
rect -876 3360 -785 3364
rect 923 3362 1015 3366
rect 1523 3365 1527 3379
rect 1611 3365 1615 3392
rect 1823 3371 1827 3380
rect 1911 3371 1915 3392
rect 1823 3367 1915 3371
rect 2123 3371 2127 3380
rect 2211 3371 2215 3392
rect 2723 3376 2727 3379
rect 2811 3376 2815 3392
rect 2723 3372 2815 3376
rect 3023 3377 3027 3380
rect 3111 3377 3115 3392
rect 3023 3373 3115 3377
rect 2123 3367 2215 3371
rect 1523 3361 1615 3365
rect -2228 3222 -2189 3282
rect 3994 3231 4024 3269
rect -1492 3211 -1470 3215
rect -1474 3128 -1470 3211
rect -1481 3124 -1470 3128
rect 3267 3211 3292 3215
rect 3267 3127 3271 3211
rect 3267 3123 3280 3127
rect -2225 2927 -2191 2972
rect 4002 2931 4032 2966
rect -1492 2911 -1467 2915
rect -1471 2828 -1467 2911
rect -1480 2824 -1467 2828
rect -2227 2624 -2202 2673
rect 3999 2625 4023 2670
rect -1492 2611 -1463 2615
rect -1467 2529 -1463 2611
rect -1479 2525 -1463 2529
rect 3263 2611 3292 2615
rect 3263 2527 3267 2611
rect 3263 2523 3279 2527
rect -2216 2334 -2187 2374
rect 4001 2328 4028 2367
rect -1493 2311 -1471 2315
rect -1475 2226 -1471 2311
rect -1481 2222 -1471 2226
rect 3266 2311 3292 2315
rect 3266 2228 3270 2311
rect 3266 2224 3281 2228
rect -1476 2215 -594 2216
rect -1476 2206 -614 2215
rect -595 2206 -594 2215
rect -1476 2205 -594 2206
rect -2211 2063 -2189 2067
rect -2216 2028 -2185 2063
rect -1476 2055 -1465 2205
rect -1495 2044 -1465 2055
rect 4003 2020 4036 2074
rect 3262 2011 3292 2015
rect 3262 1927 3266 2011
rect 3262 1923 3280 1927
rect -2216 1725 -2181 1774
rect -2218 1425 -2190 1467
rect 3992 1433 4025 1470
rect 3261 1411 3292 1415
rect 3261 1327 3265 1411
rect 3261 1323 3281 1327
rect -2213 1133 -2190 1163
rect 4000 1129 4032 1170
rect 3271 1111 3292 1115
rect 3271 1028 3275 1111
rect 3271 1024 3279 1028
rect -2212 860 -2190 864
rect -2212 836 -2189 860
rect -2208 822 -2189 836
rect 4003 833 4028 868
rect 3264 811 3292 815
rect 3264 727 3268 811
rect 3264 723 3279 727
rect 4004 563 4030 574
rect -2216 527 -2192 561
rect 3991 524 4036 563
rect 4004 523 4030 524
rect 3268 511 3292 515
rect 3268 427 3272 511
rect 3268 423 3280 427
rect 3999 231 4032 288
rect 3264 211 3292 215
rect 3264 127 3268 211
rect 3264 123 3281 127
rect -1481 71 -1472 75
rect -1476 -11 -1472 71
rect -1492 -15 -1472 -11
rect -2227 -66 -2189 -32
rect -2232 -375 -2200 -331
rect 4001 -370 4034 -324
rect -1492 -389 -1464 -385
rect -1468 -473 -1464 -389
rect -1480 -477 -1464 -473
rect 3272 -389 3292 -385
rect 3272 -473 3276 -389
rect 3272 -477 3281 -473
rect -2222 -675 -2191 -632
rect -1493 -689 -1471 -685
rect -1475 -772 -1471 -689
rect -1481 -776 -1471 -772
rect -2217 -933 -2191 -932
rect -2217 -934 -2188 -933
rect -2220 -966 -2188 -934
rect -2217 -969 -2188 -966
rect -2217 -972 -2191 -969
rect -1492 -989 -1461 -985
rect -1465 -1072 -1461 -989
rect -1480 -1076 -1461 -1072
rect -2215 -1277 -2190 -1232
rect -1492 -1289 -1472 -1285
rect -1476 -1370 -1472 -1289
rect -1480 -1374 -1472 -1370
rect -165 -1407 -142 -591
rect 3999 -666 4027 -629
rect 3265 -689 3293 -685
rect 3265 -773 3269 -689
rect 3265 -777 3279 -773
rect 3274 -989 3292 -985
rect 4007 -988 4031 -921
rect 3274 -1079 3278 -989
rect 3282 -1079 3286 -1076
rect 3274 -1083 3286 -1079
rect 3988 -1269 4024 -1227
rect 3268 -1289 3292 -1285
rect 3268 -1372 3272 -1289
rect 3268 -1376 3279 -1372
rect 430 -2097 472 -2093
rect -1382 -2130 -1313 -2100
rect -1078 -2122 -1022 -2101
rect -777 -2133 -725 -2103
rect -475 -2105 -426 -2103
rect -475 -2130 -420 -2105
rect -159 -2110 -134 -2097
rect -475 -2131 -426 -2130
rect 130 -2131 180 -2107
rect 425 -2134 484 -2097
rect 723 -2122 766 -2095
rect 1015 -2133 1073 -2107
rect 1333 -2121 1338 -2099
rect 1926 -2129 1974 -2104
rect 2225 -2129 2269 -2104
rect 2522 -2128 2583 -2105
rect 2821 -2130 2874 -2101
rect 3121 -2127 3177 -2104
<< m2contact >>
rect -1478 3381 -1472 3387
rect -1178 3378 -1172 3384
rect -877 3381 -871 3387
rect -577 3379 -571 3385
rect -277 3379 -271 3385
rect 23 3379 29 3385
rect 622 3380 628 3386
rect 922 3380 928 3386
rect 1222 3381 1228 3387
rect 1522 3379 1528 3385
rect 1822 3380 1828 3386
rect 2122 3380 2128 3386
rect 2722 3379 2728 3385
rect 3022 3380 3028 3386
rect -1487 3123 -1481 3129
rect 3280 3122 3286 3128
rect -1486 2823 -1480 2829
rect -1485 2524 -1479 2530
rect 3279 2522 3285 2528
rect -1487 2221 -1481 2227
rect 3281 2223 3287 2229
rect -614 2206 -595 2215
rect 3280 1922 3286 1928
rect 3281 1322 3287 1328
rect 3279 1023 3285 1029
rect 3279 722 3285 728
rect 3280 422 3286 428
rect 3281 122 3287 128
rect -1487 70 -1481 76
rect -1486 -478 -1480 -472
rect 3281 -478 3287 -472
rect -1487 -777 -1481 -771
rect -1486 -1077 -1480 -1071
rect -1486 -1375 -1480 -1369
rect 3279 -778 3285 -772
rect 3281 -1076 3287 -1070
rect 3279 -1377 3285 -1371
<< metal2 >>
rect -1450 3177 -1447 3386
rect -1152 3183 -1149 3384
rect -853 3190 -850 3384
rect -555 3197 -552 3384
rect -254 3207 -251 3385
rect 48 3216 51 3385
rect 645 3232 650 3387
rect 947 3251 952 3388
rect 1248 3271 1253 3387
rect 1544 3294 1549 3389
rect 1846 3313 1851 3390
rect 2145 3330 2150 3385
rect 2747 3348 2752 3387
rect 3048 3366 3053 3388
rect 3048 3361 3117 3366
rect 2747 3343 3103 3348
rect 2145 3325 3086 3330
rect 1846 3308 3067 3313
rect 1544 3289 3051 3294
rect 1248 3266 3034 3271
rect 947 3246 3017 3251
rect 645 3227 3002 3232
rect 48 3213 2193 3216
rect -254 3204 1969 3207
rect -555 3194 1913 3197
rect -853 3187 1345 3190
rect -1152 3180 1297 3183
rect -1450 3174 1201 3177
rect -1450 3157 1129 3160
rect -1450 3149 -1447 3157
rect -1485 3146 -1447 3149
rect -1437 3142 969 3145
rect -1437 2851 -1434 3142
rect -1486 2848 -1434 2851
rect -1417 3131 945 3134
rect -1417 2553 -1414 3131
rect -1484 2550 -1414 2553
rect -1396 3117 817 3120
rect -1396 2253 -1393 3117
rect -1487 2250 -1393 2253
rect -1388 3109 737 3112
rect -1486 1872 -1473 1876
rect -1477 1805 -1473 1872
rect -1388 1822 -1385 3109
rect -1374 3099 657 3102
rect -1374 1819 -1371 3099
rect -1359 3090 513 3093
rect -1359 1821 -1356 3090
rect -1345 3084 497 3087
rect -1345 1820 -1342 3084
rect -1327 3077 481 3080
rect -1327 1819 -1324 3077
rect 478 2417 481 3077
rect 494 2417 497 3084
rect 510 2417 513 3090
rect 654 2417 657 3099
rect 734 2417 737 3109
rect 814 2417 817 3117
rect 942 2417 945 3131
rect 966 2417 969 3142
rect 1126 2417 1129 3157
rect 1198 2417 1201 3174
rect 1294 2417 1297 3180
rect 1342 2417 1345 3187
rect 1910 2417 1913 3194
rect 1966 2417 1969 3204
rect 2190 2417 2193 3213
rect -595 2206 -594 2215
rect 2997 2157 3002 3227
rect 2445 2152 2446 2157
rect 2451 2152 3002 2157
rect 3012 1987 3017 3246
rect 2445 1982 3017 1987
rect -1492 1801 -1473 1805
rect -1467 1792 -672 1797
rect -1467 1641 -1462 1792
rect 3029 1707 3034 3266
rect 2449 1702 3034 1707
rect -1488 1636 -1462 1641
rect -1466 1592 -666 1597
rect -1466 1563 -1461 1592
rect -1489 1558 -1461 1563
rect -1456 1512 -669 1517
rect -1492 1395 -1466 1399
rect -1470 1327 -1466 1395
rect -1485 1323 -1466 1327
rect -1456 1265 -1451 1512
rect -1486 1260 -1451 1265
rect -1445 1492 -667 1497
rect -1492 1095 -1459 1099
rect -1463 1028 -1459 1095
rect -1484 1024 -1459 1028
rect -1445 966 -1440 1492
rect 2450 1392 2571 1397
rect -1487 961 -1440 966
rect -1434 1382 -667 1387
rect -1492 795 -1455 799
rect -1459 729 -1455 795
rect -1488 725 -1455 729
rect -1434 666 -1429 1382
rect -1488 661 -1429 666
rect -1492 495 -1461 499
rect -1465 427 -1461 495
rect -1486 423 -1461 427
rect -1388 54 -1385 1349
rect -1487 51 -1385 54
rect -1374 -450 -1371 1346
rect -1485 -453 -1371 -450
rect -1359 -749 -1356 1345
rect -1485 -752 -1356 -749
rect -1345 -1049 -1342 1344
rect -1316 1343 -677 1346
rect -1485 -1052 -1342 -1049
rect -1327 -1057 -1324 1342
rect -1458 -1060 -1324 -1057
rect -1458 -1348 -1455 -1060
rect -1485 -1351 -1455 -1348
rect -1316 -1364 -1313 1343
rect 2450 1302 2560 1307
rect 2448 1142 2544 1147
rect 2449 1052 2529 1057
rect 2449 922 2518 927
rect 2448 902 2508 907
rect 2446 832 2491 837
rect 2450 762 2481 767
rect 2449 742 2470 747
rect 2449 702 2461 707
rect 2456 607 2461 702
rect 2465 616 2470 742
rect 2476 625 2481 762
rect 2486 634 2491 832
rect 2503 647 2508 902
rect 2513 658 2518 922
rect 2524 668 2529 1052
rect 2539 683 2544 1142
rect 2555 695 2560 1302
rect 2566 706 2571 1392
rect 3046 706 3051 3289
rect 2566 701 3051 706
rect 3062 695 3067 3308
rect 2555 690 3067 695
rect 3081 683 3086 3325
rect 2539 678 3086 683
rect 3098 668 3103 3343
rect 2524 663 3103 668
rect 3112 658 3117 3361
rect 2513 653 3117 658
rect 3125 3145 3284 3150
rect 3125 647 3130 3145
rect 2503 642 3130 647
rect 3141 3059 3287 3064
rect 3141 634 3146 3059
rect 3268 2895 3292 2899
rect 3268 2828 3272 2895
rect 3268 2824 3286 2828
rect 2486 629 3146 634
rect 3151 2547 3285 2552
rect 3151 625 3156 2547
rect 2476 620 3156 625
rect 3162 2246 3285 2251
rect 3162 616 3167 2246
rect 2465 611 3167 616
rect 3173 1945 3286 1950
rect 3173 607 3178 1945
rect 2456 602 3178 607
rect 3187 1344 3286 1349
rect 3187 597 3192 1344
rect 2447 592 3192 597
rect 3199 1045 3287 1050
rect 3199 507 3204 1045
rect 2449 502 3204 507
rect 3214 743 3285 748
rect 3214 397 3219 743
rect 2449 392 3219 397
rect 3231 443 3285 448
rect 2450 356 2534 357
rect 3231 356 3236 443
rect 2450 352 3236 356
rect 2530 351 3236 352
rect 2459 332 2523 337
rect 2452 302 2514 307
rect 2453 282 2505 287
rect 2451 192 2493 197
rect 2448 162 2449 167
rect 2454 162 2482 167
rect 2456 102 2469 107
rect 2450 -138 2459 -133
rect -402 -1330 -399 -617
rect -937 -1333 -399 -1330
rect -1176 -1358 -1101 -1354
rect -1316 -1367 -1237 -1364
rect -1466 -1377 -1401 -1373
rect -1466 -1381 -1462 -1377
rect -1474 -1385 -1462 -1381
rect -1405 -1392 -1401 -1377
rect -1240 -1387 -1237 -1367
rect -1176 -1389 -1172 -1358
rect -1105 -1392 -1101 -1358
rect -937 -1386 -934 -1333
rect -330 -1340 -327 -617
rect -638 -1343 -327 -1340
rect -875 -1369 -801 -1365
rect -875 -1386 -871 -1369
rect -805 -1392 -801 -1369
rect -638 -1388 -635 -1343
rect -210 -1351 -207 -617
rect 926 -630 929 -617
rect -338 -1354 -207 -1351
rect 262 -633 929 -630
rect -576 -1367 -501 -1363
rect -576 -1384 -572 -1367
rect -505 -1394 -501 -1367
rect -338 -1386 -335 -1354
rect 24 -1368 99 -1364
rect 24 -1385 28 -1368
rect 95 -1392 99 -1368
rect 262 -1387 265 -633
rect 1070 -643 1073 -617
rect 561 -646 1073 -643
rect 324 -1369 399 -1365
rect 324 -1388 328 -1369
rect 395 -1392 399 -1369
rect 561 -1386 564 -646
rect 1102 -652 1105 -617
rect 859 -655 1105 -652
rect 623 -1365 699 -1361
rect 623 -1386 627 -1365
rect 695 -1392 699 -1365
rect 859 -1386 862 -655
rect 925 -1369 999 -1365
rect 925 -1386 929 -1369
rect 995 -1392 999 -1369
rect 1142 -1368 1145 -617
rect 1174 -1347 1177 -616
rect 1222 -1339 1225 -617
rect 2198 -1328 2201 -617
rect 2454 -1307 2459 -138
rect 2464 -1295 2469 102
rect 2477 -1284 2482 162
rect 2488 -1047 2493 192
rect 2500 -746 2505 282
rect 2509 -446 2514 302
rect 2517 150 2522 332
rect 2517 145 3283 150
rect 2509 -451 3286 -446
rect 2500 -751 3283 -746
rect 3278 -756 3283 -751
rect 2488 -1052 3285 -1047
rect 2477 -1289 3274 -1284
rect 2464 -1300 3264 -1295
rect 2454 -1312 2964 -1307
rect 2198 -1331 2660 -1328
rect 1222 -1342 2360 -1339
rect 1174 -1350 2061 -1347
rect 1142 -1371 1164 -1368
rect 1161 -1387 1164 -1371
rect 1223 -1371 1299 -1367
rect 1223 -1387 1227 -1371
rect 1295 -1392 1299 -1371
rect 1825 -1369 1899 -1365
rect 1825 -1387 1829 -1369
rect 1895 -1392 1899 -1369
rect 2058 -1387 2061 -1350
rect 2124 -1366 2199 -1362
rect 2124 -1387 2128 -1366
rect 2195 -1392 2199 -1366
rect 2357 -1385 2360 -1342
rect 2425 -1366 2499 -1362
rect 2425 -1389 2429 -1366
rect 2495 -1392 2499 -1366
rect 2657 -1384 2660 -1331
rect 2724 -1365 2799 -1361
rect 2724 -1385 2728 -1365
rect 2795 -1392 2799 -1365
rect 2959 -1387 2964 -1312
rect 3025 -1365 3099 -1361
rect 3025 -1387 3029 -1365
rect 3095 -1392 3099 -1365
rect 3259 -1386 3264 -1300
rect 3269 -1351 3274 -1289
rect 3269 -1356 3285 -1351
<< m3contact >>
rect -1389 1817 -1384 1822
rect -1375 1814 -1370 1819
rect -1360 1816 -1355 1821
rect -1346 1815 -1341 1820
rect 2446 2152 2451 2157
rect 2440 1982 2445 1987
rect -1328 1814 -1323 1819
rect -672 1792 -667 1797
rect 2444 1702 2449 1707
rect -666 1592 -661 1597
rect -669 1512 -664 1517
rect -667 1492 -662 1497
rect 2445 1392 2450 1397
rect -667 1382 -662 1387
rect -1389 1349 -1384 1354
rect -1375 1346 -1370 1351
rect -1360 1345 -1355 1350
rect -1346 1344 -1341 1349
rect -1328 1342 -1323 1347
rect -677 1342 -672 1347
rect 2445 1302 2450 1307
rect 2443 1142 2448 1147
rect 2444 1052 2449 1057
rect 2444 922 2449 927
rect 2443 902 2448 907
rect 2441 832 2446 837
rect 2445 762 2450 767
rect 2444 742 2449 747
rect 2444 702 2449 707
rect 2442 592 2447 597
rect 2444 502 2449 507
rect 2444 392 2449 397
rect 2445 352 2450 357
rect 2454 332 2459 337
rect 2447 302 2452 307
rect 2448 282 2453 287
rect 2446 192 2451 197
rect 2449 162 2454 167
rect 2451 102 2456 107
rect 2445 -138 2450 -133
<< metal3 >>
rect 2445 2157 2452 2158
rect 2430 2152 2446 2157
rect 2451 2152 2452 2157
rect 2445 2151 2452 2152
rect 2439 1987 2446 1988
rect 2431 1982 2440 1987
rect 2445 1982 2446 1987
rect 2439 1981 2446 1982
rect -1390 1822 -1383 1823
rect -1390 1817 -1389 1822
rect -1384 1817 -1383 1822
rect -1361 1821 -1354 1822
rect -1390 1816 -1383 1817
rect -1376 1819 -1369 1820
rect -1389 1355 -1384 1816
rect -1376 1814 -1375 1819
rect -1370 1814 -1369 1819
rect -1361 1816 -1360 1821
rect -1355 1816 -1354 1821
rect -1361 1815 -1354 1816
rect -1347 1820 -1340 1821
rect -1347 1815 -1346 1820
rect -1341 1815 -1340 1820
rect -1376 1813 -1369 1814
rect -1390 1354 -1383 1355
rect -1390 1349 -1389 1354
rect -1384 1349 -1383 1354
rect -1375 1352 -1370 1813
rect -1390 1348 -1383 1349
rect -1376 1351 -1369 1352
rect -1360 1351 -1355 1815
rect -1347 1814 -1340 1815
rect -1329 1819 -1322 1820
rect -1329 1814 -1328 1819
rect -1323 1814 -1322 1819
rect -1376 1346 -1375 1351
rect -1370 1346 -1369 1351
rect -1376 1345 -1369 1346
rect -1361 1350 -1354 1351
rect -1346 1350 -1341 1814
rect -1329 1813 -1322 1814
rect -1361 1345 -1360 1350
rect -1355 1345 -1354 1350
rect -1361 1344 -1354 1345
rect -1347 1349 -1340 1350
rect -1347 1344 -1346 1349
rect -1341 1344 -1340 1349
rect -1328 1348 -1323 1813
rect -673 1797 -666 1798
rect -673 1792 -672 1797
rect -667 1792 -647 1797
rect -673 1791 -666 1792
rect 2443 1707 2450 1708
rect 2431 1702 2444 1707
rect 2449 1702 2450 1707
rect 2443 1701 2450 1702
rect -667 1597 -660 1598
rect -667 1592 -666 1597
rect -661 1592 -647 1597
rect -667 1591 -660 1592
rect -670 1517 -663 1518
rect -670 1512 -669 1517
rect -664 1512 -647 1517
rect -670 1511 -663 1512
rect -668 1497 -661 1498
rect -668 1492 -667 1497
rect -662 1492 -647 1497
rect -668 1491 -661 1492
rect 2444 1397 2451 1398
rect 2431 1392 2445 1397
rect 2450 1392 2451 1397
rect 2444 1391 2451 1392
rect -668 1387 -661 1388
rect -668 1382 -667 1387
rect -662 1382 -647 1387
rect -668 1381 -661 1382
rect -1347 1343 -1340 1344
rect -1329 1347 -1322 1348
rect -1329 1342 -1328 1347
rect -1323 1342 -1322 1347
rect -1329 1341 -1322 1342
rect -678 1347 -671 1348
rect -678 1342 -677 1347
rect -672 1342 -647 1347
rect -678 1341 -671 1342
rect 2444 1307 2451 1308
rect 2431 1302 2445 1307
rect 2450 1302 2451 1307
rect 2444 1301 2451 1302
rect 2442 1147 2449 1148
rect 2431 1142 2443 1147
rect 2448 1142 2449 1147
rect 2442 1141 2449 1142
rect 2443 1057 2450 1058
rect 2431 1052 2444 1057
rect 2449 1052 2450 1057
rect 2443 1051 2450 1052
rect 2443 927 2450 928
rect 2431 922 2444 927
rect 2449 922 2450 927
rect 2443 921 2450 922
rect 2442 907 2449 908
rect 2431 902 2443 907
rect 2448 902 2449 907
rect 2442 901 2449 902
rect 2440 837 2447 838
rect 2431 832 2441 837
rect 2446 832 2447 837
rect 2440 831 2447 832
rect 2444 767 2451 768
rect 2431 762 2445 767
rect 2450 762 2451 767
rect 2444 761 2451 762
rect 2443 747 2450 748
rect 2431 742 2444 747
rect 2449 742 2450 747
rect 2443 741 2450 742
rect 2443 707 2450 708
rect 2431 702 2444 707
rect 2449 702 2450 707
rect 2443 701 2450 702
rect 2441 597 2448 598
rect 2431 592 2442 597
rect 2447 592 2448 597
rect 2441 591 2448 592
rect 2443 507 2450 508
rect 2431 502 2444 507
rect 2449 502 2450 507
rect 2443 501 2450 502
rect 2443 397 2450 398
rect 2429 392 2444 397
rect 2449 392 2450 397
rect 2443 391 2450 392
rect 2444 357 2451 358
rect 2431 352 2445 357
rect 2450 352 2451 357
rect 2444 351 2451 352
rect 2453 337 2460 338
rect 2431 332 2454 337
rect 2459 332 2460 337
rect 2453 331 2460 332
rect 2446 307 2453 308
rect 2430 302 2447 307
rect 2452 302 2453 307
rect 2446 301 2453 302
rect 2447 287 2454 288
rect 2431 282 2448 287
rect 2453 282 2454 287
rect 2447 281 2454 282
rect 2445 197 2452 198
rect 2431 192 2446 197
rect 2451 192 2452 197
rect 2445 191 2452 192
rect 2448 167 2455 168
rect 2431 162 2449 167
rect 2454 162 2455 167
rect 2448 161 2455 162
rect 2450 107 2457 108
rect 2431 102 2451 107
rect 2456 102 2457 107
rect 2450 101 2457 102
rect 2444 -133 2451 -132
rect 2429 -138 2445 -133
rect 2450 -138 2451 -133
rect 2444 -139 2451 -138
use PadFC  16_0
timestamp 1681001061
transform 1 0 -2500 0 1 3400
box 327 -3 1003 673
use PadFC  16_1
timestamp 1681001061
transform 0 1 3300 -1 0 4400
box 327 -3 1003 673
use PadFC  16_2
timestamp 1681001061
transform 0 -1 -1500 1 0 -2400
box 327 -3 1003 673
use PadFC  16_3
timestamp 1681001061
transform -1 0 4300 0 -1 -1400
box 327 -3 1003 673
use PadBiDir  17_0
timestamp 1711830429
transform 1 0 -1500 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_1
timestamp 1711830429
transform 1 0 -1200 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_2
timestamp 1711830429
transform 1 0 -900 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_3
timestamp 1711830429
transform 1 0 -600 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_4
timestamp 1711830429
transform 1 0 -300 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_5
timestamp 1711830429
transform 1 0 0 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_6
timestamp 1711830429
transform 1 0 600 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_7
timestamp 1711830429
transform 1 0 900 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_8
timestamp 1711830429
transform 1 0 1200 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_9
timestamp 1711830429
transform 0 -1 -1500 1 0 3100
box -36 -19 303 1000
use PadBiDir  17_10
timestamp 1711830429
transform 0 -1 -1500 1 0 2800
box -36 -19 303 1000
use PadBiDir  17_11
timestamp 1711830429
transform 0 -1 -1500 1 0 2500
box -36 -19 303 1000
use PadBiDir  17_12
timestamp 1711830429
transform 0 -1 -1500 1 0 2200
box -36 -19 303 1000
use PadBiDir  17_13
timestamp 1711830429
transform 0 -1 -1500 -1 0 1900
box -36 -19 303 1000
use PadBiDir  17_14
timestamp 1711830429
transform 0 -1 -1500 1 0 -500
box -36 -19 303 1000
use PadBiDir  17_15
timestamp 1711830429
transform 0 -1 -1500 1 0 -800
box -36 -19 303 1000
use PadBiDir  17_16
timestamp 1711830429
transform 0 -1 -1500 1 0 -1100
box -36 -19 303 1000
use PadBiDir  17_17
timestamp 1711830429
transform 0 1 3300 1 0 3100
box -36 -19 303 1000
use PadBiDir  17_18
timestamp 1711830429
transform 0 1 3300 1 0 2800
box -36 -19 303 1000
use PadBiDir  17_19
timestamp 1711830429
transform 0 1 3300 1 0 2500
box -36 -19 303 1000
use PadBiDir  17_20
timestamp 1711830429
transform 0 1 3300 1 0 2200
box -36 -19 303 1000
use PadBiDir  17_21
timestamp 1711830429
transform 0 1 3300 1 0 1900
box -36 -19 303 1000
use PadBiDir  17_22
timestamp 1711830429
transform 0 1 3300 1 0 -500
box -36 -19 303 1000
use PadBiDir  17_23
timestamp 1711830429
transform 0 1 3300 1 0 -800
box -36 -19 303 1000
use PadBiDir  17_24
timestamp 1711830429
transform 0 1 3300 1 0 -1100
box -36 -19 303 1000
use PadBiDir  17_25
timestamp 1711830429
transform 0 -1 -1500 1 0 -1400
box -36 -19 303 1000
use PadBiDir  17_26
timestamp 1711830429
transform 1 0 -1500 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_27
timestamp 1711830429
transform 1 0 -1200 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_28
timestamp 1711830429
transform 1 0 -900 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_29
timestamp 1711830429
transform 1 0 -600 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_30
timestamp 1711830429
transform 1 0 0 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_31
timestamp 1711830429
transform 1 0 300 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_32
timestamp 1711830429
transform 1 0 600 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_33
timestamp 1711830429
transform 1 0 900 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_34
timestamp 1711830429
transform 0 1 3300 1 0 -1400
box -36 -19 303 1000
use PadBiDir  17_35
timestamp 1711830429
transform 1 0 1200 0 -1 -1400
box -36 -19 303 1000
use PadVdd  18_0
timestamp 1711831643
transform 1 0 300 0 1 3400
box -3 -16 303 1000
use PadVdd  18_1
timestamp 1711831643
transform 1 0 -300 0 -1 -1400
box -3 -16 303 1000
use PadGnd  19_0
timestamp 1711831454
transform 0 -1 -1500 -1 0 2200
box -3 -11 303 1000
use PadGnd  19_1
timestamp 1711831454
transform 0 1 3300 -1 0 1900
box -3 -11 303 1000
use PadBiDir  PadBiDir_0
timestamp 1711830429
transform 1 0 1500 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_1
timestamp 1711830429
transform 1 0 1800 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_2
timestamp 1711830429
transform 1 0 2100 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_3
timestamp 1711830429
transform 1 0 2700 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_4
timestamp 1711830429
transform 1 0 3000 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_5
timestamp 1711830429
transform 1 0 1800 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_6
timestamp 1711830429
transform 1 0 2100 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_7
timestamp 1711830429
transform 1 0 2400 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_8
timestamp 1711830429
transform 1 0 2700 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_9
timestamp 1711830429
transform 1 0 3000 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_10
timestamp 1711830429
transform 0 -1 -1500 -1 0 100
box -36 -19 303 1000
use PadBiDir  PadBiDir_11
timestamp 1711830429
transform 0 -1 -1500 1 0 400
box -36 -19 303 1000
use PadBiDir  PadBiDir_12
timestamp 1711830429
transform 0 -1 -1500 1 0 700
box -36 -19 303 1000
use PadBiDir  PadBiDir_13
timestamp 1711830429
transform 0 -1 -1500 1 0 1000
box -36 -19 303 1000
use PadBiDir  PadBiDir_14
timestamp 1711830429
transform 0 -1 -1500 1 0 1300
box -36 -19 303 1000
use PadBiDir  PadBiDir_15
timestamp 1711830429
transform 0 1 3300 1 0 100
box -36 -19 303 1000
use PadBiDir  PadBiDir_16
timestamp 1711830429
transform 0 1 3300 1 0 400
box -36 -19 303 1000
use PadBiDir  PadBiDir_17
timestamp 1711830429
transform 0 1 3300 1 0 700
box -36 -19 303 1000
use PadBiDir  PadBiDir_18
timestamp 1711830429
transform 0 1 3300 1 0 1000
box -36 -19 303 1000
use PadBiDir  PadBiDir_19
timestamp 1711830429
transform 0 1 3300 1 0 1300
box -36 -19 303 1000
use PadGnd  PadGnd_0
timestamp 1711831454
transform 0 -1 -1500 -1 0 400
box -3 -11 303 1000
use PadGnd  PadGnd_1
timestamp 1711831454
transform 0 1 3300 -1 0 100
box -3 -11 303 1000
use PadVdd  PadVdd_0
timestamp 1711831643
transform 1 0 2400 0 1 3400
box -3 -16 303 1000
use PadVdd  PadVdd_1
timestamp 1711831643
transform 1 0 1500 0 -1 -1400
box -3 -16 303 1000
use top_module  top_module_0
timestamp 1713400504
transform 1 0 -652 0 1 -620
box 0 0 3088 3040
<< labels >>
rlabel metal1 -147 -2104 -147 -2104 1 Vdd
rlabel metal1 -2199 1754 -2199 1754 1 p_in_incr[2]
rlabel metal1 -2205 1442 -2205 1442 1 p_in_incr[1]
rlabel metal1 -2200 1148 -2200 1148 1 p_in_mult[2]
rlabel metal1 -2201 848 -2201 848 1 p_in_mult[1]
rlabel metal1 -2204 542 -2204 542 1 p_in_mult[0]
rlabel metal1 -449 -2119 -449 -2119 1 p_in_n_mines[2]
rlabel metal1 -757 -2115 -757 -2115 1 p_in_n_mines[0]
rlabel metal1 -1048 -2110 -1048 -2110 1 p_in_n_mines[1]
rlabel metal1 156 -2119 156 -2119 1 p_in_clkb
rlabel metal1 449 -2109 449 -2109 1 p_in_data[2]
rlabel metal1 742 -2107 742 -2107 1 p_in_data[1]
rlabel metal1 1045 -2120 1045 -2120 1 p_in_data[0]
rlabel metal1 2248 -2118 2248 -2118 1 p_in_data[4]
rlabel metal1 1949 -2117 1949 -2117 1 p_in_data[3]
rlabel metal1 2552 -2117 2552 -2117 1 p_in_place
rlabel metal1 2843 -2116 2843 -2116 1 p_in_data_in
rlabel metal1 3146 -2115 3146 -2115 1 p_in_restart
rlabel metal1 4008 -1250 4008 -1250 1 out_global_score[6]
rlabel metal1 4017 -952 4017 -952 1 p_global_score[5]
rlabel metal1 4012 -649 4012 -649 1 p_out_gameover
rlabel metal1 4017 -347 4017 -347 1 p_out_n_nearby[1]
rlabel metal1 4010 258 4010 258 1 p_out_global_score[7]
rlabel metal1 4012 545 4012 545 1 p_out_n_nearby[0]
rlabel metal1 4008 1449 4008 1449 1 p_out_global_score[2]
rlabel metal1 4016 1146 4016 1146 1 p_out_global_score[3]
rlabel metal1 4016 847 4016 847 1 p_out_global_score[4]
rlabel metal1 4018 2046 4018 2046 1 p_out_global_score[1]
rlabel metal1 4015 2346 4015 2346 1 p_out_win
rlabel metal1 4012 2647 4012 2647 1 p_out_global_score[0]
rlabel metal1 4016 2946 4016 2946 1 p_in_clka
rlabel metal1 4007 3249 4007 3249 1 p_out_temp_cleared[4]
rlabel metal1 3145 4107 3145 4107 1 p_out_temp_cleared[3]
rlabel metal1 2846 4108 2846 4108 1 p_out_temp_cleared[0]
rlabel metal1 2249 4117 2249 4117 1 p_out_temp_cleared[1]
rlabel metal1 1951 4109 1952 4110 1 p_out_temp_cleared[24]
rlabel metal1 1646 4114 1646 4114 1 p_out_temp_cleared[5]
rlabel metal1 1347 4110 1347 4110 1 p_out_temp_cleared[6]
rlabel metal1 746 4102 746 4102 1 p_out_temp_cleared[8]
rlabel metal1 1049 4107 1049 4107 1 p_out_temp_cleared[7]
rlabel metal1 150 4101 150 4101 1 p_out_temp_cleared[9]
rlabel metal1 -153 4117 -153 4117 1 p_out_temp_cleared[10]
rlabel metal1 -452 4105 -452 4105 1 p_out_temp_cleared[11]
rlabel metal1 -752 4109 -751 4109 1 p_out_temp_cleared[12]
rlabel metal1 -1057 4108 -1057 4108 1 p_out_temp_cleared[23]
rlabel metal1 -1361 4115 -1361 4115 1 p_out_temp_cleared[13]
rlabel metal1 -2209 3246 -2208 3246 1 p_out_temp_cleared[14]
rlabel metal1 -2209 2950 -2209 2950 1 p_out_temp_cleared[22]
rlabel metal1 -2214 2647 -2214 2647 1 p_out_temp_cleared[20]
rlabel metal1 -2201 2352 -2201 2352 1 p_out_temp_cleared[21]
rlabel metal1 -2210 -50 -2210 -50 1 p_out_temp_cleared[19]
rlabel metal1 -2219 -355 -2219 -355 1 p_out_temp_cleared[18]
rlabel metal1 -2207 -656 -2207 -656 1 p_out_temp_cleared[15]
rlabel metal1 -2204 -953 -2204 -953 1 p_out_temp_cleared[17]
rlabel metal1 -2204 -1256 -2204 -1256 1 p_out_temp_cleared[16]
rlabel metal1 -1349 -2115 -1349 -2115 1 p_in_incr[0]
rlabel metal1 -2201 2045 -2201 2046 1 GND!
<< end >>
