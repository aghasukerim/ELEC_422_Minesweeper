magic
tech scmos
timestamp 1713592123
<< nwell >>
rect -5 48 53 105
rect 6 44 33 48
<< ntransistor >>
rect 7 10 9 20
rect 15 10 17 30
rect 20 10 22 30
rect 28 10 30 30
rect 33 10 35 30
<< ptransistor >>
rect 7 70 9 90
rect 15 50 17 90
rect 20 50 22 90
rect 28 54 30 94
rect 33 54 35 94
<< ndiffusion >>
rect 12 28 15 30
rect 10 26 15 28
rect 2 19 7 20
rect 6 10 7 19
rect 9 12 10 20
rect 14 12 15 26
rect 9 10 15 12
rect 17 10 20 30
rect 22 26 28 30
rect 22 12 23 26
rect 27 12 28 26
rect 22 10 28 12
rect 30 10 33 30
rect 35 29 40 30
rect 35 10 36 29
<< pdiffusion >>
rect 23 92 28 94
rect 2 89 7 90
rect 6 70 7 89
rect 9 70 10 90
rect 14 56 15 90
rect 12 50 15 56
rect 17 50 20 90
rect 22 58 23 90
rect 27 58 28 92
rect 22 54 28 58
rect 30 54 33 94
rect 35 93 40 94
rect 35 54 36 93
rect 22 50 25 54
<< ndcontact >>
rect 2 10 6 19
rect 10 12 14 26
rect 23 12 27 26
rect 36 10 40 29
<< pdcontact >>
rect 2 70 6 89
rect 10 56 14 90
rect 23 58 27 92
rect 36 54 40 93
<< psubstratepcontact >>
rect -2 -2 2 2
rect 14 -2 18 2
rect 30 -2 34 2
<< nsubstratencontact >>
rect -2 98 2 102
rect 14 98 18 102
rect 30 98 34 102
<< polysilicon >>
rect 7 95 22 97
rect 7 90 9 95
rect 15 90 17 92
rect 20 90 22 95
rect 28 94 30 96
rect 33 94 35 96
rect 7 69 9 70
rect 4 67 9 69
rect 4 43 6 67
rect 15 49 17 50
rect 12 47 17 49
rect 20 48 22 50
rect 12 43 14 47
rect 28 40 30 54
rect 33 53 35 54
rect 33 51 36 53
rect 4 23 6 39
rect 11 33 13 39
rect 25 38 30 40
rect 20 34 24 36
rect 11 31 17 33
rect 15 30 17 31
rect 20 30 22 34
rect 34 33 36 47
rect 28 30 30 32
rect 33 31 36 33
rect 33 30 35 31
rect 4 21 9 23
rect 7 20 9 21
rect 7 5 9 10
rect 15 8 17 10
rect 20 8 22 10
rect 28 5 30 10
rect 33 8 35 10
rect 7 3 30 5
<< polycontact >>
rect 2 39 6 43
rect 10 39 14 43
rect 21 36 25 40
rect 34 47 38 51
<< metal1 >>
rect -2 102 50 103
rect 2 98 14 102
rect 18 98 30 102
rect 34 98 50 102
rect -2 97 50 98
rect 10 90 14 97
rect 2 89 6 90
rect 2 53 5 70
rect 23 92 27 94
rect 36 93 40 97
rect 27 58 31 59
rect 23 56 31 58
rect 2 50 21 53
rect 2 43 6 47
rect 10 43 14 47
rect 18 36 21 50
rect 28 37 31 56
rect 34 43 38 47
rect 18 34 23 36
rect 2 31 23 34
rect 28 33 38 37
rect 2 20 5 31
rect 28 30 31 33
rect 27 28 31 30
rect 10 26 14 28
rect 2 19 6 20
rect 10 3 14 12
rect 23 26 31 28
rect 27 25 31 26
rect 36 29 40 30
rect 23 10 27 12
rect 36 3 40 10
rect -2 2 50 3
rect 2 -2 14 2
rect 18 -2 30 2
rect 34 -2 50 2
rect -2 -3 50 -2
<< m1p >>
rect 2 43 6 47
rect 10 43 14 47
rect 34 43 38 47
rect 34 33 38 37
<< labels >>
rlabel metal1 4 45 4 45 4 S
rlabel metal1 4 100 4 100 4 vdd
rlabel metal1 4 0 4 0 4 gnd
rlabel metal1 36 35 36 35 4 Y
rlabel metal1 36 45 36 45 4 A
rlabel metal1 12 45 12 45 4 B
<< end >>
