magic
tech scmos
timestamp 1710899220
<< m2contact >>
rect -2 -2 2 2
<< end >>
