magic
tech scmos
timestamp 1713293539
use PadFrame64  PadFrame64_0
timestamp 1711836921
transform 1 0 2500 0 1 2400
box -2500 -2400 4300 4400
use top_module  top_module_0
timestamp 1710899220
transform 1 0 1948 0 1 2427
box 14 13 2730 2627
<< end >>
