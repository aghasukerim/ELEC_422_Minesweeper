magic
tech scmos
timestamp 1713400504
<< m2contact >>
rect -2 -2 2 2
<< end >>
