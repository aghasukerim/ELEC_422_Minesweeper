magic
tech scmos
timestamp 1713647636
<< metal1 >>
rect 1117 6494 1194 6529
rect 1421 6498 1485 6528
rect 1715 6489 1783 6528
rect 2019 6493 2084 6530
rect 2319 6498 2392 6528
rect 2619 6491 2690 6528
rect 3219 6495 3293 6528
rect 3511 6503 3597 6530
rect 3809 6497 3894 6528
rect 4114 6502 4185 6532
rect 4414 6497 4489 6534
rect 4720 6496 4777 6523
rect 5315 6497 5389 6528
rect 5619 6495 5691 6532
rect 1025 5767 1029 5777
rect 1111 5767 1115 5791
rect 1025 5763 1115 5767
rect 1325 5767 1329 5777
rect 1411 5767 1415 5791
rect 1325 5763 1415 5767
rect 1625 5767 1629 5777
rect 1711 5767 1715 5790
rect 1625 5763 1715 5767
rect 1925 5767 1929 5777
rect 2011 5767 2015 5791
rect 1925 5763 2015 5767
rect 2225 5767 2229 5777
rect 2311 5767 2315 5790
rect 2225 5763 2315 5767
rect 2525 5767 2529 5777
rect 2611 5767 2615 5794
rect 2525 5763 2615 5767
rect 3125 5767 3129 5777
rect 3211 5767 3215 5790
rect 3125 5763 3215 5767
rect 3425 5767 3429 5777
rect 3511 5767 3515 5790
rect 3425 5763 3515 5767
rect 3725 5767 3729 5777
rect 3811 5767 3815 5789
rect 3725 5763 3815 5767
rect 4025 5767 4029 5777
rect 4111 5767 4115 5791
rect 4025 5763 4115 5767
rect 4325 5767 4329 5777
rect 4411 5767 4415 5790
rect 4325 5763 4415 5767
rect 4625 5767 4629 5777
rect 4711 5767 4715 5790
rect 4625 5763 4715 5767
rect 5225 5767 5229 5777
rect 5311 5767 5315 5792
rect 5225 5763 5315 5767
rect 5525 5767 5529 5777
rect 5611 5767 5615 5792
rect 5525 5763 5615 5767
rect 273 5624 311 5676
rect 5762 5611 5789 5615
rect 5762 5528 5766 5611
rect 6507 5598 6533 5696
rect 5762 5524 5777 5528
rect 266 5317 310 5377
rect 1008 5311 1042 5315
rect 1038 5228 1042 5311
rect 1023 5224 1042 5228
rect 5762 5311 5790 5315
rect 5762 5228 5766 5311
rect 6502 5308 6531 5392
rect 5762 5224 5777 5228
rect 271 5010 304 5087
rect 6501 5018 6535 5098
rect 1019 5011 1042 5015
rect 1038 4928 1042 5011
rect 1023 4924 1042 4928
rect 5762 5011 5789 5015
rect 5762 4928 5766 5011
rect 5762 4924 5777 4928
rect 268 4713 303 4781
rect 1019 4711 1042 4715
rect 1038 4628 1042 4711
rect 1023 4624 1042 4628
rect 5762 4711 5788 4715
rect 6501 4714 6532 4801
rect 5762 4628 5766 4711
rect 5762 4624 5777 4628
rect 6502 4408 6534 4486
rect 1023 4272 1028 4276
rect 1024 4189 1028 4272
rect 1008 4185 1028 4189
rect 267 4116 311 4179
rect 268 3812 309 3881
rect 1008 3811 1040 3815
rect 1036 3728 1040 3811
rect 1023 3724 1040 3728
rect 5762 3811 5792 3815
rect 5762 3728 5766 3811
rect 6508 3795 6534 3889
rect 5762 3724 5777 3728
rect 267 3505 301 3584
rect 6505 3580 6533 3592
rect 6502 3517 6533 3580
rect 1009 3511 1040 3515
rect 1036 3428 1040 3511
rect 1023 3424 1040 3428
rect 5748 3511 5792 3515
rect 5748 3429 5752 3511
rect 6505 3496 6533 3517
rect 5748 3425 5777 3429
rect 267 3211 302 3280
rect 1010 3211 1040 3215
rect 1036 3128 1040 3211
rect 1023 3124 1040 3128
rect 5751 3211 5792 3215
rect 6502 3214 6532 3288
rect 5751 3128 5755 3211
rect 5751 3124 5777 3128
rect 262 2913 302 2983
rect 5741 2911 5792 2915
rect 5741 2828 5745 2911
rect 6506 2904 6532 3002
rect 5741 2824 5778 2828
rect 273 2615 316 2677
rect 1007 2646 1054 2652
rect 1048 2605 1054 2646
rect 6498 2616 6535 2692
rect 5752 2611 5792 2615
rect 1048 2599 1965 2605
rect 5752 2528 5756 2611
rect 5752 2524 5777 2528
rect 2457 1973 2463 2054
rect 2343 1967 2463 1973
rect 2343 1011 2349 1967
rect 4063 1957 4069 2057
rect 6504 2017 6535 2095
rect 5772 2011 5792 2015
rect 4063 1951 4149 1957
rect 4143 1015 4149 1951
rect 5772 1928 5776 2011
rect 5772 1924 5777 1928
rect 5770 1711 5792 1715
rect 5770 1629 5774 1711
rect 6504 1710 6533 1798
rect 5770 1625 5777 1629
rect 5756 1411 5792 1415
rect 6502 1414 6533 1490
rect 5756 1329 5760 1411
rect 5756 1325 5778 1329
rect 6501 1118 6535 1190
rect 5773 1111 5792 1115
rect 5524 1033 5615 1037
rect 5224 1025 5315 1029
rect 5311 1008 5315 1025
rect 5524 1022 5528 1033
rect 5611 1008 5615 1033
rect 5773 1029 5777 1111
rect 1112 272 1177 303
rect 1412 269 1479 307
rect 1715 267 1787 308
rect 2022 273 2078 312
rect 2310 271 2382 310
rect 2612 268 2682 313
rect 2915 270 2980 308
rect 3214 272 3285 302
rect 3514 271 3582 306
rect 3817 272 3883 304
rect 4112 270 4186 314
rect 4417 270 4484 304
rect 4713 264 4791 304
rect 5013 267 5088 307
rect 5318 267 5392 303
rect 5610 265 5688 303
<< m2contact >>
rect 1025 5777 1029 5781
rect 1325 5777 1329 5781
rect 1625 5777 1629 5781
rect 1925 5777 1929 5781
rect 2225 5777 2229 5781
rect 2525 5777 2529 5781
rect 3125 5777 3129 5781
rect 3425 5777 3429 5781
rect 3725 5777 3729 5781
rect 4025 5777 4029 5781
rect 4325 5777 4329 5781
rect 4625 5777 4629 5781
rect 5225 5777 5229 5781
rect 5525 5777 5529 5781
rect 5777 5524 5781 5528
rect 1019 5224 1023 5228
rect 5777 5224 5781 5228
rect 1019 4924 1023 4928
rect 5777 4924 5781 4928
rect 1019 4624 1023 4628
rect 5777 4624 5781 4628
rect 1019 4272 1023 4276
rect 1019 3724 1023 3728
rect 5777 3724 5781 3728
rect 1019 3424 1023 3428
rect 5777 3425 5781 3429
rect 1019 3124 1023 3128
rect 5777 3124 5781 3128
rect 5778 2824 5782 2828
rect 5777 2524 5781 2528
rect 5777 1924 5781 1928
rect 5777 1625 5781 1629
rect 5778 1325 5782 1329
rect 5224 1021 5228 1025
rect 5524 1018 5528 1022
rect 5773 1025 5777 1029
<< metal2 >>
rect 1019 5756 1024 5760
rect 1008 5595 1033 5599
rect 1029 5529 1033 5595
rect 1047 5550 1050 5781
rect 1347 5559 1350 5781
rect 1647 5568 1650 5781
rect 1947 5579 1950 5781
rect 2247 5588 2250 5781
rect 2547 5599 2550 5781
rect 3147 5610 3150 5781
rect 3447 5623 3450 5781
rect 3747 5756 3750 5781
rect 4047 5756 4050 5781
rect 4347 5756 4350 5781
rect 4647 5756 4650 5781
rect 5247 5756 5250 5781
rect 5547 5756 5550 5783
rect 3447 5620 4770 5623
rect 3147 5607 4546 5610
rect 2547 5596 4490 5599
rect 2247 5585 3922 5588
rect 1947 5576 3874 5579
rect 1647 5565 3778 5568
rect 1347 5556 3706 5559
rect 1047 5547 3546 5550
rect 1015 5525 1033 5529
rect 1019 5247 3522 5250
rect 1063 5238 3394 5241
rect 1063 4950 1066 5238
rect 1019 4947 1066 4950
rect 1083 5229 3314 5232
rect 1083 4650 1086 5229
rect 1019 4647 1086 4650
rect 1101 5222 3234 5225
rect 1101 4253 1104 5222
rect 1017 4250 1104 4253
rect 1121 5214 3090 5217
rect 1010 3751 1051 3753
rect 1121 3751 1124 5214
rect 1010 3748 1124 3751
rect 1135 5205 3074 5208
rect 1010 3744 1051 3748
rect 1019 3452 1051 3453
rect 1135 3452 1138 5205
rect 1019 3449 1138 3452
rect 1153 5198 3058 5201
rect 1019 3444 1051 3449
rect 1019 3151 1051 3153
rect 1153 3151 1156 5198
rect 3055 5064 3058 5198
rect 3071 5064 3074 5205
rect 3087 5063 3090 5214
rect 3231 5065 3234 5222
rect 3311 5064 3314 5229
rect 3391 5064 3394 5238
rect 3519 5064 3522 5247
rect 3543 5063 3546 5547
rect 3703 5063 3706 5556
rect 3775 5065 3778 5565
rect 3871 5062 3874 5576
rect 3919 5064 3922 5585
rect 4487 5064 4490 5596
rect 4543 5063 4546 5607
rect 4767 5063 4770 5620
rect 5774 5546 5781 5551
rect 5774 5246 5781 5251
rect 5774 4946 5781 4951
rect 5774 4646 5781 4651
rect 5762 4395 5792 4399
rect 5762 4328 5766 4395
rect 5762 4324 5783 4328
rect 5774 3746 5781 3751
rect 5781 3660 5785 3665
rect 5782 3495 5792 3499
rect 5763 3446 5781 3450
rect 5781 3424 5785 3428
rect 1019 3148 1156 3151
rect 1019 3144 1051 3148
rect 5763 3146 5781 3150
rect 1019 3060 1024 3064
rect 1008 2895 1035 2899
rect 1031 2828 1035 2895
rect 5763 2847 5781 2851
rect 1017 2824 1035 2828
rect 5763 2546 5781 2550
rect 2175 1985 2178 2038
rect 1260 1982 2178 1985
rect 1025 1024 1099 1028
rect 1025 1017 1029 1024
rect 1095 1008 1099 1024
rect 1260 1019 1263 1982
rect 2247 1969 2250 2038
rect 1560 1966 2250 1969
rect 1324 1029 1399 1033
rect 1324 1016 1328 1029
rect 1395 1008 1399 1029
rect 1560 1018 1563 1966
rect 2367 1956 2370 2038
rect 3503 2022 3506 2038
rect 1860 1953 2370 1956
rect 2431 2019 3506 2022
rect 1623 1029 1699 1033
rect 1623 1016 1627 1029
rect 1695 1008 1699 1029
rect 1860 1018 1863 1953
rect 2431 1926 2434 2019
rect 3647 2008 3650 2038
rect 2160 1923 2434 1926
rect 2760 2005 3650 2008
rect 1924 1032 1999 1036
rect 1924 1015 1928 1032
rect 1995 1008 1999 1032
rect 2160 1019 2163 1923
rect 2524 1028 2599 1032
rect 2524 1017 2528 1028
rect 2595 1008 2599 1028
rect 2760 1019 2763 2005
rect 3679 1996 3682 2038
rect 3060 1993 3682 1996
rect 2825 1028 2899 1032
rect 2825 1018 2829 1028
rect 2895 1008 2899 1028
rect 3060 1019 3063 1993
rect 3719 1969 3722 2038
rect 3360 1966 3722 1969
rect 3124 1030 3199 1034
rect 3124 1016 3128 1030
rect 3195 1008 3199 1030
rect 3360 1019 3363 1966
rect 3751 1941 3754 2037
rect 3660 1938 3754 1941
rect 3424 1028 3499 1032
rect 3424 1014 3428 1028
rect 3495 1008 3499 1028
rect 3660 1019 3663 1938
rect 3799 1838 3802 2038
rect 4775 1875 4778 2037
rect 5763 1946 5781 1950
rect 4560 1872 4778 1875
rect 3799 1835 3963 1838
rect 3724 1029 3799 1033
rect 3724 1018 3728 1029
rect 3795 1008 3799 1029
rect 3960 1019 3963 1835
rect 4324 1031 4399 1035
rect 4324 1015 4328 1031
rect 4395 1008 4399 1031
rect 4560 1019 4563 1872
rect 5763 1650 5781 1651
rect 5763 1647 5783 1650
rect 5781 1646 5783 1647
rect 5771 1347 5785 1351
rect 5766 1047 5782 1051
rect 4925 1031 4999 1035
rect 4625 1027 4699 1031
rect 4625 1015 4629 1027
rect 4695 1008 4699 1027
rect 4860 1019 4864 1023
rect 4925 1016 4929 1031
rect 4995 1008 4999 1031
rect 5160 1018 5164 1024
rect 5224 1019 5228 1021
rect 5247 1019 5250 1039
rect 5547 1019 5550 1047
rect 5777 1025 5784 1029
<< m3contact >>
rect 1024 5756 1028 5760
rect 3747 5752 3751 5756
rect 4047 5752 4051 5756
rect 4347 5752 4351 5756
rect 4647 5752 4651 5756
rect 5247 5752 5251 5756
rect 5547 5752 5551 5756
rect 5770 5547 5774 5551
rect 5770 5247 5774 5251
rect 5770 4947 5774 4951
rect 5770 4647 5774 4651
rect 5776 4560 5781 4565
rect 5770 3747 5774 3751
rect 5759 3446 5763 3450
rect 5759 3146 5763 3150
rect 1024 3060 1028 3064
rect 5759 2847 5763 2851
rect 5759 2546 5763 2550
rect 5759 1946 5763 1950
rect 5759 1647 5763 1651
rect 5767 1347 5771 1351
rect 5547 1047 5551 1051
rect 5762 1047 5766 1051
rect 5247 1039 5251 1043
rect 4860 1023 4864 1027
rect 5160 1024 5164 1028
<< metal3 >>
rect 1023 5760 1029 5761
rect 1023 5756 1024 5760
rect 1028 5757 1032 5760
rect 1028 5756 1033 5757
rect 3746 5756 3752 5757
rect 4046 5756 4052 5757
rect 1023 5755 1185 5756
rect 1027 5751 1185 5755
rect 3745 5752 3747 5756
rect 3751 5752 3753 5756
rect 4046 5753 4047 5756
rect 3745 5751 3753 5752
rect 4045 5752 4047 5753
rect 4051 5753 4052 5756
rect 4346 5756 4352 5757
rect 4051 5752 4053 5753
rect 1180 4449 1185 5751
rect 3746 5633 3751 5751
rect 4045 5748 4053 5752
rect 4346 5752 4347 5756
rect 4351 5752 4352 5756
rect 4346 5751 4352 5752
rect 4646 5756 4652 5757
rect 4646 5752 4647 5756
rect 4651 5752 4652 5756
rect 4047 5663 4052 5748
rect 4345 5690 4353 5751
rect 4646 5728 4652 5752
rect 5246 5756 5252 5757
rect 5246 5752 5247 5756
rect 5251 5752 5252 5756
rect 5246 5751 5252 5752
rect 5546 5756 5552 5757
rect 5546 5752 5547 5756
rect 5551 5752 5552 5756
rect 5546 5751 5552 5752
rect 4646 5723 5236 5728
rect 4345 5685 5221 5690
rect 4047 5658 5201 5663
rect 3746 5628 5176 5633
rect 5171 4809 5176 5628
rect 5004 4804 5176 4809
rect 5196 4639 5201 5658
rect 5003 4634 5201 4639
rect 1180 4444 1937 4449
rect 5216 4359 5221 5685
rect 5003 4354 5221 4359
rect 5231 4339 5236 5723
rect 5002 4334 5236 4339
rect 1169 4244 1939 4249
rect 1169 3065 1174 4244
rect 1935 4164 1939 4169
rect 1934 4144 1938 4149
rect 5247 4062 5252 5751
rect 5547 5744 5552 5751
rect 5544 5739 5552 5744
rect 5008 4057 5252 4062
rect 5504 5624 5509 5626
rect 5544 5624 5549 5739
rect 5504 5619 5549 5624
rect 1934 4034 1938 4039
rect 5008 4038 5013 4057
rect 1934 3994 1938 3999
rect 5504 3959 5509 5619
rect 5747 5551 5775 5552
rect 5003 3954 5509 3959
rect 5530 5547 5770 5551
rect 5774 5547 5775 5551
rect 5530 5546 5752 5547
rect 5765 5546 5775 5547
rect 5530 3799 5535 5546
rect 5003 3794 5535 3799
rect 5556 5251 5775 5252
rect 5556 5247 5770 5251
rect 5774 5247 5775 5251
rect 5556 3709 5561 5247
rect 5765 5246 5775 5247
rect 5002 3704 5561 3709
rect 5590 4951 5775 4952
rect 5590 4947 5770 4951
rect 5774 4947 5775 4951
rect 5590 3579 5595 4947
rect 5765 4946 5775 4947
rect 5748 4651 5775 4652
rect 5004 3574 5595 3579
rect 5632 4647 5770 4651
rect 5774 4647 5775 4651
rect 5632 4646 5754 4647
rect 5765 4646 5775 4647
rect 5632 3559 5637 4646
rect 5775 4565 5782 4566
rect 5003 3554 5637 3559
rect 5664 4560 5776 4565
rect 5781 4560 5782 4565
rect 5664 3489 5669 4560
rect 5775 4559 5782 4560
rect 5004 3484 5669 3489
rect 5700 3751 5775 3752
rect 5700 3747 5770 3751
rect 5774 3747 5775 3751
rect 5700 3399 5705 3747
rect 5765 3746 5775 3747
rect 5758 3450 5764 3451
rect 5002 3394 5705 3399
rect 5721 3446 5759 3450
rect 5763 3446 5764 3450
rect 5721 3445 5764 3446
rect 5721 3359 5726 3445
rect 5002 3354 5726 3359
rect 5003 3244 5475 3249
rect 5002 3154 5411 3159
rect 1023 3064 1174 3065
rect 1023 3060 1024 3064
rect 1028 3060 1174 3064
rect 1023 3059 1030 3060
rect 5004 3044 5362 3049
rect 5003 3004 5348 3009
rect 5002 2984 5323 2989
rect 5004 2954 5308 2959
rect 5004 2934 5291 2939
rect 5003 2844 5269 2849
rect 5002 2814 5252 2819
rect 5004 2754 5165 2759
rect 5004 2514 5016 2519
rect 5011 2017 5016 2514
rect 4860 2012 5016 2017
rect 4860 1028 4865 2012
rect 5160 1029 5165 2754
rect 5247 1044 5252 2814
rect 5264 1084 5269 2844
rect 5286 1120 5291 2934
rect 5303 1352 5308 2954
rect 5318 1652 5323 2984
rect 5343 1951 5348 3004
rect 5357 2550 5362 3044
rect 5406 2850 5411 3154
rect 5470 3151 5475 3244
rect 5470 3150 5764 3151
rect 5470 3146 5759 3150
rect 5763 3146 5764 3150
rect 5758 3145 5764 3146
rect 5758 2851 5764 2852
rect 5754 2850 5759 2851
rect 5406 2847 5759 2850
rect 5763 2847 5764 2851
rect 5406 2846 5764 2847
rect 5406 2845 5759 2846
rect 5758 2550 5764 2551
rect 5357 2546 5759 2550
rect 5763 2546 5764 2550
rect 5357 2545 5764 2546
rect 5343 1950 5764 1951
rect 5343 1946 5759 1950
rect 5763 1946 5764 1950
rect 5758 1945 5764 1946
rect 5318 1651 5764 1652
rect 5318 1647 5759 1651
rect 5763 1647 5764 1651
rect 5758 1646 5764 1647
rect 5303 1351 5772 1352
rect 5303 1347 5767 1351
rect 5771 1347 5772 1351
rect 5766 1346 5772 1347
rect 5286 1115 5578 1120
rect 5264 1079 5552 1084
rect 5547 1052 5552 1079
rect 5546 1051 5552 1052
rect 5546 1047 5547 1051
rect 5551 1047 5552 1051
rect 5573 1052 5578 1115
rect 5573 1051 5767 1052
rect 5573 1047 5762 1051
rect 5766 1047 5767 1051
rect 5546 1046 5552 1047
rect 5761 1046 5767 1047
rect 5246 1043 5252 1044
rect 5246 1039 5247 1043
rect 5251 1039 5252 1043
rect 5246 1038 5252 1039
rect 4859 1027 4865 1028
rect 4859 1023 4860 1027
rect 4864 1023 4865 1027
rect 5159 1028 5165 1029
rect 5159 1024 5160 1028
rect 5164 1024 5165 1028
rect 5159 1023 5165 1024
rect 4859 1022 4865 1023
use PadFrame64  PadFrame64_0
timestamp 1713593144
transform 1 0 2500 0 1 2400
box -2500 -2400 4300 4400
use top_module  top_module_0
timestamp 1713592123
transform 1 0 1925 0 1 2032
box 0 0 3088 3040
<< labels >>
rlabel metal1 2310 271 2382 310 0 Vdd!
rlabel metal1 273 2615 316 2677 0 GND!
rlabel space 0 0 6800 6800 1 in_n_mines1unexpand
rlabel metal2 2175 2034 2178 2038 1 in_n_mines1
rlabel metal1 1112 272 1177 303 0 p_in_n_mines1
rlabel metal2 2247 2034 2250 2038 1 in_n_mines0
rlabel metal1 1412 269 1479 307 1 p_in_n_mines0
rlabel metal2 2367 2034 2370 2038 1 in_n_mines2
rlabel metal1 1715 267 1787 308 0 p_in_n_mines2
rlabel metal2 3503 2035 3506 2038 1 in_clkb
rlabel metal1 2022 273 2078 312 0 p_in_clkb
rlabel metal2 3647 2035 3650 2038 1 in_data2
rlabel metal1 2612 268 2682 313 0 p_in_data2
rlabel metal2 3679 2035 3682 2038 1 in_data1
rlabel metal1 2915 270 2980 308 0 p_in_data1
rlabel metal2 3719 2034 3722 2038 1 in_data0
rlabel metal1 3214 272 3285 302 1 p_in_data0
rlabel metal3 5004 3484 5009 3489 1 in_clka
rlabel metal2 3751 2034 3754 2037 1 in_data3
rlabel metal1 3514 271 3582 306 1 p_in_data3
rlabel metal2 3799 2035 3802 2038 1 in_data4
rlabel metal1 3817 272 3883 304 0 p_in_data4
rlabel metal2 4775 2034 4778 2037 1 in_place
rlabel metal1 4417 270 4484 304 0 p_in_place
rlabel metal1 4112 270 4186 314 0 Vdd!
rlabel metal3 5004 2514 5008 2519 1 in_data_in
rlabel metal1 4713 264 4791 304 0 p_in_data_in
rlabel metal3 5004 2754 5009 2759 1 in_restart
rlabel metal1 5013 267 5088 307 0 p_in_restart
rlabel metal3 5003 2814 5007 2819 1 out_global_score6
rlabel metal3 5003 2844 5007 2849 1 out_global_score5
rlabel metal1 5318 267 5392 303 0 p_out_global_score6
rlabel metal1 5610 265 5688 303 1 p_out_global_score5
rlabel metal3 5004 2934 5008 2939 1 out_gameover
rlabel metal1 6501 1118 6535 1190 0 p_out_gameover
rlabel metal3 5005 2954 5009 2959 1 out_n_nearby1
rlabel metal1 6502 1414 6533 1490 0 p_out_n_nearby1
rlabel metal3 5003 2984 5007 2989 1 out_global_score7
rlabel metal3 5004 3004 5008 3009 1 out_n_nearby0
rlabel metal3 5005 3044 5009 3049 1 out_global_score4
rlabel metal1 6504 1710 6533 1798 0 p_out_global_score7
rlabel metal1 6504 2017 6535 2095 0 p_out_n_nearby0
rlabel metal1 6498 2616 6535 2692 0 p_out_global_score4
rlabel metal3 5003 3154 5008 3159 1 out_global_score3
rlabel metal1 6506 2904 6532 3002 0 p_out_global_score3
rlabel metal3 5003 3244 5008 3249 1 out_global_score2
rlabel metal1 6502 3214 6532 3288 1 p_out_global_score2
rlabel metal3 5003 3354 5007 3359 1 out_global_score1
rlabel metal1 6505 3496 6533 3592 0 p_out_global_score1
rlabel metal3 5002 3394 5008 3399 1 out_win
rlabel metal1 6508 3795 6534 3889 0 p_out_win
rlabel metal1 6502 4408 6534 4486 0 p_in_clka
rlabel metal3 5003 3554 5008 3559 1 out_temp_cleared4
rlabel metal1 6501 4714 6532 4801 0 p_out_temp_cleared4
rlabel metal3 5004 3574 5008 3579 1 out_temp_cleared3
rlabel metal1 6501 5018 6535 5098 0 p_out_temp_cleared3
rlabel metal3 5003 3704 5007 3709 1 out_temp_cleared0
rlabel metal1 6502 5308 6531 5392 0 p_out_temp_cleared0
rlabel metal3 5003 3794 5008 3799 1 out_temp_cleared1
rlabel metal1 6507 5598 6533 5696 0 p_out_temp_cleared1
rlabel metal3 5003 3954 5009 3959 1 out_temp_cleared24
rlabel metal3 5008 4038 5013 4043 1 out_temp_cleared5
rlabel metal3 5002 4334 5007 4339 1 out_temp_cleared2
rlabel metal1 5619 6495 5691 6532 1 p_out_temp_cleared24
rlabel metal1 5315 6497 5389 6528 1 p_out_temp_cleared5
rlabel metal1 4720 6496 4777 6523 1 p_out_temp_cleared2
rlabel metal3 5003 4354 5007 4359 1 out_temp_cleared6
rlabel metal1 4414 6497 4489 6534 0 p_out_temp_cleared6
rlabel metal3 5003 4634 5007 4639 1 out_temp_cleared7
rlabel metal1 4114 6502 4185 6532 0 p_out_temp_cleared7
rlabel metal3 5004 4804 5009 4809 1 out_temp_cleared8
rlabel metal1 3809 6497 3894 6528 0 p_out_temp_cleared8
rlabel metal2 4767 5063 4770 5067 1 out_temp_cleared9
rlabel metal1 3511 6503 3597 6530 0 p_out_temp_cleared9
rlabel metal2 4543 5063 4546 5066 1 out_temp_cleared10
rlabel metal1 3219 6495 3293 6528 0 p_out_temp_cleared10
rlabel metal2 4487 5064 4490 5067 1 out_temp_cleared11
rlabel metal1 2619 6491 2690 6528 0 p_out_temp_cleared11
rlabel metal2 3919 5064 3922 5067 1 out_temp_cleared12
rlabel metal1 2319 6498 2392 6528 0 p_out_temp_cleared12
rlabel metal2 3871 5062 3874 5066 1 out_temp_cleared23
rlabel metal1 2019 6493 2084 6530 0 p_out_temp_cleared23
rlabel metal2 3775 5065 3778 5068 1 out_temp_cleared13
rlabel metal1 1715 6489 1783 6528 0 p_out_temp_cleared13
rlabel metal2 3703 5063 3706 5066 1 out_temp_cleared14
rlabel metal1 1421 6498 1485 6528 0 p_out_temp_cleared14
rlabel metal2 3543 5063 3546 5067 1 out_temp_cleared22
rlabel metal1 1117 6494 1194 6529 0 p_out_temp_cleared22
rlabel metal2 3519 5064 3522 5067 1 out_temp_cleared20
rlabel metal1 266 5317 310 5377 0 p_out_temp_cleared20
rlabel metal2 3391 5064 3394 5067 1 out_temp_cleared21
rlabel metal1 271 5010 304 5087 0 p_out_temp_cleared21
rlabel metal2 3311 5065 3314 5068 1 out_temp_cleared19
rlabel metal1 268 4713 303 4781 0 p_out_temp_cleared19
rlabel metal2 3231 5066 3234 5068 1 out_temp_cleared18
rlabel metal1 267 4116 311 4179 0 p_out_temp_cleared18
rlabel metal2 3087 5063 3090 5066 1 out_temp_cleared15
rlabel metal1 268 3812 309 3881 0 p_out_temp_cleared15
rlabel metal2 3071 5064 3074 5067 1 out_temp_cleared17
rlabel metal2 3055 5064 3058 5067 1 out_temp_cleared16
rlabel metal1 267 3505 301 3584 0 p_out_temp_cleared17
rlabel metal1 267 3211 302 3280 0 p_out_temp_cleared16
rlabel metal3 1933 4444 1937 4449 1 in_incr2
rlabel metal3 1935 4244 1939 4249 1 in_incr1
rlabel metal3 1935 4164 1939 4169 1 in_mult2
rlabel metal3 1934 4144 1938 4149 1 in_mult1
rlabel metal3 1934 4034 1938 4039 1 in_mult0
rlabel metal3 1934 3994 1938 3999 1 in_incr0
rlabel metal1 273 5624 311 5676 0 p_in_incr2
rlabel metal1 262 2913 302 2983 0 p_in_incr1
<< end >>
