magic
tech scmos
timestamp 1713592123
<< m2contact >>
rect -2 -2 2 2
<< end >>
