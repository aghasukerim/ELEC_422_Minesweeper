magic
tech scmos
timestamp 1713400504
<< metal1 >>
rect 14 3007 3074 3027
rect 38 2983 3050 3003
rect 38 2967 3050 2973
rect 290 2933 324 2936
rect 394 2933 436 2936
rect 554 2933 572 2936
rect 658 2933 684 2936
rect 826 2933 844 2936
rect 914 2933 940 2936
rect 1162 2933 1172 2936
rect 1258 2933 1292 2936
rect 1314 2933 1332 2936
rect 1364 2933 1381 2936
rect 1162 2926 1165 2933
rect 1378 2926 1381 2933
rect 1754 2926 1757 2935
rect 1946 2926 1949 2935
rect 2706 2926 2709 2935
rect 2722 2933 2748 2936
rect 178 2923 204 2926
rect 284 2923 325 2926
rect 458 2923 500 2926
rect 506 2923 516 2926
rect 580 2923 613 2926
rect 658 2923 692 2926
rect 818 2923 852 2926
rect 1004 2923 1029 2926
rect 1100 2923 1125 2926
rect 1156 2923 1165 2926
rect 1180 2923 1228 2926
rect 1300 2923 1340 2926
rect 1378 2923 1420 2926
rect 1468 2923 1485 2926
rect 1530 2923 1540 2926
rect 1588 2923 1613 2926
rect 1684 2923 1709 2926
rect 1740 2923 1757 2926
rect 1764 2923 1796 2926
rect 1876 2923 1901 2926
rect 1932 2923 1949 2926
rect 1956 2923 1996 2926
rect 2076 2923 2101 2926
rect 2138 2923 2164 2926
rect 2348 2923 2365 2926
rect 2434 2923 2444 2926
rect 2628 2923 2653 2926
rect 2684 2923 2709 2926
rect 2716 2923 2756 2926
rect 348 2913 357 2916
rect 708 2913 717 2916
rect 868 2913 877 2916
rect 14 2867 3074 2873
rect 1162 2833 1196 2836
rect 2426 2833 2444 2836
rect 2634 2833 2652 2836
rect 1162 2816 1165 2833
rect 1204 2823 1261 2826
rect 1356 2823 1365 2826
rect 2132 2823 2141 2826
rect 2156 2823 2173 2826
rect 2252 2823 2261 2826
rect 2428 2823 2437 2826
rect 2452 2823 2493 2826
rect 2636 2823 2645 2826
rect 116 2813 149 2816
rect 218 2813 252 2816
rect 258 2813 284 2816
rect 418 2813 452 2816
rect 466 2813 484 2816
rect 522 2813 572 2816
rect 700 2813 717 2816
rect 722 2813 748 2816
rect 754 2813 788 2816
rect 820 2813 837 2816
rect 842 2813 876 2816
rect 882 2813 908 2816
rect 940 2813 949 2816
rect 962 2813 1012 2816
rect 1124 2813 1165 2816
rect 1266 2813 1276 2816
rect 1290 2813 1348 2816
rect 1458 2813 1500 2816
rect 1572 2813 1597 2816
rect 1706 2806 1709 2814
rect 1780 2813 1789 2816
rect 1922 2813 1940 2816
rect 1956 2813 1981 2816
rect 2020 2813 2045 2816
rect 2108 2813 2125 2816
rect 2178 2813 2229 2816
rect 2314 2813 2340 2816
rect 2370 2813 2436 2816
rect 2514 2813 2540 2816
rect 2666 2813 2716 2816
rect 2746 2813 2796 2816
rect 122 2803 148 2806
rect 322 2803 348 2806
rect 1098 2803 1116 2806
rect 1210 2803 1268 2806
rect 1292 2803 1309 2806
rect 1354 2803 1420 2806
rect 1450 2803 1492 2806
rect 1674 2803 1684 2806
rect 1706 2803 1772 2806
rect 1850 2803 1876 2806
rect 1890 2803 1932 2806
rect 2090 2803 2100 2806
rect 2226 2805 2229 2813
rect 2266 2803 2292 2806
rect 2306 2803 2332 2806
rect 2356 2803 2365 2806
rect 2458 2803 2500 2806
rect 38 2767 3050 2773
rect 570 2743 588 2746
rect 714 2736 717 2745
rect 1722 2736 1725 2756
rect 2146 2743 2156 2746
rect 2594 2743 2620 2746
rect 138 2733 148 2736
rect 338 2733 356 2736
rect 404 2733 412 2736
rect 506 2733 516 2736
rect 578 2733 613 2736
rect 708 2733 717 2736
rect 724 2733 757 2736
rect 842 2733 860 2736
rect 940 2733 956 2736
rect 1066 2733 1100 2736
rect 1116 2733 1133 2736
rect 1162 2733 1180 2736
rect 1204 2733 1237 2736
rect 1316 2733 1341 2736
rect 1394 2733 1412 2736
rect 1490 2733 1516 2736
rect 1546 2733 1580 2736
rect 1604 2733 1613 2736
rect 1674 2733 1692 2736
rect 890 2726 893 2733
rect 116 2723 149 2726
rect 218 2723 236 2726
rect 242 2723 268 2726
rect 306 2723 332 2726
rect 500 2723 517 2726
rect 610 2723 628 2726
rect 692 2723 717 2726
rect 796 2723 821 2726
rect 868 2723 893 2726
rect 916 2723 949 2726
rect 978 2723 1004 2726
rect 1036 2723 1045 2726
rect 1058 2723 1092 2726
rect 1124 2723 1149 2726
rect 1178 2723 1188 2726
rect 172 2713 181 2716
rect 876 2713 885 2716
rect 1204 2713 1237 2716
rect 1234 2706 1237 2713
rect 1338 2706 1341 2733
rect 1450 2726 1468 2727
rect 1706 2726 1709 2736
rect 1722 2733 1756 2736
rect 1772 2733 1837 2736
rect 1866 2733 1885 2736
rect 1890 2733 1932 2736
rect 1948 2733 1957 2736
rect 2082 2733 2108 2736
rect 2164 2733 2197 2736
rect 2298 2733 2308 2736
rect 2404 2733 2453 2736
rect 2514 2733 2540 2736
rect 2628 2733 2645 2736
rect 1394 2724 1468 2726
rect 1394 2723 1453 2724
rect 1538 2723 1588 2726
rect 1602 2723 1652 2726
rect 1700 2723 1709 2726
rect 1780 2723 1813 2726
rect 1826 2723 1836 2726
rect 1866 2725 1869 2733
rect 2834 2726 2837 2735
rect 2858 2733 2884 2736
rect 2916 2733 2933 2736
rect 1874 2723 1924 2726
rect 2020 2723 2045 2726
rect 2082 2723 2116 2726
rect 2418 2723 2468 2726
rect 2636 2723 2653 2726
rect 2804 2723 2837 2726
rect 2850 2723 2892 2726
rect 2922 2723 2988 2726
rect 1388 2713 1397 2716
rect 1484 2713 1509 2716
rect 1540 2713 1573 2716
rect 1604 2713 1621 2716
rect 2484 2713 2493 2716
rect 1234 2703 1253 2706
rect 1338 2703 1380 2706
rect 1442 2703 1476 2706
rect 14 2667 3074 2673
rect 1730 2633 1748 2636
rect 170 2623 189 2626
rect 186 2616 189 2623
rect 92 2613 101 2616
rect 148 2613 181 2616
rect 186 2613 196 2616
rect 276 2613 309 2616
rect 418 2613 428 2616
rect 466 2613 476 2616
rect 508 2613 548 2616
rect 596 2613 605 2616
rect 708 2613 733 2616
rect 772 2613 797 2616
rect 826 2613 853 2616
rect 884 2613 909 2616
rect 98 2603 116 2606
rect 164 2603 188 2606
rect 282 2603 308 2606
rect 356 2603 389 2606
rect 652 2603 661 2606
rect 738 2603 748 2606
rect 794 2605 797 2613
rect 850 2606 853 2613
rect 850 2603 860 2606
rect 906 2603 909 2613
rect 914 2606 917 2626
rect 1596 2623 1605 2626
rect 1722 2623 1732 2626
rect 1756 2623 1781 2626
rect 2076 2623 2085 2626
rect 2212 2623 2253 2626
rect 2756 2623 2765 2626
rect 2780 2623 2821 2626
rect 1778 2616 1781 2623
rect 940 2613 965 2616
rect 988 2613 997 2616
rect 1028 2613 1045 2616
rect 1092 2613 1109 2616
rect 1148 2613 1173 2616
rect 1180 2613 1228 2616
rect 1324 2613 1349 2616
rect 1394 2613 1412 2616
rect 1492 2613 1517 2616
rect 1554 2613 1580 2616
rect 1778 2613 1789 2616
rect 1842 2613 1852 2616
rect 1858 2613 1884 2616
rect 1898 2613 1932 2616
rect 1954 2613 1980 2616
rect 1994 2613 2005 2616
rect 2034 2613 2060 2616
rect 2116 2613 2133 2616
rect 2172 2613 2181 2616
rect 2204 2613 2245 2616
rect 2260 2613 2301 2616
rect 2308 2613 2349 2616
rect 914 2603 932 2606
rect 938 2603 980 2606
rect 994 2605 997 2613
rect 1044 2603 1053 2606
rect 1170 2605 1173 2613
rect 2002 2606 2005 2613
rect 2394 2606 2397 2616
rect 2492 2613 2533 2616
rect 2564 2613 2597 2616
rect 2666 2613 2708 2616
rect 2786 2613 2836 2616
rect 2866 2613 2900 2616
rect 2956 2613 2965 2616
rect 3012 2613 3021 2616
rect 1394 2603 1404 2606
rect 1428 2603 1453 2606
rect 1554 2603 1572 2606
rect 1796 2603 1829 2606
rect 1834 2603 1844 2606
rect 1946 2603 1972 2606
rect 2002 2603 2052 2606
rect 2146 2603 2164 2606
rect 2178 2603 2196 2606
rect 2226 2603 2252 2606
rect 2380 2603 2397 2606
rect 362 2593 388 2596
rect 1762 2593 1788 2596
rect 2530 2595 2533 2613
rect 2724 2603 2749 2606
rect 2794 2603 2828 2606
rect 2866 2603 2869 2613
rect 38 2567 3050 2573
rect 162 2543 196 2546
rect 1450 2543 1477 2546
rect 1930 2543 1948 2546
rect 2090 2543 2108 2546
rect 2154 2543 2164 2546
rect 1474 2536 1477 2543
rect 2178 2536 2181 2546
rect 2194 2543 2220 2546
rect 2234 2543 2268 2546
rect 2514 2543 2540 2546
rect 2554 2543 2604 2546
rect 178 2526 181 2536
rect 186 2533 204 2536
rect 346 2533 380 2536
rect 426 2533 436 2536
rect 490 2533 508 2536
rect 626 2533 644 2536
rect 674 2533 708 2536
rect 820 2533 845 2536
rect 906 2533 916 2536
rect 1028 2533 1061 2536
rect 1066 2533 1092 2536
rect 1124 2533 1141 2536
rect 1266 2533 1284 2536
rect 1394 2533 1412 2536
rect 1444 2533 1469 2536
rect 1474 2533 1484 2536
rect 1602 2533 1628 2536
rect 1714 2533 1732 2536
rect 1764 2533 1805 2536
rect 1946 2533 1956 2536
rect 1970 2533 2012 2536
rect 2172 2533 2181 2536
rect 490 2526 493 2533
rect 570 2526 573 2533
rect 626 2526 629 2533
rect 1466 2526 1469 2533
rect 74 2523 100 2526
rect 132 2523 181 2526
rect 218 2523 252 2526
rect 258 2523 308 2526
rect 340 2523 388 2526
rect 466 2523 493 2526
rect 532 2523 573 2526
rect 602 2523 629 2526
rect 668 2523 685 2526
rect 706 2523 716 2526
rect 876 2523 917 2526
rect 962 2523 1004 2526
rect 1034 2523 1100 2526
rect 1196 2523 1221 2526
rect 1258 2523 1292 2526
rect 1364 2523 1420 2526
rect 1466 2523 1501 2526
rect 1540 2523 1565 2526
rect 1676 2523 1740 2526
rect 1802 2523 1805 2533
rect 1810 2523 1828 2526
rect 1866 2523 1916 2526
rect 1964 2523 2005 2526
rect 2068 2523 2085 2526
rect 2234 2525 2237 2543
rect 2276 2533 2293 2536
rect 2298 2533 2324 2536
rect 2338 2533 2372 2536
rect 2538 2533 2548 2536
rect 2594 2533 2612 2536
rect 2290 2526 2293 2533
rect 2290 2523 2325 2526
rect 2332 2523 2373 2526
rect 2380 2523 2421 2526
rect 2516 2523 2525 2526
rect 2538 2523 2541 2533
rect 2620 2523 2653 2526
rect 2658 2523 2661 2535
rect 2684 2533 2717 2536
rect 2818 2533 2852 2536
rect 2882 2533 2948 2536
rect 2980 2533 2989 2536
rect 1652 2513 1661 2516
rect 1836 2513 1845 2516
rect 1860 2513 1893 2516
rect 2076 2513 2101 2516
rect 2340 2513 2373 2516
rect 2394 2513 2428 2516
rect 2818 2513 2821 2533
rect 2898 2523 2956 2526
rect 2884 2513 2893 2516
rect 2434 2503 2444 2506
rect 14 2467 3074 2473
rect 1210 2433 1276 2436
rect 2514 2433 2533 2436
rect 2578 2433 2612 2436
rect 2626 2433 2669 2436
rect 884 2423 949 2426
rect 1234 2423 1260 2426
rect 1284 2423 1349 2426
rect 1844 2423 1869 2426
rect 2090 2423 2108 2426
rect 1234 2416 1237 2423
rect 2514 2416 2517 2433
rect 74 2413 140 2416
rect 172 2413 221 2416
rect 274 2413 324 2416
rect 914 2413 964 2416
rect 1010 2413 1076 2416
rect 1180 2413 1189 2416
rect 1196 2413 1237 2416
rect 1338 2413 1356 2416
rect 1388 2413 1445 2416
rect 1626 2413 1668 2416
rect 1732 2413 1757 2416
rect 1900 2413 1933 2416
rect 2012 2413 2045 2416
rect 2204 2413 2245 2416
rect 2316 2413 2341 2416
rect 2372 2413 2413 2416
rect 2492 2413 2517 2416
rect 2530 2415 2533 2433
rect 2620 2423 2653 2426
rect 2666 2415 2669 2433
rect 2954 2433 2973 2436
rect 2954 2426 2957 2433
rect 2908 2423 2957 2426
rect 2690 2413 2748 2416
rect 2780 2413 2829 2416
rect 2874 2413 2892 2416
rect 178 2403 220 2406
rect 644 2403 677 2406
rect 884 2403 893 2406
rect 938 2403 956 2406
rect 994 2403 1068 2406
rect 1092 2403 1157 2406
rect 1290 2403 1364 2406
rect 1380 2403 1421 2406
rect 1506 2403 1548 2406
rect 1554 2403 1604 2406
rect 1628 2403 1653 2406
rect 1802 2403 1820 2406
rect 1850 2403 1892 2406
rect 1906 2403 1948 2406
rect 1970 2403 2004 2406
rect 2138 2403 2196 2406
rect 2252 2403 2301 2406
rect 2314 2403 2364 2406
rect 2474 2403 2484 2406
rect 2754 2403 2772 2406
rect 2802 2403 2828 2406
rect 2858 2403 2884 2406
rect 1922 2393 1940 2396
rect 1962 2393 1996 2396
rect 2010 2393 2052 2396
rect 2170 2393 2188 2396
rect 2226 2393 2244 2396
rect 2266 2393 2300 2396
rect 2410 2393 2428 2396
rect 38 2367 3050 2373
rect 1244 2343 1261 2346
rect 1874 2343 1892 2346
rect 1922 2343 1964 2346
rect 66 2333 108 2336
rect 218 2333 268 2336
rect 324 2333 372 2336
rect 484 2333 509 2336
rect 658 2333 676 2336
rect 690 2333 724 2336
rect 884 2333 925 2336
rect 930 2333 940 2336
rect 90 2323 116 2326
rect 122 2323 132 2326
rect 154 2323 180 2326
rect 212 2323 276 2326
rect 332 2323 357 2326
rect 684 2323 717 2326
rect 748 2313 757 2316
rect 978 2313 981 2336
rect 1044 2333 1117 2336
rect 1146 2326 1149 2335
rect 1154 2333 1228 2336
rect 1242 2333 1316 2336
rect 1364 2333 1413 2336
rect 1418 2333 1444 2336
rect 1858 2333 1900 2336
rect 1972 2333 2020 2336
rect 2170 2333 2196 2336
rect 2244 2333 2293 2336
rect 2330 2333 2356 2336
rect 2564 2333 2581 2336
rect 2762 2333 2796 2336
rect 2834 2326 2837 2336
rect 1002 2323 1020 2326
rect 1106 2323 1132 2326
rect 1146 2323 1220 2326
rect 1250 2323 1341 2326
rect 1372 2323 1436 2326
rect 1468 2323 1525 2326
rect 1148 2313 1157 2316
rect 1482 2313 1532 2316
rect 1538 2306 1541 2325
rect 1636 2323 1661 2326
rect 1740 2323 1765 2326
rect 1796 2323 1805 2326
rect 1852 2323 1869 2326
rect 1908 2323 1925 2326
rect 2028 2323 2069 2326
rect 2108 2323 2117 2326
rect 2204 2323 2221 2326
rect 2324 2323 2349 2326
rect 2578 2323 2628 2326
rect 2634 2323 2652 2326
rect 2698 2323 2724 2326
rect 2834 2323 2852 2326
rect 2882 2323 2916 2326
rect 3012 2323 3021 2326
rect 1860 2313 1869 2316
rect 2460 2313 2469 2316
rect 2524 2313 2533 2316
rect 2634 2313 2637 2323
rect 2668 2313 2717 2316
rect 1474 2303 1541 2306
rect 2442 2303 2452 2306
rect 2506 2303 2540 2306
rect 14 2267 3074 2273
rect 1930 2233 1988 2236
rect 2306 2233 2324 2236
rect 2562 2233 2588 2236
rect 116 2213 133 2216
rect 148 2213 157 2216
rect 210 2213 236 2216
rect 498 2213 532 2216
rect 700 2213 725 2216
rect 730 2206 733 2226
rect 868 2223 885 2226
rect 1596 2223 1645 2226
rect 1804 2223 1845 2226
rect 1946 2223 1972 2226
rect 1996 2223 2021 2226
rect 2266 2223 2308 2226
rect 2546 2223 2572 2226
rect 1842 2216 1845 2223
rect 860 2213 869 2216
rect 874 2213 956 2216
rect 1196 2213 1237 2216
rect 1266 2213 1276 2216
rect 1396 2213 1421 2216
rect 1508 2213 1557 2216
rect 1564 2213 1581 2216
rect 1594 2213 1660 2216
rect 1714 2213 1781 2216
rect 1842 2213 1868 2216
rect 2050 2213 2060 2216
rect 2106 2213 2117 2216
rect 2186 2213 2196 2216
rect 2388 2213 2429 2216
rect 2436 2213 2445 2216
rect 2540 2213 2557 2216
rect 2652 2213 2661 2216
rect 2844 2213 2869 2216
rect 2876 2213 2893 2216
rect 1234 2206 1237 2213
rect 380 2203 428 2206
rect 514 2203 524 2206
rect 636 2203 645 2206
rect 730 2203 764 2206
rect 930 2203 948 2206
rect 980 2203 997 2206
rect 1002 2203 1076 2206
rect 1234 2203 1284 2206
rect 1300 2203 1349 2206
rect 1500 2203 1541 2206
rect 1578 2205 1581 2213
rect 1714 2206 1717 2213
rect 1602 2203 1652 2206
rect 1684 2203 1717 2206
rect 1778 2205 1781 2213
rect 2106 2206 2109 2213
rect 1874 2203 1916 2206
rect 2002 2203 2052 2206
rect 2076 2203 2109 2206
rect 2252 2203 2293 2206
rect 2338 2203 2380 2206
rect 2484 2203 2517 2206
rect 2602 2203 2644 2206
rect 2674 2203 2692 2206
rect 2716 2203 2749 2206
rect 2866 2205 2869 2213
rect 346 2193 372 2196
rect 658 2193 684 2196
rect 698 2193 756 2196
rect 1482 2193 1492 2196
rect 1890 2193 1908 2196
rect 2234 2193 2244 2196
rect 2442 2193 2476 2196
rect 38 2167 3050 2173
rect 474 2143 492 2146
rect 538 2136 541 2146
rect 562 2143 604 2146
rect 642 2143 668 2146
rect 1188 2143 1197 2146
rect 1714 2143 1740 2146
rect 1898 2143 1909 2146
rect 2010 2143 2044 2146
rect 2732 2143 2741 2146
rect 212 2133 221 2136
rect 226 2133 276 2136
rect 356 2133 373 2136
rect 538 2133 556 2136
rect 612 2133 669 2136
rect 676 2133 701 2136
rect 988 2133 1045 2136
rect 1098 2133 1172 2136
rect 1268 2133 1325 2136
rect 218 2126 221 2133
rect 370 2126 373 2133
rect 698 2126 701 2133
rect 1330 2126 1333 2135
rect 1356 2133 1389 2136
rect 1484 2133 1493 2136
rect 1578 2133 1604 2136
rect 1628 2133 1653 2136
rect 1658 2133 1684 2136
rect 1698 2133 1748 2136
rect 162 2123 180 2126
rect 218 2123 237 2126
rect 300 2123 349 2126
rect 370 2123 396 2126
rect 698 2123 709 2126
rect 914 2123 964 2126
rect 1042 2123 1068 2126
rect 1146 2123 1164 2126
rect 1188 2123 1252 2126
rect 1298 2123 1333 2126
rect 1412 2123 1460 2126
rect 108 2113 117 2116
rect 148 2113 173 2116
rect 412 2113 421 2116
rect 452 2113 461 2116
rect 1268 2113 1325 2116
rect 1490 2106 1493 2133
rect 1898 2126 1901 2143
rect 1906 2133 1924 2136
rect 2002 2133 2052 2136
rect 2348 2133 2396 2136
rect 2570 2133 2580 2136
rect 2866 2133 2900 2136
rect 2932 2133 2957 2136
rect 1498 2113 1540 2116
rect 1546 2106 1549 2125
rect 1570 2123 1612 2126
rect 1700 2123 1733 2126
rect 1762 2123 1772 2126
rect 1836 2123 1861 2126
rect 1898 2123 1932 2126
rect 1978 2123 1996 2126
rect 2100 2123 2156 2126
rect 2404 2123 2437 2126
rect 2546 2123 2588 2126
rect 1978 2116 1981 2123
rect 1564 2113 1597 2116
rect 1948 2113 1981 2116
rect 2634 2106 2637 2125
rect 2898 2123 2908 2126
rect 2938 2123 3004 2126
rect 1490 2103 1549 2106
rect 2610 2103 2637 2106
rect 14 2067 3074 2073
rect 1506 2033 1540 2036
rect 148 2023 181 2026
rect 860 2023 893 2026
rect 1156 2023 1213 2026
rect 1244 2023 1253 2026
rect 1506 2016 1509 2033
rect 162 2013 188 2016
rect 332 2013 349 2016
rect 468 2013 477 2016
rect 524 2013 533 2016
rect 596 2013 645 2016
rect 698 2006 701 2016
rect 722 2013 732 2016
rect 914 2013 948 2016
rect 1074 2013 1133 2016
rect 1410 2013 1452 2016
rect 1476 2013 1509 2016
rect 1562 2016 1565 2036
rect 1986 2033 2037 2036
rect 2010 2023 2028 2026
rect 1562 2013 1620 2016
rect 1652 2013 1717 2016
rect 1756 2013 1765 2016
rect 1828 2013 1861 2016
rect 1908 2013 1933 2016
rect 1964 2013 2021 2016
rect 2034 2015 2037 2033
rect 2052 2023 2125 2026
rect 2364 2023 2381 2026
rect 2892 2023 2925 2026
rect 2956 2023 2973 2026
rect 2970 2016 2973 2023
rect 2082 2013 2132 2016
rect 2220 2013 2285 2016
rect 2356 2013 2421 2016
rect 2450 2013 2541 2016
rect 1130 2006 1133 2013
rect 2562 2006 2565 2014
rect 2588 2013 2597 2016
rect 2714 2013 2748 2016
rect 2820 2013 2853 2016
rect 2890 2013 2948 2016
rect 2970 2013 2988 2016
rect 220 2003 269 2006
rect 306 2003 324 2006
rect 338 2003 388 2006
rect 442 2003 460 2006
rect 466 2003 516 2006
rect 522 2003 588 2006
rect 652 2003 701 2006
rect 714 2003 724 2006
rect 762 2003 836 2006
rect 906 2003 940 2006
rect 1082 2003 1100 2006
rect 1130 2003 1140 2006
rect 1194 2003 1220 2006
rect 1346 2003 1372 2006
rect 1396 2003 1445 2006
rect 1450 2003 1460 2006
rect 1578 2003 1628 2006
rect 1644 2003 1661 2006
rect 1666 2003 1732 2006
rect 1754 2003 1820 2006
rect 1842 2003 1892 2006
rect 1938 2003 1956 2006
rect 2212 2003 2277 2006
rect 2298 2003 2348 2006
rect 2452 2003 2485 2006
rect 2514 2003 2556 2006
rect 2562 2003 2580 2006
rect 2730 2003 2740 2006
rect 2764 2003 2805 2006
rect 2842 2003 2868 2006
rect 2898 2003 2940 2006
rect 1658 1996 1661 2003
rect 346 1993 380 1996
rect 394 1993 452 1996
rect 466 1993 508 1996
rect 522 1993 580 1996
rect 594 1993 644 1996
rect 1658 1993 1701 1996
rect 1874 1993 1884 1996
rect 2154 1993 2204 1996
rect 2258 1993 2284 1996
rect 38 1967 3050 1973
rect 1146 1953 1173 1956
rect 1170 1946 1173 1953
rect 218 1943 236 1946
rect 1124 1943 1165 1946
rect 1170 1943 1188 1946
rect 1282 1943 1316 1946
rect 1162 1936 1165 1943
rect 114 1933 156 1936
rect 204 1933 244 1936
rect 274 1933 300 1936
rect 426 1933 436 1936
rect 450 1933 492 1936
rect 506 1933 556 1936
rect 706 1933 732 1936
rect 890 1933 948 1936
rect 978 1933 1020 1936
rect 1034 1933 1101 1936
rect 1162 1933 1244 1936
rect 1324 1933 1357 1936
rect 1426 1933 1444 1936
rect 1466 1933 1516 1936
rect 1532 1933 1588 1936
rect 1698 1933 1748 1936
rect 90 1923 108 1926
rect 114 1915 117 1933
rect 354 1923 396 1926
rect 444 1923 477 1926
rect 500 1923 549 1926
rect 564 1923 661 1926
rect 722 1923 740 1926
rect 770 1923 852 1926
rect 882 1923 956 1926
rect 962 1923 1028 1926
rect 1098 1925 1101 1933
rect 1826 1926 1829 1945
rect 2250 1943 2284 1946
rect 2524 1943 2549 1946
rect 1204 1923 1213 1926
rect 1252 1923 1317 1926
rect 1396 1923 1421 1926
rect 1452 1923 1501 1926
rect 1554 1923 1596 1926
rect 1668 1923 1701 1926
rect 1706 1923 1740 1926
rect 1772 1923 1829 1926
rect 1842 1933 1876 1936
rect 1890 1933 1924 1936
rect 2292 1933 2332 1936
rect 2362 1933 2396 1936
rect 2460 1933 2493 1936
rect 2522 1933 2557 1936
rect 2602 1933 2636 1936
rect 1842 1925 1845 1933
rect 1850 1923 1884 1926
rect 1932 1923 1965 1926
rect 1986 1924 2004 1927
rect 964 1913 1021 1916
rect 1036 1913 1085 1916
rect 1698 1906 1701 1923
rect 1986 1916 1989 1924
rect 2026 1923 2092 1926
rect 2188 1923 2197 1926
rect 2300 1923 2309 1926
rect 2340 1923 2397 1926
rect 2404 1923 2429 1926
rect 2522 1925 2525 1933
rect 2538 1923 2572 1926
rect 2586 1923 2644 1926
rect 2682 1923 2732 1926
rect 2860 1923 2877 1926
rect 1962 1913 1989 1916
rect 2020 1913 2037 1916
rect 2348 1913 2381 1916
rect 2874 1913 2900 1916
rect 2906 1906 2909 1925
rect 2954 1923 2964 1926
rect 1698 1903 1733 1906
rect 1946 1903 2012 1906
rect 2898 1903 2909 1906
rect 634 1893 717 1896
rect 14 1867 3074 1873
rect 2714 1853 2733 1856
rect 756 1823 781 1826
rect 940 1823 989 1826
rect 1004 1823 1037 1826
rect 1034 1816 1037 1823
rect 92 1813 109 1816
rect 156 1813 181 1816
rect 228 1813 253 1816
rect 298 1813 348 1816
rect 380 1813 436 1816
rect 468 1813 533 1816
rect 570 1813 644 1816
rect 932 1813 973 1816
rect 986 1813 996 1816
rect 1034 1813 1052 1816
rect 1074 1813 1100 1816
rect 1146 1813 1164 1816
rect 1170 1806 1173 1825
rect 1450 1816 1453 1836
rect 1794 1833 1836 1836
rect 1874 1833 1893 1836
rect 1938 1833 1972 1836
rect 2010 1833 2036 1836
rect 1874 1826 1877 1833
rect 1802 1823 1820 1826
rect 1844 1823 1877 1826
rect 1908 1823 1917 1826
rect 1922 1823 1956 1826
rect 1986 1823 2020 1826
rect 2044 1823 2077 1826
rect 2596 1823 2621 1826
rect 1922 1816 1925 1823
rect 1266 1813 1284 1816
rect 1388 1813 1405 1816
rect 1450 1813 1476 1816
rect 1514 1813 1596 1816
rect 1626 1813 1700 1816
rect 1788 1813 1813 1816
rect 1914 1813 1925 1816
rect 2058 1813 2117 1816
rect 2194 1813 2204 1816
rect 2308 1813 2357 1816
rect 2506 1813 2524 1816
rect 2706 1813 2756 1816
rect 2874 1813 2932 1816
rect 2978 1813 2996 1816
rect 292 1803 325 1806
rect 386 1803 428 1806
rect 498 1803 532 1806
rect 564 1803 581 1806
rect 674 1803 732 1806
rect 860 1803 877 1806
rect 882 1803 924 1806
rect 978 1803 988 1806
rect 1058 1803 1092 1806
rect 1106 1803 1156 1806
rect 1170 1803 1212 1806
rect 1290 1803 1324 1806
rect 1346 1803 1380 1806
rect 1394 1803 1404 1806
rect 1418 1803 1468 1806
rect 1498 1803 1532 1806
rect 1620 1803 1637 1806
rect 1738 1803 1780 1806
rect 2066 1803 2084 1806
rect 2132 1803 2141 1806
rect 2260 1803 2300 1806
rect 2380 1803 2397 1806
rect 2540 1803 2565 1806
rect 2596 1803 2629 1806
rect 2706 1803 2748 1806
rect 2826 1803 2836 1806
rect 2882 1803 2924 1806
rect 1290 1793 1316 1796
rect 2098 1793 2124 1796
rect 2226 1793 2252 1796
rect 2602 1793 2628 1796
rect 38 1767 3050 1773
rect 1114 1743 1141 1746
rect 1490 1743 1556 1746
rect 1586 1743 1597 1746
rect 1786 1743 1844 1746
rect 2314 1743 2324 1746
rect 1114 1736 1117 1743
rect 1594 1736 1597 1743
rect 66 1733 212 1736
rect 226 1733 348 1736
rect 668 1733 740 1736
rect 860 1733 917 1736
rect 922 1733 948 1736
rect 980 1733 997 1736
rect 1002 1733 1068 1736
rect 1100 1733 1117 1736
rect 1122 1733 1180 1736
rect 1204 1733 1213 1736
rect 1322 1733 1356 1736
rect 1386 1733 1460 1736
rect 1564 1733 1589 1736
rect 1594 1733 1620 1736
rect 1658 1733 1676 1736
rect 1690 1733 1756 1736
rect 1780 1733 1789 1736
rect 1852 1733 1900 1736
rect 1922 1733 1956 1736
rect 1986 1733 2028 1736
rect 2138 1733 2156 1736
rect 2252 1733 2309 1736
rect 2322 1733 2332 1736
rect 2404 1733 2421 1736
rect 2650 1733 2676 1736
rect 2786 1733 2796 1736
rect 210 1723 220 1726
rect 748 1723 829 1726
rect 946 1723 956 1726
rect 1018 1723 1076 1726
rect 1130 1723 1188 1726
rect 1434 1723 1452 1726
rect 1484 1723 1549 1726
rect 1628 1723 1637 1726
rect 1706 1723 1764 1726
rect 1908 1723 1917 1726
rect 1964 1723 2021 1726
rect 2036 1723 2093 1726
rect 2178 1723 2236 1726
rect 2322 1723 2325 1733
rect 2698 1726 2716 1727
rect 2858 1726 2861 1736
rect 2340 1723 2397 1726
rect 2642 1724 2716 1726
rect 2642 1723 2701 1724
rect 2738 1723 2804 1726
rect 2858 1723 2884 1726
rect 210 1703 213 1723
rect 228 1713 349 1716
rect 364 1713 509 1716
rect 668 1713 741 1716
rect 1018 1713 1021 1723
rect 1204 1713 1261 1716
rect 1972 1713 1981 1716
rect 2018 1713 2021 1723
rect 2044 1713 2085 1716
rect 2708 1713 2717 1716
rect 14 1667 3074 1673
rect 2322 1633 2348 1636
rect 2362 1633 2381 1636
rect 2610 1633 2676 1636
rect 2378 1626 2381 1633
rect 204 1623 213 1626
rect 1060 1623 1101 1626
rect 1258 1623 1293 1626
rect 1844 1623 1877 1626
rect 2060 1623 2093 1626
rect 2298 1623 2332 1626
rect 2356 1623 2373 1626
rect 2378 1623 2404 1626
rect 2540 1623 2573 1626
rect 2604 1623 2613 1626
rect 2618 1623 2660 1626
rect 1258 1616 1261 1623
rect 2610 1616 2613 1623
rect 108 1613 133 1616
rect 170 1613 188 1616
rect 260 1613 285 1616
rect 322 1613 348 1616
rect 362 1613 373 1616
rect 500 1613 533 1616
rect 778 1613 812 1616
rect 834 1613 852 1616
rect 1026 1613 1044 1616
rect 1074 1613 1132 1616
rect 1210 1613 1228 1616
rect 1252 1613 1261 1616
rect 1266 1613 1308 1616
rect 1428 1613 1445 1616
rect 1476 1613 1509 1616
rect 1540 1613 1565 1616
rect 1754 1613 1796 1616
rect 1802 1613 1836 1616
rect 1916 1613 1965 1616
rect 1980 1613 2021 1616
rect 2122 1613 2156 1616
rect 2434 1613 2484 1616
rect 2538 1613 2596 1616
rect 2610 1613 2629 1616
rect 2690 1613 2724 1616
rect 330 1603 340 1606
rect 362 1605 365 1613
rect 474 1603 492 1606
rect 506 1603 532 1606
rect 690 1603 716 1606
rect 754 1603 804 1606
rect 818 1603 844 1606
rect 868 1603 933 1606
rect 978 1603 1036 1606
rect 1060 1603 1093 1606
rect 1162 1603 1236 1606
rect 690 1593 693 1603
rect 1266 1596 1269 1613
rect 1252 1593 1269 1596
rect 1282 1603 1300 1606
rect 1378 1603 1412 1606
rect 1642 1603 1700 1606
rect 1738 1603 1788 1606
rect 1842 1603 1908 1606
rect 1282 1586 1285 1603
rect 1378 1593 1404 1596
rect 1962 1595 1965 1613
rect 1972 1603 1989 1606
rect 2172 1603 2197 1606
rect 2498 1603 2516 1606
rect 2540 1603 2549 1606
rect 2578 1603 2588 1606
rect 2738 1603 2788 1606
rect 1258 1583 1285 1586
rect 38 1567 3050 1573
rect 1082 1543 1125 1546
rect 1180 1543 1253 1546
rect 1746 1543 1781 1546
rect 2314 1543 2340 1546
rect 1122 1536 1125 1543
rect 1778 1536 1781 1543
rect 226 1533 260 1536
rect 314 1533 332 1536
rect 674 1533 708 1536
rect 740 1533 773 1536
rect 794 1533 820 1536
rect 858 1533 940 1536
rect 964 1533 1037 1536
rect 1076 1533 1117 1536
rect 1122 1533 1164 1536
rect 1290 1533 1364 1536
rect 1388 1533 1453 1536
rect 1484 1533 1525 1536
rect 1580 1533 1637 1536
rect 1652 1533 1708 1536
rect 1732 1533 1773 1536
rect 1778 1533 1796 1536
rect 1834 1533 1908 1536
rect 2106 1533 2116 1536
rect 2180 1533 2189 1536
rect 2348 1533 2373 1536
rect 2434 1533 2476 1536
rect 2506 1533 2572 1536
rect 1450 1526 1453 1533
rect 164 1523 189 1526
rect 234 1523 268 1526
rect 314 1523 340 1526
rect 532 1523 549 1526
rect 626 1523 716 1526
rect 1018 1523 1052 1526
rect 1180 1523 1237 1526
rect 1242 1523 1260 1526
rect 1298 1523 1372 1526
rect 1450 1523 1461 1526
rect 1594 1523 1621 1526
rect 1660 1523 1669 1526
rect 1738 1523 1804 1526
rect 1932 1523 1949 1526
rect 2012 1523 2037 1526
rect 2186 1523 2285 1526
rect 2292 1523 2341 1526
rect 314 1516 317 1523
rect 1594 1516 1597 1523
rect 284 1513 317 1516
rect 1388 1513 1445 1516
rect 1580 1513 1597 1516
rect 2370 1506 2373 1533
rect 2500 1523 2565 1526
rect 2610 1523 2668 1526
rect 2698 1523 2740 1526
rect 2858 1523 2884 1526
rect 2370 1503 2420 1506
rect 14 1467 3074 1473
rect 420 1423 453 1426
rect 556 1423 565 1426
rect 916 1423 981 1426
rect 1108 1423 1165 1426
rect 450 1416 453 1423
rect 1178 1416 1181 1425
rect 1498 1423 1533 1426
rect 2532 1423 2557 1426
rect 1498 1416 1501 1423
rect 116 1413 141 1416
rect 178 1413 212 1416
rect 340 1413 404 1416
rect 450 1413 468 1416
rect 530 1413 540 1416
rect 634 1413 708 1416
rect 762 1413 796 1416
rect 834 1413 900 1416
rect 970 1413 996 1416
rect 1146 1413 1172 1416
rect 1178 1413 1221 1416
rect 218 1403 260 1406
rect 306 1403 332 1406
rect 628 1403 653 1406
rect 748 1403 757 1406
rect 770 1403 788 1406
rect 826 1403 892 1406
rect 916 1403 925 1406
rect 930 1403 988 1406
rect 1020 1403 1037 1406
rect 1050 1403 1092 1406
rect 1218 1405 1221 1413
rect 1266 1413 1301 1416
rect 1332 1413 1357 1416
rect 1442 1413 1460 1416
rect 1492 1413 1501 1416
rect 1506 1413 1572 1416
rect 1610 1413 1652 1416
rect 1676 1413 1725 1416
rect 1732 1413 1781 1416
rect 1266 1405 1269 1413
rect 1354 1406 1357 1413
rect 1274 1403 1308 1406
rect 1354 1403 1380 1406
rect 1402 1403 1468 1406
rect 1484 1403 1501 1406
rect 1554 1403 1564 1406
rect 1588 1403 1613 1406
rect 1618 1403 1660 1406
rect 1698 1403 1724 1406
rect 1778 1405 1781 1413
rect 1802 1413 1853 1416
rect 1866 1413 1924 1416
rect 2140 1413 2181 1416
rect 2242 1413 2284 1416
rect 2330 1413 2381 1416
rect 2452 1413 2493 1416
rect 2506 1413 2516 1416
rect 2658 1413 2668 1416
rect 1802 1405 1805 1413
rect 2802 1406 2805 1414
rect 2810 1413 2876 1416
rect 2892 1413 2901 1416
rect 1810 1403 1852 1406
rect 1882 1403 1932 1406
rect 2068 1403 2116 1406
rect 2242 1403 2276 1406
rect 2370 1403 2388 1406
rect 2498 1403 2508 1406
rect 2532 1403 2541 1406
rect 2714 1403 2780 1406
rect 2802 1403 2868 1406
rect 306 1396 309 1403
rect 1618 1396 1621 1403
rect 276 1393 309 1396
rect 314 1393 324 1396
rect 1346 1393 1372 1396
rect 1594 1393 1621 1396
rect 1676 1393 1685 1396
rect 38 1367 3050 1373
rect 378 1343 412 1346
rect 994 1343 1029 1346
rect 2082 1343 2101 1346
rect 2418 1343 2436 1346
rect 994 1336 997 1343
rect 66 1333 92 1336
rect 146 1333 156 1336
rect 180 1333 189 1336
rect 242 1333 260 1336
rect 370 1333 420 1336
rect 426 1333 460 1336
rect 482 1333 516 1336
rect 722 1333 812 1336
rect 858 1333 932 1336
rect 964 1333 997 1336
rect 1002 1333 1044 1336
rect 1068 1333 1093 1336
rect 1186 1333 1220 1336
rect 1316 1333 1333 1336
rect 1338 1333 1348 1336
rect 1402 1333 1460 1336
rect 1546 1333 1556 1336
rect 1580 1333 1621 1336
rect 1330 1326 1333 1333
rect 1626 1326 1629 1335
rect 1650 1333 1700 1336
rect 1762 1333 1788 1336
rect 1812 1333 1860 1336
rect 1898 1333 1924 1336
rect 1962 1333 2020 1336
rect 2098 1333 2108 1336
rect 2284 1333 2293 1336
rect 2330 1333 2340 1336
rect 2356 1333 2437 1336
rect 2444 1333 2461 1336
rect 1898 1326 1901 1333
rect 2554 1326 2557 1336
rect 2676 1333 2685 1336
rect 2714 1333 2748 1336
rect 2764 1333 2797 1336
rect 2882 1333 2892 1336
rect 100 1323 157 1326
rect 202 1323 228 1326
rect 258 1323 268 1326
rect 108 1313 149 1316
rect 284 1313 333 1316
rect 346 1306 349 1325
rect 468 1323 477 1326
rect 524 1323 533 1326
rect 850 1323 940 1326
rect 970 1323 1052 1326
rect 1098 1323 1148 1326
rect 1218 1323 1228 1326
rect 1330 1323 1349 1326
rect 1442 1323 1452 1326
rect 1484 1323 1493 1326
rect 1506 1323 1564 1326
rect 1602 1323 1629 1326
rect 1636 1323 1645 1326
rect 1730 1323 1796 1326
rect 1868 1323 1901 1326
rect 2044 1323 2077 1326
rect 2090 1323 2116 1326
rect 2180 1323 2237 1326
rect 2266 1323 2332 1326
rect 2538 1323 2548 1326
rect 2554 1323 2612 1326
rect 2682 1323 2685 1333
rect 2810 1326 2813 1333
rect 2772 1323 2813 1326
rect 2900 1323 2917 1326
rect 850 1313 853 1323
rect 1068 1313 1077 1316
rect 1156 1313 1205 1316
rect 1580 1313 1589 1316
rect 2836 1313 2845 1316
rect 306 1303 349 1306
rect 14 1267 3074 1273
rect 372 1223 381 1226
rect 578 1223 605 1226
rect 644 1223 677 1226
rect 972 1223 981 1226
rect 1332 1223 1373 1226
rect 1804 1223 1837 1226
rect 1852 1223 1893 1226
rect 2940 1223 2949 1226
rect 602 1216 605 1223
rect 674 1216 677 1223
rect 1362 1216 1365 1223
rect 140 1213 188 1216
rect 300 1213 333 1216
rect 370 1213 428 1216
rect 564 1213 597 1216
rect 602 1213 628 1216
rect 674 1213 692 1216
rect 818 1213 868 1216
rect 970 1213 1036 1216
rect 1060 1213 1093 1216
rect 1098 1213 1124 1216
rect 1170 1213 1212 1216
rect 1250 1213 1316 1216
rect 1362 1213 1388 1216
rect 1442 1213 1468 1216
rect 1530 1213 1572 1216
rect 1618 1213 1676 1216
rect 1698 1213 1748 1216
rect 1754 1213 1796 1216
rect 1802 1213 1853 1216
rect 1898 1213 1916 1216
rect 1946 1213 2004 1216
rect 2084 1213 2117 1216
rect 2140 1213 2196 1216
rect 2300 1213 2325 1216
rect 2348 1213 2397 1216
rect 330 1206 333 1213
rect 594 1206 597 1213
rect 2114 1207 2117 1213
rect 2402 1206 2405 1214
rect 2436 1213 2453 1216
rect 2482 1213 2500 1216
rect 2506 1213 2524 1216
rect 2548 1213 2573 1216
rect 2612 1213 2637 1216
rect 2708 1213 2733 1216
rect 2770 1213 2796 1216
rect 2866 1206 2869 1214
rect 2874 1213 2924 1216
rect 132 1203 157 1206
rect 266 1203 292 1206
rect 330 1203 348 1206
rect 372 1203 397 1206
rect 444 1203 485 1206
rect 490 1203 500 1206
rect 524 1203 556 1206
rect 594 1203 620 1206
rect 644 1203 653 1206
rect 794 1203 860 1206
rect 922 1203 956 1206
rect 1194 1203 1220 1206
rect 1266 1203 1308 1206
rect 1332 1203 1373 1206
rect 1410 1203 1476 1206
rect 1522 1203 1580 1206
rect 1596 1203 1605 1206
rect 1642 1203 1668 1206
rect 1692 1203 1709 1206
rect 1858 1203 1908 1206
rect 1986 1203 1996 1206
rect 2028 1203 2045 1206
rect 2050 1203 2060 1206
rect 2164 1203 2197 1206
rect 2242 1203 2268 1206
rect 2378 1203 2405 1206
rect 2442 1203 2492 1206
rect 2514 1203 2532 1206
rect 2802 1203 2844 1206
rect 2866 1203 2916 1206
rect 1194 1196 1197 1203
rect 98 1193 124 1196
rect 194 1193 236 1196
rect 1060 1193 1077 1196
rect 1148 1193 1197 1196
rect 2042 1193 2045 1203
rect 38 1167 3050 1173
rect 178 1143 204 1146
rect 140 1133 205 1136
rect 212 1133 221 1136
rect 242 1133 252 1136
rect 266 1133 308 1136
rect 346 1133 372 1136
rect 386 1133 412 1136
rect 442 1133 492 1136
rect 516 1133 549 1136
rect 570 1133 596 1136
rect 666 1133 732 1136
rect 756 1133 773 1136
rect 898 1133 940 1136
rect 964 1133 973 1136
rect 978 1133 1052 1136
rect 1106 1133 1140 1136
rect 1172 1133 1277 1136
rect 1434 1133 1508 1136
rect 1532 1133 1597 1136
rect 1628 1133 1709 1136
rect 1732 1133 1804 1136
rect 108 1123 133 1126
rect 220 1123 229 1126
rect 234 1123 260 1126
rect 330 1123 420 1126
rect 514 1123 564 1126
rect 604 1123 653 1126
rect 660 1123 733 1126
rect 828 1123 837 1126
rect 890 1123 948 1126
rect 978 1116 981 1133
rect 1826 1126 1829 1145
rect 2460 1143 2485 1146
rect 2626 1143 2653 1146
rect 2626 1136 2629 1143
rect 2650 1136 2653 1143
rect 1954 1133 1996 1136
rect 2138 1133 2156 1136
rect 2194 1133 2228 1136
rect 2282 1133 2292 1136
rect 2370 1126 2373 1136
rect 2618 1133 2629 1136
rect 994 1123 1060 1126
rect 1138 1123 1148 1126
rect 1340 1123 1397 1126
rect 1428 1123 1501 1126
rect 1506 1123 1516 1126
rect 1586 1123 1604 1126
rect 1698 1123 1708 1126
rect 1812 1123 1829 1126
rect 1844 1123 1853 1126
rect 1866 1123 1924 1126
rect 2020 1123 2029 1126
rect 2076 1123 2085 1126
rect 2324 1123 2373 1126
rect 2378 1123 2388 1126
rect 2394 1123 2436 1126
rect 2460 1123 2485 1126
rect 2586 1123 2596 1126
rect 2618 1125 2621 1133
rect 2634 1126 2637 1136
rect 2650 1133 2660 1136
rect 2714 1133 2740 1136
rect 2756 1133 2781 1136
rect 2882 1133 2892 1136
rect 2810 1126 2813 1133
rect 2634 1123 2668 1126
rect 2764 1123 2813 1126
rect 2900 1123 2917 1126
rect 332 1113 357 1116
rect 436 1113 453 1116
rect 516 1113 525 1116
rect 964 1113 981 1116
rect 2466 1103 2525 1106
rect 14 1067 3074 1073
rect 1394 1053 1437 1056
rect 338 1033 365 1036
rect 322 1023 356 1026
rect 108 1013 133 1016
rect 212 1013 269 1016
rect 362 1015 365 1033
rect 508 1023 541 1026
rect 972 1023 997 1026
rect 1068 1023 1077 1026
rect 1714 1023 1733 1026
rect 2452 1023 2461 1026
rect 2844 1023 2853 1026
rect 538 1016 541 1023
rect 1730 1016 1733 1023
rect 428 1013 485 1016
rect 538 1013 564 1016
rect 636 1013 661 1016
rect 794 1013 860 1016
rect 898 1013 956 1016
rect 978 1013 1052 1016
rect 1106 1013 1148 1016
rect 1162 1013 1252 1016
rect 1282 1013 1364 1016
rect 1500 1013 1525 1016
rect 1530 1013 1580 1016
rect 1612 1013 1621 1016
rect 1692 1013 1725 1016
rect 1730 1013 1740 1016
rect 1764 1013 1813 1016
rect 1850 1013 1876 1016
rect 2034 1013 2052 1016
rect 2116 1013 2149 1016
rect 2188 1013 2221 1016
rect 2228 1013 2269 1016
rect 2292 1013 2341 1016
rect 2372 1013 2429 1016
rect 2450 1013 2492 1016
rect 2660 1013 2685 1016
rect 2788 1013 2821 1016
rect 2908 1013 2917 1016
rect 194 1003 204 1006
rect 218 1003 268 1006
rect 482 1005 485 1013
rect 722 1003 748 1006
rect 780 1003 813 1006
rect 890 1003 948 1006
rect 1068 1003 1101 1006
rect 1164 1003 1181 1006
rect 1314 1003 1356 1006
rect 1562 1003 1588 1006
rect 1610 1003 1668 1006
rect 1738 1003 1748 1006
rect 1810 1005 1813 1013
rect 2426 1007 2429 1013
rect 2818 1007 2821 1013
rect 1858 1003 1868 1006
rect 1900 1003 1909 1006
rect 2140 1003 2180 1006
rect 2210 1003 2220 1006
rect 2316 1003 2325 1006
rect 2508 1003 2525 1006
rect 2746 1003 2764 1006
rect 2890 1003 2900 1006
rect 1764 993 1773 996
rect 2372 993 2381 996
rect 38 967 3050 973
rect 2770 953 2853 956
rect 370 943 380 946
rect 1780 943 1797 946
rect 162 933 188 936
rect 378 933 388 936
rect 394 933 404 936
rect 578 933 588 936
rect 634 933 644 936
rect 834 933 860 936
rect 892 933 917 936
rect 1004 933 1077 936
rect 1116 933 1173 936
rect 1178 933 1188 936
rect 1226 933 1300 936
rect 1338 933 1412 936
rect 1428 933 1453 936
rect 1618 933 1676 936
rect 1698 933 1764 936
rect 1852 933 1893 936
rect 378 926 381 933
rect 1898 926 1901 935
rect 1924 933 1957 936
rect 2012 933 2028 936
rect 2050 933 2100 936
rect 2138 933 2180 936
rect 2234 933 2276 936
rect 2314 933 2356 936
rect 2698 933 2876 936
rect 170 923 196 926
rect 276 923 293 926
rect 362 923 381 926
rect 402 923 412 926
rect 492 923 509 926
rect 548 923 557 926
rect 596 923 645 926
rect 740 923 765 926
rect 842 923 868 926
rect 898 923 980 926
rect 1018 923 1092 926
rect 1162 923 1196 926
rect 1282 923 1308 926
rect 1500 923 1557 926
rect 1658 923 1668 926
rect 1706 923 1756 926
rect 1810 923 1836 926
rect 1850 923 1901 926
rect 1988 923 2029 926
rect 2058 923 2108 926
rect 2204 923 2284 926
rect 2452 923 2461 926
rect 2602 923 2628 926
rect 2756 923 2789 926
rect 2900 923 2941 926
rect 2954 923 2957 935
rect 170 916 173 923
rect 140 913 173 916
rect 604 913 637 916
rect 1852 913 1885 916
rect 14 867 3074 873
rect 220 823 253 826
rect 276 823 309 826
rect 364 823 389 826
rect 420 823 453 826
rect 522 823 549 826
rect 1052 823 1117 826
rect 250 816 253 823
rect 306 816 309 823
rect 546 816 549 823
rect 108 813 133 816
rect 164 813 197 816
rect 250 813 268 816
rect 306 813 324 816
rect 460 813 501 816
rect 508 813 541 816
rect 546 813 556 816
rect 634 813 652 816
rect 700 813 741 816
rect 748 813 821 816
rect 994 813 1044 816
rect 1114 806 1117 823
rect 1154 823 1189 826
rect 2788 823 2797 826
rect 1154 816 1157 823
rect 1124 813 1157 816
rect 1162 813 1284 816
rect 1354 813 1396 816
rect 1466 813 1492 816
rect 1708 813 1717 816
rect 1810 813 1876 816
rect 1964 813 2045 816
rect 2060 813 2077 816
rect 2124 813 2173 816
rect 2204 813 2229 816
rect 2252 813 2293 816
rect 2348 813 2389 816
rect 2404 813 2429 816
rect 226 803 260 806
rect 370 803 404 806
rect 466 803 500 806
rect 562 803 604 806
rect 626 803 644 806
rect 658 803 692 806
rect 754 803 820 806
rect 1098 805 1117 806
rect 1098 803 1116 805
rect 1178 803 1196 806
rect 1234 803 1276 806
rect 1420 803 1485 806
rect 1490 803 1500 806
rect 1570 803 1612 806
rect 1626 803 1700 806
rect 1706 803 1788 806
rect 1842 803 1868 806
rect 1882 803 1940 806
rect 1650 793 1692 796
rect 1706 793 1780 796
rect 2042 795 2045 813
rect 2226 807 2229 813
rect 2458 806 2461 816
rect 2466 813 2476 816
rect 2516 813 2541 816
rect 2580 813 2605 816
rect 2642 813 2668 816
rect 2724 813 2765 816
rect 2762 807 2765 813
rect 2898 806 2901 814
rect 2906 813 2940 816
rect 2052 803 2085 806
rect 2354 803 2461 806
rect 2492 803 2508 806
rect 2716 803 2757 806
rect 2850 803 2876 806
rect 2898 803 2932 806
rect 38 767 3050 773
rect 1290 753 1381 756
rect 546 743 581 746
rect 578 736 581 743
rect 2626 743 2660 746
rect 2674 743 2732 746
rect 298 733 340 736
rect 370 733 420 736
rect 458 733 516 736
rect 540 733 573 736
rect 578 733 596 736
rect 620 733 653 736
rect 674 733 684 736
rect 708 733 748 736
rect 818 733 876 736
rect 900 733 917 736
rect 1114 733 1164 736
rect 1250 733 1260 736
rect 1284 733 1301 736
rect 1564 733 1581 736
rect 1586 733 1636 736
rect 298 726 301 733
rect 1586 726 1589 733
rect 1650 726 1653 736
rect 1802 733 1836 736
rect 1860 733 1917 736
rect 1970 733 2004 736
rect 2170 733 2212 736
rect 2234 733 2284 736
rect 2298 733 2348 736
rect 2372 733 2381 736
rect 2450 733 2476 736
rect 2490 733 2532 736
rect 2570 733 2612 736
rect 1802 726 1805 733
rect 2626 726 2629 743
rect 2650 733 2740 736
rect 210 723 228 726
rect 276 723 301 726
rect 306 723 348 726
rect 410 723 428 726
rect 482 723 524 726
rect 594 723 604 726
rect 618 723 692 726
rect 756 723 805 726
rect 812 723 877 726
rect 988 723 1005 726
rect 1044 723 1077 726
rect 1092 723 1117 726
rect 1162 723 1172 726
rect 1186 723 1268 726
rect 1572 723 1589 726
rect 1644 723 1653 726
rect 1732 723 1749 726
rect 1788 723 1805 726
rect 1826 723 1844 726
rect 1906 723 1932 726
rect 1962 723 2012 726
rect 2068 723 2077 726
rect 2220 723 2285 726
rect 2292 723 2356 726
rect 2410 723 2444 726
rect 2466 723 2484 726
rect 2562 723 2629 726
rect 2676 723 2725 726
rect 2828 723 2853 726
rect 2410 716 2413 723
rect 2466 716 2469 723
rect 284 713 325 716
rect 364 713 397 716
rect 1284 713 1317 716
rect 2076 713 2140 716
rect 2164 713 2213 716
rect 2372 713 2413 716
rect 2452 713 2469 716
rect 2556 713 2581 716
rect 2098 703 2156 706
rect 14 667 3074 673
rect 2194 633 2245 636
rect 2674 633 2725 636
rect 228 623 253 626
rect 556 623 589 626
rect 620 623 653 626
rect 996 623 1045 626
rect 1292 623 1325 626
rect 1532 623 1573 626
rect 1612 623 1621 626
rect 1756 623 1797 626
rect 1836 623 1853 626
rect 2202 623 2236 626
rect 250 616 253 623
rect 586 616 589 623
rect 650 616 653 623
rect 1042 616 1045 623
rect 1570 616 1573 623
rect 116 613 141 616
rect 172 613 205 616
rect 250 613 268 616
rect 298 613 340 616
rect 346 613 364 616
rect 444 613 469 616
rect 500 613 517 616
rect 522 613 540 616
rect 586 613 612 616
rect 650 613 668 616
rect 674 613 716 616
rect 746 613 804 616
rect 892 613 973 616
rect 1042 613 1084 616
rect 1162 613 1172 616
rect 1306 613 1364 616
rect 1388 613 1421 616
rect 1466 613 1516 616
rect 1570 613 1596 616
rect 1676 613 1685 616
rect 1714 613 1740 616
rect 1762 613 1820 616
rect 2068 613 2101 616
rect 2108 613 2117 616
rect 2154 613 2229 616
rect 2242 615 2245 633
rect 2260 623 2293 626
rect 2682 623 2716 626
rect 2316 613 2325 616
rect 2484 613 2509 616
rect 2540 613 2565 616
rect 2722 615 2725 633
rect 2740 623 2749 626
rect 2810 623 2844 626
rect 234 603 260 606
rect 322 603 332 606
rect 570 603 604 606
rect 674 603 708 606
rect 738 603 796 606
rect 820 603 884 606
rect 970 605 973 613
rect 2746 606 2749 623
rect 2874 613 2924 616
rect 2930 613 2956 616
rect 2978 606 2981 614
rect 996 603 1005 606
rect 1292 603 1372 606
rect 1386 603 1420 606
rect 1468 603 1477 606
rect 1490 603 1508 606
rect 1532 603 1565 606
rect 1570 603 1588 606
rect 1836 603 1845 606
rect 2082 603 2100 606
rect 2122 603 2140 606
rect 2266 603 2308 606
rect 2570 603 2580 606
rect 2634 603 2652 606
rect 2746 603 2780 606
rect 2978 603 2989 606
rect 1570 596 1573 603
rect 1388 593 1413 596
rect 1538 593 1573 596
rect 2290 593 2300 596
rect 2668 593 2709 596
rect 2986 593 2989 603
rect 38 567 3050 573
rect 1418 553 1437 556
rect 1434 536 1437 553
rect 1578 543 1644 546
rect 2732 543 2757 546
rect 346 533 372 536
rect 396 533 453 536
rect 484 533 516 536
rect 538 533 572 536
rect 596 533 636 536
rect 722 526 725 535
rect 748 533 781 536
rect 930 533 956 536
rect 980 533 1005 536
rect 1154 533 1188 536
rect 1220 533 1245 536
rect 1250 533 1284 536
rect 1316 533 1341 536
rect 1378 533 1388 536
rect 1412 533 1429 536
rect 1434 533 1452 536
rect 1474 533 1532 536
rect 1570 533 1652 536
rect 1706 533 1748 536
rect 1956 533 2013 536
rect 2218 533 2252 536
rect 2276 533 2309 536
rect 2618 533 2652 536
rect 2658 533 2709 536
rect 2858 533 2876 536
rect 2946 533 2957 536
rect 1474 526 1477 533
rect 116 523 141 526
rect 172 523 197 526
rect 202 523 236 526
rect 322 523 380 526
rect 514 523 524 526
rect 660 523 725 526
rect 778 523 796 526
rect 930 523 964 526
rect 1002 523 1020 526
rect 1170 523 1196 526
rect 1234 523 1292 526
rect 1322 523 1396 526
rect 1460 523 1477 526
rect 1668 523 1693 526
rect 1714 523 1756 526
rect 1954 523 2028 526
rect 2108 523 2133 526
rect 778 516 781 523
rect 1002 516 1005 523
rect 748 513 781 516
rect 980 513 1005 516
rect 1956 513 2021 516
rect 2036 513 2077 516
rect 2130 506 2133 523
rect 2138 513 2164 516
rect 2170 506 2173 525
rect 2194 523 2260 526
rect 2460 523 2485 526
rect 2556 523 2581 526
rect 2612 523 2621 526
rect 2660 523 2701 526
rect 2706 525 2709 533
rect 2954 526 2957 533
rect 2796 523 2821 526
rect 2884 523 2909 526
rect 2954 523 2996 526
rect 2188 513 2245 516
rect 2130 503 2173 506
rect 14 467 3074 473
rect 2258 433 2308 436
rect 242 416 245 426
rect 556 423 589 426
rect 700 423 733 426
rect 1060 423 1101 426
rect 1140 423 1149 426
rect 1364 423 1389 426
rect 1804 423 1829 426
rect 2020 423 2069 426
rect 2100 423 2125 426
rect 2292 423 2301 426
rect 2820 423 2837 426
rect 586 416 589 423
rect 1098 416 1101 423
rect 92 413 157 416
rect 194 413 260 416
rect 436 413 461 416
rect 492 413 533 416
rect 554 413 565 416
rect 586 413 612 416
rect 618 413 684 416
rect 706 413 780 416
rect 852 413 869 416
rect 972 413 1037 416
rect 1098 413 1132 416
rect 1170 413 1236 416
rect 1266 413 1348 416
rect 1426 413 1444 416
rect 1468 413 1493 416
rect 1506 413 1580 416
rect 1676 413 1701 416
rect 1738 413 1788 416
rect 1938 413 1996 416
rect 2026 413 2092 416
rect 2180 413 2197 416
rect 2202 413 2228 416
rect 2410 413 2428 416
rect 2508 413 2533 416
rect 2620 413 2685 416
rect 74 403 84 406
rect 154 405 157 413
rect 562 406 565 413
rect 188 403 205 406
rect 514 403 532 406
rect 562 403 604 406
rect 658 403 676 406
rect 700 403 765 406
rect 796 403 805 406
rect 810 403 844 406
rect 858 403 892 406
rect 930 403 964 406
rect 1034 405 1037 413
rect 1060 403 1069 406
rect 1170 403 1173 413
rect 2690 406 2693 414
rect 2898 413 2908 416
rect 1178 403 1228 406
rect 1330 403 1340 406
rect 1364 403 1452 406
rect 1482 403 1572 406
rect 1804 403 1837 406
rect 1962 403 1988 406
rect 2074 403 2084 406
rect 2106 403 2164 406
rect 2578 403 2612 406
rect 2674 403 2693 406
rect 2754 403 2796 406
rect 2820 403 2829 406
rect 2906 403 2916 406
rect 1178 386 1181 403
rect 2594 393 2604 396
rect 1146 383 1181 386
rect 38 367 3050 373
rect 1978 343 1988 346
rect 2138 343 2196 346
rect 2258 343 2300 346
rect 2402 343 2428 346
rect 2818 343 2837 346
rect 2834 336 2837 343
rect 106 333 148 336
rect 202 333 236 336
rect 460 333 508 336
rect 572 333 613 336
rect 618 333 628 336
rect 652 333 685 336
rect 722 333 764 336
rect 788 333 805 336
rect 810 333 828 336
rect 866 333 876 336
rect 900 333 925 336
rect 1130 333 1164 336
rect 1300 333 1333 336
rect 1354 333 1364 336
rect 1388 333 1437 336
rect 1468 333 1524 336
rect 1666 333 1692 336
rect 1778 333 1820 336
rect 1834 333 1852 336
rect 1970 333 1996 336
rect 2178 333 2204 336
rect 2258 333 2308 336
rect 2314 333 2348 336
rect 2410 333 2436 336
rect 618 326 621 333
rect 90 323 100 326
rect 178 323 228 326
rect 252 323 293 326
rect 306 323 340 326
rect 362 323 372 326
rect 516 323 549 326
rect 570 323 621 326
rect 626 323 636 326
rect 650 323 700 326
rect 746 323 772 326
rect 836 323 877 326
rect 1234 323 1276 326
rect 1306 323 1372 326
rect 1386 323 1452 326
rect 1522 323 1532 326
rect 1764 323 1773 326
rect 1786 323 1828 326
rect 172 313 197 316
rect 460 313 485 316
rect 572 313 597 316
rect 716 313 733 316
rect 1468 313 1509 316
rect 1716 313 1733 316
rect 1772 313 1813 316
rect 1834 315 1837 333
rect 2098 326 2116 327
rect 2682 326 2685 335
rect 2714 333 2788 336
rect 2804 333 2829 336
rect 2834 333 2876 336
rect 2900 333 2909 336
rect 2004 323 2060 326
rect 2066 324 2116 326
rect 2066 323 2101 324
rect 2218 323 2252 326
rect 2316 323 2333 326
rect 2652 323 2685 326
rect 2692 323 2701 326
rect 2708 323 2725 326
rect 2818 323 2884 326
rect 2908 323 2917 326
rect 1866 313 1916 316
rect 2066 315 2069 323
rect 2074 313 2108 316
rect 2090 303 2124 306
rect 14 267 3074 273
rect 154 233 173 236
rect 250 233 292 236
rect 1426 233 1452 236
rect 2426 233 2477 236
rect 2770 233 2797 236
rect 154 226 157 233
rect 116 223 157 226
rect 250 206 253 233
rect 266 223 276 226
rect 300 223 349 226
rect 572 223 597 226
rect 594 216 597 223
rect 306 213 364 216
rect 378 213 396 216
rect 538 213 556 216
rect 594 213 612 216
rect 700 213 757 216
rect 770 206 773 225
rect 916 223 925 226
rect 1346 223 1436 226
rect 1460 223 1477 226
rect 1554 216 1557 225
rect 1562 223 1636 226
rect 1740 223 1773 226
rect 1812 223 1861 226
rect 2268 223 2325 226
rect 2450 223 2468 226
rect 2450 216 2453 223
rect 786 213 828 216
rect 908 213 957 216
rect 1122 213 1172 216
rect 1506 213 1548 216
rect 1554 213 1644 216
rect 1794 213 1804 216
rect 1818 213 1884 216
rect 1964 213 1973 216
rect 2084 213 2117 216
rect 2122 213 2140 216
rect 228 203 253 206
rect 314 203 356 206
rect 578 203 604 206
rect 618 203 676 206
rect 770 203 820 206
rect 922 203 956 206
rect 980 203 1021 206
rect 1298 203 1316 206
rect 1698 203 1724 206
rect 1786 203 1796 206
rect 1810 203 1876 206
rect 2066 203 2076 206
rect 2138 203 2148 206
rect 2162 203 2244 206
rect 2268 203 2325 206
rect 2330 205 2333 216
rect 2354 213 2413 216
rect 2420 213 2453 216
rect 2474 215 2477 233
rect 2778 223 2788 226
rect 2634 213 2652 216
rect 2410 205 2413 213
rect 2634 203 2644 206
rect 2698 203 2701 214
rect 2724 213 2741 216
rect 2794 215 2797 233
rect 2898 206 2901 214
rect 2818 203 2892 206
rect 2898 203 2948 206
rect 194 193 220 196
rect 2826 193 2884 196
rect 38 167 3050 173
rect 882 143 916 146
rect 2546 143 2556 146
rect 2946 143 2972 146
rect 186 126 189 135
rect 266 133 276 136
rect 386 133 396 136
rect 682 133 692 136
rect 722 133 732 136
rect 882 133 924 136
rect 1020 133 1061 136
rect 1274 133 1284 136
rect 1396 133 1421 136
rect 1602 133 1612 136
rect 1650 133 1660 136
rect 1818 133 1828 136
rect 2050 133 2068 136
rect 2092 133 2109 136
rect 2138 133 2156 136
rect 2564 133 2589 136
rect 2706 133 2756 136
rect 2772 133 2781 136
rect 172 123 189 126
rect 236 123 277 126
rect 308 123 349 126
rect 346 106 349 123
rect 362 106 365 125
rect 500 123 525 126
rect 556 123 565 126
rect 604 123 629 126
rect 660 123 693 126
rect 730 123 740 126
rect 820 123 845 126
rect 962 123 1004 126
rect 1058 123 1084 126
rect 1220 123 1261 126
rect 1292 123 1380 126
rect 1394 123 1436 126
rect 1562 123 1596 126
rect 1668 123 1693 126
rect 1796 123 1805 126
rect 1884 123 1893 126
rect 2122 123 2164 126
rect 2468 123 2477 126
rect 2524 123 2557 126
rect 2572 123 2581 126
rect 730 116 733 123
rect 1058 116 1061 123
rect 716 113 733 116
rect 1020 113 1061 116
rect 1092 113 1125 116
rect 1396 113 1405 116
rect 1676 113 1685 116
rect 1844 113 1861 116
rect 2092 113 2149 116
rect 2202 113 2252 116
rect 2586 106 2589 133
rect 2674 123 2700 126
rect 2780 123 2789 126
rect 2802 123 2860 126
rect 2898 123 2932 126
rect 2898 116 2901 123
rect 2610 113 2620 116
rect 2876 113 2901 116
rect 346 103 365 106
rect 2186 103 2268 106
rect 2586 103 2636 106
rect 14 67 3074 73
rect 38 37 3050 57
rect 14 13 3074 33
<< metal2 >>
rect 2 3033 77 3036
rect 2 1883 5 3033
rect 14 13 34 3027
rect 38 37 58 3003
rect 74 2946 77 3033
rect 66 2943 77 2946
rect 146 2943 181 2946
rect 66 2773 69 2943
rect 82 2906 85 2926
rect 154 2916 157 2936
rect 162 2923 173 2926
rect 178 2923 181 2943
rect 194 2933 197 2956
rect 282 2933 285 2956
rect 426 2943 461 2946
rect 290 2926 293 2936
rect 354 2933 397 2936
rect 154 2913 173 2916
rect 82 2903 93 2906
rect 90 2836 93 2903
rect 82 2833 93 2836
rect 66 2333 69 2756
rect 82 2676 85 2833
rect 90 2813 125 2816
rect 146 2813 149 2836
rect 170 2823 173 2913
rect 210 2823 213 2836
rect 250 2816 253 2926
rect 258 2923 293 2926
rect 322 2903 325 2926
rect 114 2753 117 2806
rect 122 2803 125 2813
rect 154 2776 157 2816
rect 210 2813 221 2816
rect 250 2813 261 2816
rect 242 2793 245 2806
rect 250 2786 253 2813
rect 242 2783 253 2786
rect 290 2786 293 2816
rect 314 2813 317 2836
rect 330 2826 333 2926
rect 354 2913 357 2933
rect 386 2903 389 2916
rect 450 2883 453 2926
rect 458 2923 461 2943
rect 314 2793 317 2806
rect 322 2786 325 2826
rect 330 2823 373 2826
rect 410 2823 413 2836
rect 290 2783 325 2786
rect 154 2773 181 2776
rect 90 2723 93 2746
rect 74 2673 85 2676
rect 74 2506 77 2673
rect 90 2606 93 2636
rect 98 2613 101 2626
rect 114 2613 117 2736
rect 138 2733 141 2746
rect 146 2703 149 2726
rect 154 2666 157 2726
rect 178 2713 181 2773
rect 210 2726 213 2746
rect 226 2733 229 2746
rect 210 2723 221 2726
rect 210 2703 213 2716
rect 154 2663 173 2666
rect 170 2623 173 2663
rect 82 2603 101 2606
rect 98 2526 101 2596
rect 98 2523 109 2526
rect 114 2506 117 2596
rect 74 2503 85 2506
rect 82 2436 85 2503
rect 74 2433 85 2436
rect 106 2503 117 2506
rect 74 2353 77 2433
rect 106 2406 109 2503
rect 130 2406 133 2536
rect 162 2416 165 2546
rect 178 2533 181 2616
rect 186 2533 189 2606
rect 202 2593 205 2636
rect 242 2596 245 2783
rect 298 2733 301 2746
rect 354 2743 357 2816
rect 418 2813 421 2826
rect 442 2793 445 2806
rect 322 2733 341 2736
rect 274 2716 277 2726
rect 290 2723 301 2726
rect 306 2716 309 2726
rect 274 2713 309 2716
rect 338 2703 341 2733
rect 378 2723 389 2726
rect 306 2633 341 2636
rect 250 2613 285 2616
rect 306 2613 309 2633
rect 338 2613 341 2633
rect 402 2626 405 2736
rect 418 2723 421 2746
rect 426 2703 429 2716
rect 394 2623 405 2626
rect 242 2593 261 2596
rect 274 2593 277 2606
rect 282 2603 285 2613
rect 194 2543 221 2546
rect 210 2446 213 2526
rect 218 2523 221 2543
rect 242 2533 245 2546
rect 258 2523 261 2593
rect 354 2566 357 2606
rect 362 2593 365 2616
rect 386 2596 389 2606
rect 394 2603 397 2623
rect 402 2596 405 2616
rect 418 2613 421 2626
rect 466 2613 469 2936
rect 490 2933 493 2976
rect 626 2963 661 2966
rect 506 2933 509 2956
rect 498 2923 509 2926
rect 490 2823 525 2826
rect 490 2813 493 2823
rect 506 2813 517 2816
rect 522 2813 525 2823
rect 514 2793 517 2806
rect 554 2756 557 2936
rect 610 2916 613 2926
rect 618 2923 621 2936
rect 626 2923 629 2963
rect 650 2933 653 2956
rect 658 2933 661 2963
rect 642 2923 653 2926
rect 658 2916 661 2926
rect 586 2836 589 2916
rect 610 2913 661 2916
rect 578 2833 589 2836
rect 682 2836 685 2936
rect 714 2913 725 2916
rect 746 2913 749 2926
rect 778 2923 781 2936
rect 810 2933 813 2976
rect 786 2896 789 2926
rect 810 2903 813 2926
rect 818 2913 821 2926
rect 826 2896 829 2936
rect 874 2933 917 2936
rect 874 2913 877 2933
rect 906 2903 909 2916
rect 786 2893 845 2896
rect 682 2833 725 2836
rect 578 2806 581 2833
rect 594 2813 613 2816
rect 666 2813 669 2826
rect 562 2803 581 2806
rect 578 2793 581 2803
rect 626 2766 629 2806
rect 610 2763 629 2766
rect 554 2753 581 2756
rect 490 2733 501 2736
rect 506 2726 509 2736
rect 474 2723 509 2726
rect 514 2706 517 2726
rect 546 2706 549 2726
rect 514 2703 549 2706
rect 562 2716 565 2736
rect 570 2723 573 2746
rect 578 2733 581 2753
rect 610 2733 613 2763
rect 674 2756 677 2816
rect 698 2793 701 2806
rect 658 2753 677 2756
rect 602 2716 605 2726
rect 562 2713 605 2716
rect 610 2713 613 2726
rect 618 2716 621 2736
rect 658 2733 661 2753
rect 618 2713 661 2716
rect 562 2616 565 2713
rect 482 2613 565 2616
rect 602 2613 605 2626
rect 618 2613 621 2656
rect 386 2593 405 2596
rect 418 2593 421 2606
rect 506 2593 509 2606
rect 346 2563 357 2566
rect 338 2533 341 2546
rect 346 2526 349 2563
rect 314 2523 349 2526
rect 202 2443 213 2446
rect 146 2413 181 2416
rect 106 2403 125 2406
rect 130 2403 141 2406
rect 122 2333 125 2403
rect 90 2193 93 2326
rect 122 2306 125 2326
rect 114 2303 125 2306
rect 114 2226 117 2303
rect 114 2223 125 2226
rect 98 2203 117 2206
rect 82 2133 85 2176
rect 90 2096 93 2126
rect 114 2113 117 2203
rect 122 2173 125 2223
rect 90 2093 109 2096
rect 106 2023 109 2093
rect 82 1983 85 2006
rect 90 1923 93 2016
rect 130 2006 133 2216
rect 138 2203 141 2403
rect 154 2323 157 2356
rect 170 2226 173 2406
rect 178 2403 181 2413
rect 202 2386 205 2443
rect 218 2433 253 2436
rect 218 2413 221 2433
rect 250 2413 253 2433
rect 274 2413 277 2426
rect 202 2383 213 2386
rect 210 2346 213 2383
rect 186 2343 221 2346
rect 186 2323 189 2343
rect 194 2333 213 2336
rect 146 2223 173 2226
rect 146 2196 149 2223
rect 122 2003 133 2006
rect 142 2193 149 2196
rect 154 2196 157 2216
rect 194 2203 197 2333
rect 154 2193 165 2196
rect 98 1933 101 1946
rect 82 1913 117 1916
rect 82 1803 85 1913
rect 106 1786 109 1816
rect 122 1813 125 2003
rect 142 1996 145 2193
rect 162 2146 165 2193
rect 138 1993 145 1996
rect 154 2143 165 2146
rect 138 1933 141 1993
rect 154 1983 157 2143
rect 162 2093 165 2126
rect 186 2123 189 2176
rect 202 2146 205 2216
rect 210 2213 213 2226
rect 218 2183 221 2343
rect 266 2333 269 2406
rect 314 2403 317 2436
rect 322 2413 325 2523
rect 426 2506 429 2536
rect 482 2533 517 2536
rect 458 2513 461 2526
rect 466 2506 469 2526
rect 426 2503 469 2506
rect 314 2233 317 2346
rect 330 2336 333 2416
rect 418 2393 421 2416
rect 426 2403 429 2503
rect 474 2343 477 2436
rect 514 2376 517 2533
rect 538 2513 541 2613
rect 626 2606 629 2646
rect 650 2613 653 2626
rect 586 2603 629 2606
rect 658 2603 661 2713
rect 706 2643 709 2736
rect 714 2723 717 2816
rect 722 2813 725 2833
rect 754 2813 757 2826
rect 738 2793 741 2806
rect 794 2786 797 2816
rect 818 2793 821 2806
rect 794 2783 821 2786
rect 730 2613 733 2756
rect 754 2753 813 2756
rect 754 2733 757 2753
rect 762 2733 765 2746
rect 810 2706 813 2753
rect 818 2733 821 2783
rect 818 2716 821 2726
rect 826 2723 829 2746
rect 834 2716 837 2816
rect 842 2813 845 2893
rect 930 2866 933 2946
rect 954 2923 957 2936
rect 978 2923 981 2936
rect 1026 2913 1029 2926
rect 1058 2876 1061 2966
rect 1130 2963 1133 3040
rect 1050 2873 1061 2876
rect 930 2863 965 2866
rect 882 2813 885 2826
rect 866 2793 869 2806
rect 914 2756 917 2816
rect 938 2793 941 2806
rect 818 2713 837 2716
rect 842 2706 845 2736
rect 810 2703 845 2706
rect 794 2633 829 2636
rect 570 2506 573 2526
rect 594 2513 597 2526
rect 602 2506 605 2526
rect 570 2503 605 2506
rect 618 2506 621 2536
rect 626 2513 629 2603
rect 658 2533 677 2536
rect 634 2523 653 2526
rect 634 2506 637 2523
rect 618 2503 637 2506
rect 634 2436 637 2503
rect 634 2433 645 2436
rect 642 2416 645 2433
rect 514 2373 525 2376
rect 530 2353 533 2406
rect 538 2403 541 2416
rect 506 2343 533 2346
rect 546 2343 549 2416
rect 634 2413 645 2416
rect 634 2393 637 2413
rect 618 2343 621 2376
rect 330 2333 341 2336
rect 506 2333 509 2343
rect 226 2203 229 2216
rect 202 2143 221 2146
rect 210 2116 213 2126
rect 170 2113 213 2116
rect 218 2046 221 2143
rect 226 2113 229 2136
rect 234 2096 237 2126
rect 242 2116 245 2216
rect 338 2203 341 2333
rect 330 2183 333 2196
rect 282 2123 285 2136
rect 290 2133 293 2146
rect 338 2136 341 2196
rect 346 2166 349 2236
rect 354 2193 357 2326
rect 378 2303 381 2326
rect 386 2243 389 2326
rect 450 2223 453 2306
rect 514 2303 517 2336
rect 458 2226 461 2246
rect 458 2223 469 2226
rect 362 2213 389 2216
rect 346 2163 357 2166
rect 346 2143 349 2156
rect 338 2133 349 2136
rect 242 2113 301 2116
rect 346 2113 349 2133
rect 234 2093 245 2096
rect 218 2043 229 2046
rect 162 2013 165 2026
rect 178 2023 221 2026
rect 194 1983 197 2016
rect 218 2013 221 2023
rect 226 1946 229 2043
rect 242 1946 245 2093
rect 282 2013 285 2026
rect 298 2013 301 2113
rect 202 1933 205 1946
rect 218 1943 229 1946
rect 234 1943 245 1946
rect 130 1786 133 1816
rect 106 1783 133 1786
rect 66 1733 69 1766
rect 154 1703 157 1806
rect 170 1746 173 1866
rect 186 1856 189 1926
rect 178 1853 189 1856
rect 178 1813 181 1853
rect 218 1836 221 1943
rect 234 1863 237 1943
rect 242 1923 253 1926
rect 194 1833 221 1836
rect 194 1803 197 1833
rect 218 1813 221 1833
rect 242 1803 245 1923
rect 250 1913 253 1923
rect 250 1813 253 1826
rect 258 1813 261 1846
rect 266 1826 269 2006
rect 274 1933 277 2006
rect 298 2003 309 2006
rect 338 1976 341 2026
rect 354 2016 357 2163
rect 362 2123 365 2213
rect 386 2033 389 2136
rect 418 2083 421 2116
rect 434 2036 437 2216
rect 466 2176 469 2223
rect 490 2213 493 2226
rect 458 2173 469 2176
rect 458 2113 461 2173
rect 434 2033 445 2036
rect 346 1993 349 2016
rect 354 2013 397 2016
rect 354 1996 357 2013
rect 442 2003 445 2033
rect 458 2006 461 2036
rect 458 2003 469 2006
rect 354 1993 365 1996
rect 378 1993 397 1996
rect 450 1993 469 1996
rect 338 1973 349 1976
rect 346 1933 349 1973
rect 362 1946 365 1993
rect 354 1943 365 1946
rect 322 1913 325 1926
rect 354 1923 357 1943
rect 266 1823 285 1826
rect 266 1813 277 1816
rect 282 1806 285 1823
rect 290 1813 293 1826
rect 298 1813 301 1846
rect 354 1816 357 1916
rect 386 1826 389 1936
rect 386 1823 405 1826
rect 354 1813 389 1816
rect 266 1803 285 1806
rect 170 1743 189 1746
rect 66 1496 69 1646
rect 82 1526 85 1606
rect 130 1603 133 1616
rect 162 1613 165 1736
rect 186 1636 189 1743
rect 226 1733 229 1746
rect 266 1726 269 1803
rect 266 1723 277 1726
rect 170 1633 189 1636
rect 170 1606 173 1633
rect 210 1623 213 1706
rect 162 1603 173 1606
rect 82 1523 93 1526
rect 138 1523 141 1536
rect 162 1533 165 1603
rect 66 1493 77 1496
rect 74 1446 77 1493
rect 66 1443 77 1446
rect 66 1333 69 1443
rect 90 1336 93 1523
rect 138 1413 141 1426
rect 170 1413 173 1596
rect 178 1586 181 1606
rect 194 1603 205 1606
rect 178 1583 229 1586
rect 226 1533 229 1583
rect 234 1563 237 1606
rect 258 1596 261 1716
rect 274 1666 277 1723
rect 298 1716 301 1806
rect 250 1593 261 1596
rect 270 1663 277 1666
rect 290 1713 301 1716
rect 290 1666 293 1713
rect 290 1663 301 1666
rect 178 1413 181 1426
rect 82 1333 93 1336
rect 82 636 85 1333
rect 98 1133 101 1216
rect 114 1093 117 1346
rect 146 1313 149 1346
rect 154 1333 181 1336
rect 186 1333 189 1526
rect 218 1513 221 1526
rect 234 1506 237 1526
rect 230 1503 237 1506
rect 202 1403 205 1426
rect 218 1403 221 1446
rect 154 1323 157 1333
rect 162 1216 165 1326
rect 178 1313 181 1333
rect 202 1323 205 1346
rect 218 1333 221 1346
rect 210 1246 213 1306
rect 210 1243 221 1246
rect 138 1186 141 1216
rect 162 1213 169 1216
rect 130 1183 141 1186
rect 130 1143 133 1183
rect 130 1123 149 1126
rect 146 1113 149 1123
rect 154 1036 157 1206
rect 166 1136 169 1213
rect 178 1196 181 1206
rect 178 1193 197 1196
rect 178 1143 181 1193
rect 202 1186 205 1236
rect 194 1183 205 1186
rect 166 1133 173 1136
rect 150 1033 157 1036
rect 130 976 133 1016
rect 130 973 141 976
rect 114 923 117 936
rect 122 923 125 936
rect 138 933 141 973
rect 150 926 153 1033
rect 162 933 165 1026
rect 150 923 157 926
rect 130 813 133 826
rect 154 806 157 923
rect 170 816 173 1133
rect 194 1126 197 1183
rect 218 1156 221 1243
rect 230 1216 233 1503
rect 230 1213 237 1216
rect 242 1213 245 1536
rect 250 1506 253 1593
rect 270 1586 273 1663
rect 266 1583 273 1586
rect 266 1523 269 1583
rect 282 1533 285 1616
rect 298 1513 301 1663
rect 306 1526 309 1706
rect 322 1686 325 1806
rect 346 1733 365 1736
rect 322 1683 333 1686
rect 314 1533 317 1676
rect 330 1636 333 1683
rect 322 1633 333 1636
rect 306 1523 317 1526
rect 250 1503 261 1506
rect 258 1436 261 1503
rect 314 1496 317 1523
rect 250 1433 261 1436
rect 306 1493 317 1496
rect 250 1396 253 1433
rect 274 1413 277 1426
rect 306 1416 309 1493
rect 306 1413 317 1416
rect 250 1393 261 1396
rect 258 1346 261 1393
rect 250 1343 261 1346
rect 234 1193 237 1213
rect 242 1183 245 1206
rect 250 1196 253 1343
rect 258 1296 261 1326
rect 274 1316 277 1396
rect 282 1333 285 1346
rect 314 1336 317 1413
rect 322 1406 325 1633
rect 330 1556 333 1606
rect 346 1596 349 1733
rect 354 1706 357 1726
rect 362 1713 365 1733
rect 354 1703 365 1706
rect 362 1623 365 1703
rect 378 1636 381 1806
rect 386 1803 389 1813
rect 402 1736 405 1823
rect 426 1743 429 1936
rect 450 1816 453 1936
rect 474 1923 477 2156
rect 498 2133 501 2216
rect 522 2213 525 2326
rect 530 2323 533 2343
rect 626 2333 629 2346
rect 506 2113 509 2126
rect 514 2006 517 2206
rect 538 2143 541 2216
rect 626 2193 629 2216
rect 642 2203 645 2356
rect 658 2333 661 2533
rect 682 2523 685 2606
rect 730 2586 733 2606
rect 738 2593 741 2606
rect 754 2586 757 2616
rect 794 2613 797 2633
rect 818 2613 821 2626
rect 826 2613 829 2633
rect 850 2623 853 2756
rect 914 2753 941 2756
rect 882 2713 885 2746
rect 890 2703 893 2726
rect 914 2623 917 2656
rect 938 2616 941 2753
rect 946 2723 949 2816
rect 962 2813 965 2863
rect 954 2706 957 2786
rect 842 2613 869 2616
rect 914 2613 941 2616
rect 950 2703 957 2706
rect 730 2583 757 2586
rect 706 2506 709 2526
rect 698 2503 709 2506
rect 698 2456 701 2503
rect 698 2453 709 2456
rect 706 2433 709 2453
rect 722 2433 725 2526
rect 754 2523 757 2583
rect 842 2546 845 2613
rect 810 2543 845 2546
rect 674 2423 701 2426
rect 674 2403 677 2423
rect 690 2406 693 2416
rect 698 2413 701 2423
rect 666 2236 669 2346
rect 682 2343 685 2406
rect 690 2403 701 2406
rect 658 2233 669 2236
rect 546 2143 565 2146
rect 546 2016 549 2143
rect 562 2123 565 2136
rect 618 2113 621 2186
rect 530 2013 549 2016
rect 554 2013 597 2016
rect 514 2003 525 2006
rect 506 1993 525 1996
rect 442 1813 453 1816
rect 394 1733 405 1736
rect 394 1713 397 1733
rect 442 1696 445 1813
rect 442 1693 453 1696
rect 450 1676 453 1693
rect 442 1673 453 1676
rect 370 1613 373 1636
rect 378 1633 389 1636
rect 386 1613 389 1633
rect 410 1613 413 1636
rect 346 1593 357 1596
rect 330 1553 337 1556
rect 334 1496 337 1553
rect 354 1536 357 1593
rect 386 1563 389 1606
rect 346 1533 357 1536
rect 346 1513 349 1533
rect 394 1523 397 1536
rect 334 1493 349 1496
rect 346 1436 349 1493
rect 338 1433 349 1436
rect 338 1413 341 1433
rect 322 1403 341 1406
rect 306 1333 317 1336
rect 274 1313 285 1316
rect 258 1293 269 1296
rect 266 1236 269 1293
rect 258 1233 269 1236
rect 258 1213 261 1233
rect 250 1193 257 1196
rect 266 1193 269 1206
rect 210 1153 221 1156
rect 186 1123 197 1126
rect 186 1026 189 1123
rect 202 1106 205 1136
rect 198 1103 205 1106
rect 198 1046 201 1103
rect 198 1043 205 1046
rect 186 1023 197 1026
rect 194 983 197 1023
rect 202 963 205 1043
rect 210 936 213 1153
rect 218 1123 221 1136
rect 242 1133 245 1166
rect 254 1126 257 1193
rect 266 1133 269 1186
rect 226 1113 229 1126
rect 234 1096 237 1126
rect 218 1093 237 1096
rect 250 1123 257 1126
rect 218 1003 221 1093
rect 250 956 253 1123
rect 266 1013 269 1036
rect 274 1003 277 1016
rect 234 953 253 956
rect 186 933 229 936
rect 186 836 189 933
rect 186 833 197 836
rect 170 813 181 816
rect 194 813 197 833
rect 202 826 205 926
rect 202 823 213 826
rect 154 803 173 806
rect 178 786 181 813
rect 194 793 197 806
rect 202 786 205 816
rect 178 783 205 786
rect 202 766 205 783
rect 186 763 205 766
rect 186 636 189 763
rect 210 723 213 823
rect 218 803 221 826
rect 226 803 229 933
rect 234 906 237 953
rect 282 946 285 1313
rect 306 1303 309 1333
rect 338 1326 341 1403
rect 378 1343 381 1416
rect 394 1403 397 1416
rect 418 1403 421 1526
rect 394 1373 429 1376
rect 314 1323 341 1326
rect 314 1286 317 1323
rect 306 1283 317 1286
rect 306 1106 309 1283
rect 322 1176 325 1306
rect 330 1296 333 1316
rect 338 1313 341 1323
rect 354 1333 373 1336
rect 354 1303 357 1333
rect 394 1316 397 1373
rect 426 1333 429 1373
rect 434 1326 437 1616
rect 458 1603 461 1806
rect 498 1786 501 1806
rect 490 1783 501 1786
rect 466 1613 469 1746
rect 490 1736 493 1783
rect 506 1763 509 1936
rect 530 1813 533 2013
rect 554 1966 557 2013
rect 578 1993 597 1996
rect 546 1963 557 1966
rect 546 1923 549 1963
rect 618 1906 621 2106
rect 642 2013 645 2146
rect 658 2106 661 2233
rect 690 2203 693 2336
rect 698 2283 701 2403
rect 738 2386 741 2406
rect 786 2393 789 2406
rect 794 2403 797 2426
rect 818 2403 821 2526
rect 842 2523 845 2536
rect 850 2533 853 2546
rect 898 2523 901 2536
rect 906 2533 909 2606
rect 914 2523 917 2613
rect 938 2596 941 2606
rect 922 2593 941 2596
rect 922 2523 925 2593
rect 950 2576 953 2703
rect 962 2613 965 2726
rect 970 2703 973 2716
rect 978 2653 981 2826
rect 1002 2736 1005 2806
rect 1050 2756 1053 2873
rect 1074 2796 1077 2936
rect 1122 2923 1125 2946
rect 1146 2826 1149 3040
rect 1162 3026 1165 3040
rect 1162 3023 1173 3026
rect 1170 2956 1173 3023
rect 1162 2953 1173 2956
rect 1162 2933 1165 2953
rect 1138 2823 1149 2826
rect 1074 2793 1085 2796
rect 1050 2753 1061 2756
rect 1002 2733 1037 2736
rect 1010 2636 1013 2726
rect 994 2633 1013 2636
rect 994 2613 997 2633
rect 1042 2613 1045 2726
rect 1058 2723 1061 2753
rect 1066 2733 1069 2786
rect 1082 2706 1085 2793
rect 1066 2703 1085 2706
rect 1050 2603 1053 2626
rect 1066 2583 1069 2703
rect 946 2573 953 2576
rect 946 2556 949 2573
rect 942 2553 949 2556
rect 930 2513 933 2526
rect 942 2476 945 2553
rect 922 2473 945 2476
rect 922 2426 925 2473
rect 866 2413 869 2426
rect 922 2423 929 2426
rect 858 2403 869 2406
rect 738 2383 757 2386
rect 698 2186 701 2196
rect 666 2183 701 2186
rect 714 2183 717 2326
rect 730 2296 733 2326
rect 754 2313 757 2383
rect 802 2376 805 2396
rect 802 2373 813 2376
rect 786 2313 789 2346
rect 810 2316 813 2373
rect 850 2316 853 2356
rect 866 2333 869 2403
rect 802 2313 813 2316
rect 842 2313 853 2316
rect 802 2296 805 2313
rect 730 2293 741 2296
rect 738 2246 741 2293
rect 730 2243 741 2246
rect 794 2293 805 2296
rect 730 2223 733 2243
rect 666 2143 669 2183
rect 674 2143 717 2146
rect 674 2136 677 2143
rect 666 2133 677 2136
rect 682 2123 685 2136
rect 698 2133 709 2136
rect 658 2103 669 2106
rect 666 2036 669 2103
rect 658 2033 669 2036
rect 658 1923 661 2033
rect 666 1996 669 2016
rect 698 2013 701 2133
rect 706 2116 709 2126
rect 714 2123 717 2143
rect 722 2133 725 2216
rect 770 2183 773 2216
rect 794 2166 797 2293
rect 794 2163 805 2166
rect 802 2146 805 2163
rect 802 2143 813 2146
rect 818 2133 821 2286
rect 842 2216 845 2313
rect 858 2236 861 2326
rect 874 2323 877 2336
rect 890 2316 893 2406
rect 882 2313 893 2316
rect 858 2233 877 2236
rect 834 2213 845 2216
rect 866 2213 869 2226
rect 874 2213 877 2233
rect 882 2223 885 2313
rect 722 2116 725 2126
rect 706 2113 725 2116
rect 834 2103 837 2213
rect 666 1993 685 1996
rect 610 1903 621 1906
rect 538 1833 565 1836
rect 538 1813 541 1833
rect 554 1813 557 1826
rect 562 1816 565 1833
rect 562 1813 573 1816
rect 546 1753 549 1806
rect 578 1766 581 1856
rect 610 1826 613 1903
rect 570 1763 581 1766
rect 602 1823 613 1826
rect 490 1733 501 1736
rect 474 1603 477 1716
rect 498 1676 501 1733
rect 506 1696 509 1716
rect 506 1693 517 1696
rect 490 1673 501 1676
rect 490 1656 493 1673
rect 486 1653 493 1656
rect 486 1566 489 1653
rect 514 1646 517 1693
rect 506 1643 517 1646
rect 506 1623 509 1643
rect 530 1623 557 1626
rect 530 1613 533 1623
rect 538 1613 549 1616
rect 474 1563 489 1566
rect 506 1566 509 1606
rect 546 1603 557 1606
rect 506 1563 533 1566
rect 474 1436 477 1563
rect 530 1546 533 1563
rect 570 1556 573 1763
rect 602 1716 605 1823
rect 626 1796 629 1816
rect 618 1793 629 1796
rect 618 1736 621 1793
rect 618 1733 629 1736
rect 602 1713 621 1716
rect 618 1693 621 1713
rect 570 1553 589 1556
rect 530 1543 537 1546
rect 506 1523 509 1536
rect 534 1496 537 1543
rect 426 1323 437 1326
rect 458 1433 477 1436
rect 530 1493 537 1496
rect 426 1316 429 1323
rect 362 1296 365 1316
rect 330 1293 341 1296
rect 338 1226 341 1293
rect 330 1223 341 1226
rect 354 1293 365 1296
rect 386 1313 397 1316
rect 410 1313 429 1316
rect 354 1236 357 1293
rect 386 1256 389 1313
rect 386 1253 397 1256
rect 354 1233 389 1236
rect 330 1186 333 1223
rect 354 1213 357 1233
rect 362 1213 373 1216
rect 362 1206 365 1213
rect 346 1203 365 1206
rect 378 1196 381 1226
rect 370 1193 381 1196
rect 370 1186 373 1193
rect 330 1183 373 1186
rect 322 1173 341 1176
rect 330 1133 333 1166
rect 314 1123 333 1126
rect 306 1103 317 1106
rect 314 1046 317 1103
rect 314 1043 325 1046
rect 290 1023 293 1036
rect 322 1006 325 1043
rect 250 933 253 946
rect 274 943 285 946
rect 234 903 253 906
rect 218 733 229 736
rect 250 716 253 903
rect 274 896 277 943
rect 290 923 293 1006
rect 318 1003 325 1006
rect 318 916 321 1003
rect 330 923 333 986
rect 318 913 325 916
rect 242 713 253 716
rect 266 893 277 896
rect 242 646 245 713
rect 242 643 253 646
rect 82 633 93 636
rect 186 633 213 636
rect 90 533 93 633
rect 138 603 141 616
rect 202 613 205 626
rect 138 406 141 526
rect 194 426 197 526
rect 202 523 205 606
rect 210 586 213 633
rect 218 603 229 606
rect 234 603 237 626
rect 210 583 217 586
rect 214 506 217 583
rect 226 533 229 546
rect 242 516 245 536
rect 250 523 253 643
rect 266 633 269 893
rect 282 793 285 826
rect 314 773 317 806
rect 306 706 309 726
rect 298 703 309 706
rect 298 636 301 703
rect 298 633 309 636
rect 274 583 277 626
rect 306 616 309 633
rect 298 533 301 616
rect 306 613 313 616
rect 322 613 325 913
rect 338 906 341 1173
rect 346 1096 349 1136
rect 354 1113 357 1183
rect 346 1093 353 1096
rect 350 986 353 1093
rect 346 983 353 986
rect 362 1033 373 1036
rect 346 946 349 983
rect 346 943 353 946
rect 334 903 341 906
rect 334 816 337 903
rect 350 896 353 943
rect 362 923 365 1033
rect 378 1023 381 1186
rect 386 1133 389 1233
rect 394 1203 397 1253
rect 410 1116 413 1313
rect 458 1306 461 1433
rect 450 1303 461 1306
rect 450 1246 453 1303
rect 450 1243 457 1246
rect 418 1183 421 1206
rect 442 1166 445 1226
rect 454 1186 457 1243
rect 466 1186 469 1326
rect 474 1323 477 1426
rect 530 1413 533 1493
rect 546 1416 549 1526
rect 586 1436 589 1553
rect 594 1546 597 1606
rect 618 1603 621 1616
rect 594 1543 605 1546
rect 602 1446 605 1543
rect 626 1523 629 1733
rect 634 1716 637 1896
rect 682 1866 685 1993
rect 666 1863 685 1866
rect 658 1813 661 1826
rect 650 1736 653 1806
rect 642 1733 653 1736
rect 634 1713 641 1716
rect 650 1713 653 1726
rect 638 1526 641 1713
rect 666 1646 669 1863
rect 674 1753 677 1806
rect 690 1656 693 1846
rect 706 1676 709 1936
rect 714 1893 717 2006
rect 722 1923 725 2016
rect 738 1993 741 2006
rect 746 1996 749 2016
rect 754 2003 757 2016
rect 746 1993 757 1996
rect 762 1993 765 2006
rect 746 1933 749 1956
rect 754 1923 757 1993
rect 722 1686 725 1826
rect 738 1813 741 1826
rect 738 1696 741 1716
rect 754 1713 757 1806
rect 738 1693 753 1696
rect 722 1683 741 1686
rect 706 1673 717 1676
rect 662 1643 669 1646
rect 686 1653 693 1656
rect 634 1523 641 1526
rect 634 1503 637 1523
rect 570 1433 589 1436
rect 594 1443 605 1446
rect 546 1413 557 1416
rect 482 1316 485 1336
rect 530 1316 533 1406
rect 554 1403 557 1413
rect 554 1333 557 1386
rect 562 1323 565 1426
rect 570 1383 573 1433
rect 482 1313 493 1316
rect 530 1313 573 1316
rect 490 1236 493 1313
rect 578 1296 581 1426
rect 594 1423 597 1443
rect 586 1413 637 1416
rect 594 1403 605 1406
rect 570 1293 581 1296
rect 594 1296 597 1386
rect 650 1366 653 1526
rect 662 1456 665 1643
rect 674 1613 677 1636
rect 686 1606 689 1653
rect 698 1626 701 1646
rect 698 1623 705 1626
rect 674 1603 689 1606
rect 662 1453 669 1456
rect 666 1433 669 1453
rect 626 1363 653 1366
rect 594 1293 605 1296
rect 570 1246 573 1293
rect 570 1243 581 1246
rect 482 1233 493 1236
rect 482 1203 485 1233
rect 454 1183 461 1186
rect 466 1183 477 1186
rect 490 1183 493 1206
rect 506 1196 509 1216
rect 498 1193 509 1196
rect 458 1166 461 1183
rect 442 1163 453 1166
rect 458 1163 465 1166
rect 434 1126 437 1136
rect 442 1133 445 1156
rect 402 1113 413 1116
rect 426 1123 437 1126
rect 402 996 405 1113
rect 426 1006 429 1123
rect 450 1113 453 1163
rect 462 1106 465 1163
rect 458 1103 465 1106
rect 458 1053 461 1103
rect 474 1056 477 1183
rect 466 1053 477 1056
rect 418 1003 429 1006
rect 466 996 469 1053
rect 482 1013 485 1036
rect 490 1003 493 1136
rect 498 1126 501 1193
rect 498 1123 517 1126
rect 498 1096 501 1116
rect 498 1093 509 1096
rect 506 1026 509 1093
rect 498 1023 509 1026
rect 402 993 413 996
rect 466 993 493 996
rect 410 946 413 993
rect 370 933 373 946
rect 394 943 413 946
rect 394 936 397 943
rect 386 933 397 936
rect 330 813 337 816
rect 346 893 353 896
rect 346 836 349 893
rect 346 833 373 836
rect 330 716 333 813
rect 346 803 349 833
rect 354 796 357 816
rect 370 803 373 833
rect 386 823 389 933
rect 394 913 397 926
rect 402 906 405 936
rect 466 933 469 946
rect 402 903 413 906
rect 410 846 413 903
rect 402 843 413 846
rect 402 826 405 843
rect 402 823 421 826
rect 450 823 461 826
rect 466 823 469 836
rect 458 816 461 823
rect 346 793 357 796
rect 338 733 341 746
rect 346 723 349 793
rect 354 733 365 736
rect 370 733 373 746
rect 410 723 413 816
rect 458 813 469 816
rect 450 803 461 806
rect 466 803 469 813
rect 490 786 493 993
rect 498 913 501 1023
rect 506 923 509 1006
rect 522 976 525 1226
rect 546 1143 573 1146
rect 546 1133 549 1143
rect 554 1096 557 1136
rect 570 1133 573 1143
rect 578 1113 581 1243
rect 546 1093 557 1096
rect 546 1066 549 1093
rect 586 1086 589 1256
rect 602 1236 605 1293
rect 598 1233 605 1236
rect 598 1136 601 1233
rect 626 1226 629 1363
rect 666 1346 669 1366
rect 662 1343 669 1346
rect 626 1223 637 1226
rect 618 1203 621 1216
rect 634 1166 637 1223
rect 650 1203 653 1326
rect 662 1246 665 1343
rect 674 1253 677 1603
rect 690 1576 693 1596
rect 686 1573 693 1576
rect 686 1376 689 1573
rect 702 1566 705 1623
rect 714 1603 717 1673
rect 698 1563 705 1566
rect 698 1386 701 1563
rect 722 1556 725 1616
rect 730 1593 733 1606
rect 738 1566 741 1683
rect 750 1636 753 1693
rect 750 1633 757 1636
rect 714 1553 725 1556
rect 730 1563 741 1566
rect 746 1596 749 1606
rect 754 1603 757 1633
rect 762 1596 765 1936
rect 770 1923 773 1966
rect 794 1836 797 2036
rect 850 2016 853 2206
rect 898 2146 901 2336
rect 914 2246 917 2416
rect 926 2356 929 2423
rect 922 2353 929 2356
rect 922 2333 925 2353
rect 930 2313 933 2336
rect 910 2243 917 2246
rect 910 2166 913 2243
rect 910 2163 917 2166
rect 898 2143 905 2146
rect 866 2026 869 2136
rect 882 2133 893 2136
rect 874 2103 877 2126
rect 882 2113 893 2116
rect 866 2023 873 2026
rect 890 2023 893 2113
rect 902 2026 905 2143
rect 898 2023 905 2026
rect 842 2003 845 2016
rect 850 2013 861 2016
rect 858 2003 861 2013
rect 870 1976 873 2023
rect 898 2006 901 2023
rect 914 2013 917 2163
rect 866 1973 873 1976
rect 890 2003 901 2006
rect 866 1953 869 1973
rect 890 1946 893 2003
rect 866 1943 893 1946
rect 842 1843 845 1936
rect 858 1923 861 1936
rect 866 1923 869 1943
rect 794 1833 805 1836
rect 770 1786 773 1816
rect 778 1806 781 1826
rect 778 1803 789 1806
rect 770 1783 777 1786
rect 774 1666 777 1783
rect 746 1593 765 1596
rect 770 1663 777 1666
rect 714 1523 717 1553
rect 722 1533 725 1546
rect 730 1523 733 1563
rect 706 1393 709 1416
rect 698 1383 709 1386
rect 686 1373 693 1376
rect 690 1303 693 1373
rect 662 1243 669 1246
rect 666 1196 669 1243
rect 698 1213 701 1226
rect 706 1206 709 1383
rect 682 1203 709 1206
rect 594 1133 601 1136
rect 618 1163 637 1166
rect 650 1193 669 1196
rect 594 1113 597 1133
rect 618 1106 621 1163
rect 650 1133 653 1193
rect 706 1163 709 1203
rect 714 1146 717 1426
rect 730 1413 733 1466
rect 738 1406 741 1516
rect 722 1403 741 1406
rect 746 1386 749 1593
rect 770 1516 773 1663
rect 786 1646 789 1803
rect 778 1643 789 1646
rect 778 1596 781 1643
rect 802 1626 805 1833
rect 826 1793 829 1806
rect 826 1733 829 1746
rect 826 1673 829 1726
rect 834 1626 837 1816
rect 842 1803 845 1826
rect 858 1816 861 1836
rect 842 1713 845 1736
rect 850 1656 853 1816
rect 858 1813 865 1816
rect 874 1813 877 1936
rect 882 1923 885 1943
rect 890 1826 893 1936
rect 882 1823 893 1826
rect 862 1746 865 1813
rect 874 1763 877 1806
rect 862 1743 869 1746
rect 794 1623 805 1626
rect 826 1623 837 1626
rect 846 1653 853 1656
rect 778 1593 785 1596
rect 782 1526 785 1593
rect 754 1513 773 1516
rect 778 1523 785 1526
rect 754 1423 757 1513
rect 762 1503 773 1506
rect 778 1503 781 1523
rect 754 1393 757 1406
rect 762 1396 765 1416
rect 770 1403 773 1503
rect 762 1393 773 1396
rect 738 1383 749 1386
rect 722 1283 725 1336
rect 738 1256 741 1383
rect 762 1376 765 1393
rect 762 1373 769 1376
rect 722 1236 725 1256
rect 738 1253 749 1256
rect 722 1233 733 1236
rect 730 1156 733 1233
rect 698 1143 717 1146
rect 722 1153 733 1156
rect 666 1126 669 1136
rect 538 1063 549 1066
rect 554 1083 589 1086
rect 610 1103 621 1106
rect 538 986 541 1063
rect 538 983 545 986
rect 522 973 533 976
rect 498 793 501 816
rect 514 803 517 826
rect 490 783 501 786
rect 442 733 445 776
rect 458 733 461 746
rect 330 713 337 716
rect 310 546 313 613
rect 322 593 325 606
rect 334 566 337 713
rect 394 713 445 716
rect 394 636 397 713
rect 442 703 445 713
rect 482 656 485 726
rect 498 706 501 783
rect 522 723 525 826
rect 530 736 533 973
rect 542 916 545 983
rect 554 923 557 1083
rect 570 1023 573 1036
rect 610 973 613 1103
rect 578 933 581 966
rect 542 913 549 916
rect 538 746 541 816
rect 546 806 549 913
rect 562 813 565 826
rect 618 823 621 836
rect 546 803 565 806
rect 538 743 549 746
rect 530 733 541 736
rect 498 703 509 706
rect 538 703 541 733
rect 482 653 489 656
rect 346 623 349 636
rect 386 633 397 636
rect 330 563 337 566
rect 306 543 313 546
rect 306 526 309 543
rect 322 533 325 546
rect 306 523 325 526
rect 210 503 217 506
rect 234 513 245 516
rect 210 483 213 503
rect 234 446 237 513
rect 234 443 245 446
rect 162 423 189 426
rect 194 423 205 426
rect 242 423 245 443
rect 162 413 165 423
rect 186 416 189 423
rect 74 323 77 406
rect 138 403 173 406
rect 178 386 181 416
rect 186 413 197 416
rect 154 383 181 386
rect 90 333 93 346
rect 90 203 93 326
rect 106 323 109 336
rect 154 323 157 383
rect 186 376 189 406
rect 162 373 189 376
rect 162 306 165 373
rect 170 333 173 346
rect 154 303 165 306
rect 154 246 157 303
rect 154 243 165 246
rect 162 223 165 243
rect 170 226 173 236
rect 178 233 181 356
rect 194 313 197 413
rect 202 403 205 423
rect 170 223 189 226
rect 98 203 101 216
rect 170 206 173 216
rect 202 206 205 336
rect 234 213 237 406
rect 250 403 253 496
rect 322 493 325 516
rect 266 403 269 426
rect 322 353 325 426
rect 330 413 333 563
rect 346 546 349 616
rect 354 603 357 616
rect 386 586 389 633
rect 386 583 397 586
rect 338 543 349 546
rect 338 433 341 543
rect 346 423 349 536
rect 394 493 397 583
rect 418 506 421 606
rect 466 583 469 616
rect 486 596 489 653
rect 506 636 509 703
rect 482 593 489 596
rect 498 633 509 636
rect 482 576 485 593
rect 466 573 485 576
rect 410 503 421 506
rect 362 466 365 486
rect 362 463 373 466
rect 370 416 373 463
rect 362 413 373 416
rect 242 343 253 346
rect 290 333 309 336
rect 354 333 357 356
rect 362 333 365 413
rect 410 403 413 503
rect 434 446 437 566
rect 450 533 453 546
rect 458 533 461 566
rect 466 453 469 573
rect 434 443 445 446
rect 442 396 445 443
rect 434 393 445 396
rect 90 133 93 146
rect 114 123 117 206
rect 170 203 205 206
rect 186 116 189 126
rect 194 123 197 203
rect 202 116 205 136
rect 186 113 205 116
rect 186 0 189 113
rect 250 0 253 136
rect 266 133 269 326
rect 290 236 293 326
rect 298 313 301 326
rect 306 323 309 333
rect 338 323 365 326
rect 434 313 437 393
rect 458 383 461 416
rect 442 323 453 326
rect 482 313 485 516
rect 290 233 317 236
rect 498 233 501 633
rect 546 626 549 743
rect 570 733 573 776
rect 546 623 565 626
rect 514 593 517 616
rect 514 403 517 526
rect 522 483 525 616
rect 530 603 533 616
rect 546 603 557 606
rect 546 583 549 603
rect 538 523 541 536
rect 562 436 565 623
rect 570 593 573 606
rect 578 523 581 736
rect 594 723 597 746
rect 602 626 605 646
rect 594 623 605 626
rect 594 536 597 623
rect 610 546 613 816
rect 634 813 637 936
rect 642 933 645 1126
rect 650 1123 669 1126
rect 666 1113 669 1123
rect 698 1036 701 1143
rect 698 1033 717 1036
rect 658 976 661 1016
rect 658 973 669 976
rect 642 916 645 926
rect 650 923 653 946
rect 666 933 669 973
rect 690 963 693 1016
rect 714 993 717 1033
rect 714 933 717 976
rect 722 963 725 1153
rect 730 1116 733 1126
rect 738 1123 741 1136
rect 746 1123 749 1253
rect 754 1203 757 1366
rect 766 1236 769 1373
rect 762 1233 769 1236
rect 730 1113 757 1116
rect 762 1106 765 1233
rect 770 1193 773 1206
rect 770 1133 773 1146
rect 778 1116 781 1406
rect 786 1373 789 1406
rect 786 1203 789 1216
rect 794 1203 797 1623
rect 818 1593 821 1606
rect 826 1523 829 1623
rect 834 1533 837 1616
rect 846 1586 849 1653
rect 866 1646 869 1743
rect 842 1583 849 1586
rect 858 1643 869 1646
rect 842 1523 845 1583
rect 858 1576 861 1643
rect 866 1613 869 1626
rect 850 1573 861 1576
rect 850 1496 853 1573
rect 858 1533 861 1546
rect 866 1536 869 1576
rect 882 1553 885 1823
rect 898 1776 901 1796
rect 894 1773 901 1776
rect 894 1536 897 1773
rect 866 1533 877 1536
rect 842 1493 853 1496
rect 802 1396 805 1406
rect 810 1403 813 1416
rect 818 1403 821 1436
rect 826 1396 829 1406
rect 802 1393 829 1396
rect 802 1356 805 1376
rect 802 1353 809 1356
rect 806 1216 809 1353
rect 834 1336 837 1416
rect 842 1413 845 1493
rect 826 1333 837 1336
rect 842 1333 845 1346
rect 858 1336 861 1526
rect 874 1366 877 1533
rect 890 1533 897 1536
rect 890 1436 893 1533
rect 890 1433 901 1436
rect 866 1363 877 1366
rect 866 1343 869 1363
rect 858 1333 869 1336
rect 882 1326 885 1346
rect 802 1213 809 1216
rect 818 1213 821 1326
rect 834 1323 885 1326
rect 842 1313 853 1316
rect 826 1266 829 1286
rect 826 1263 833 1266
rect 802 1196 805 1213
rect 830 1206 833 1263
rect 754 1103 765 1106
rect 770 1113 781 1116
rect 786 1193 805 1196
rect 826 1203 833 1206
rect 754 1013 757 1103
rect 762 1003 765 1016
rect 770 1013 773 1113
rect 786 956 789 1193
rect 794 1013 797 1036
rect 802 973 805 1136
rect 826 1086 829 1203
rect 842 1156 845 1313
rect 882 1306 885 1323
rect 874 1303 885 1306
rect 874 1246 877 1303
rect 874 1243 885 1246
rect 842 1153 849 1156
rect 834 1123 837 1146
rect 822 1083 829 1086
rect 810 993 813 1036
rect 786 953 797 956
rect 642 913 669 916
rect 754 816 757 826
rect 738 813 757 816
rect 762 813 765 926
rect 626 773 629 806
rect 658 766 661 806
rect 650 763 661 766
rect 618 723 621 746
rect 650 733 653 763
rect 618 703 621 716
rect 674 646 677 796
rect 738 793 741 806
rect 754 803 757 813
rect 794 793 797 953
rect 810 806 813 946
rect 822 886 825 1083
rect 834 893 837 1096
rect 846 1076 849 1153
rect 866 1126 869 1226
rect 874 1136 877 1206
rect 882 1203 885 1243
rect 890 1203 893 1416
rect 898 1276 901 1433
rect 906 1283 909 2006
rect 922 1963 925 2236
rect 938 2216 941 2416
rect 946 2323 949 2436
rect 954 2306 957 2566
rect 1098 2536 1101 2806
rect 1138 2756 1141 2823
rect 1138 2753 1149 2756
rect 1106 2703 1109 2726
rect 1130 2656 1133 2736
rect 1146 2706 1149 2753
rect 1162 2733 1165 2816
rect 1178 2723 1181 2926
rect 1186 2813 1189 2826
rect 1202 2706 1205 3006
rect 1274 2976 1277 3040
rect 1274 2973 1285 2976
rect 1218 2906 1221 2936
rect 1234 2933 1237 2946
rect 1242 2923 1245 2936
rect 1218 2903 1229 2906
rect 1210 2783 1213 2806
rect 1226 2756 1229 2903
rect 1250 2823 1253 2936
rect 1258 2933 1261 2966
rect 1282 2926 1285 2973
rect 1274 2923 1285 2926
rect 1258 2823 1261 2836
rect 1266 2813 1269 2826
rect 1146 2703 1157 2706
rect 1130 2653 1137 2656
rect 1106 2613 1109 2626
rect 1134 2596 1137 2653
rect 1154 2636 1157 2703
rect 1146 2633 1157 2636
rect 1194 2703 1205 2706
rect 1218 2753 1229 2756
rect 1146 2613 1149 2633
rect 1130 2593 1137 2596
rect 1130 2566 1133 2593
rect 1194 2586 1197 2703
rect 1126 2563 1133 2566
rect 962 2413 965 2526
rect 970 2403 973 2426
rect 978 2333 981 2516
rect 994 2473 997 2536
rect 1010 2413 1013 2536
rect 1018 2513 1021 2526
rect 1034 2503 1037 2526
rect 1058 2486 1061 2536
rect 1042 2483 1061 2486
rect 986 2383 989 2406
rect 994 2326 997 2406
rect 1042 2366 1045 2483
rect 1066 2376 1069 2536
rect 1090 2533 1101 2536
rect 1066 2373 1077 2376
rect 950 2303 957 2306
rect 962 2323 997 2326
rect 950 2236 953 2303
rect 950 2233 957 2236
rect 938 2213 945 2216
rect 930 1946 933 2206
rect 942 2026 945 2213
rect 954 2033 957 2233
rect 962 2203 965 2323
rect 970 2213 973 2226
rect 962 2073 965 2126
rect 970 2103 973 2136
rect 978 2046 981 2316
rect 962 2043 981 2046
rect 922 1943 933 1946
rect 938 2023 945 2026
rect 922 1846 925 1943
rect 922 1843 933 1846
rect 914 1573 917 1736
rect 922 1716 925 1776
rect 930 1736 933 1843
rect 938 1793 941 2023
rect 962 2013 965 2043
rect 986 2026 989 2136
rect 982 2023 989 2026
rect 946 2003 957 2006
rect 962 1986 965 2006
rect 954 1983 965 1986
rect 946 1933 949 1946
rect 954 1836 957 1983
rect 962 1923 965 1966
rect 970 1906 973 2006
rect 982 1956 985 2023
rect 994 2003 997 2246
rect 1002 2233 1005 2326
rect 1010 2226 1013 2366
rect 1042 2363 1057 2366
rect 1026 2333 1029 2346
rect 1034 2323 1037 2336
rect 1018 2246 1021 2296
rect 1018 2243 1029 2246
rect 1010 2223 1017 2226
rect 1002 1996 1005 2206
rect 1014 2066 1017 2223
rect 1026 2083 1029 2243
rect 1042 2133 1045 2326
rect 1054 2296 1057 2363
rect 1054 2293 1061 2296
rect 1058 2153 1061 2293
rect 1074 2236 1077 2373
rect 1090 2346 1093 2436
rect 1090 2343 1101 2346
rect 1066 2233 1077 2236
rect 1014 2063 1021 2066
rect 994 1993 1005 1996
rect 982 1953 989 1956
rect 950 1833 957 1836
rect 966 1903 973 1906
rect 950 1746 953 1833
rect 966 1826 969 1903
rect 962 1823 969 1826
rect 950 1743 957 1746
rect 962 1743 965 1823
rect 930 1733 941 1736
rect 922 1713 929 1716
rect 926 1626 929 1713
rect 922 1623 929 1626
rect 922 1546 925 1623
rect 930 1553 933 1606
rect 922 1543 933 1546
rect 930 1476 933 1543
rect 938 1486 941 1733
rect 946 1603 949 1726
rect 954 1643 957 1743
rect 962 1723 965 1736
rect 970 1706 973 1816
rect 978 1803 981 1936
rect 986 1833 989 1953
rect 994 1923 997 1993
rect 1018 1986 1021 2063
rect 1042 2013 1045 2126
rect 1058 2116 1061 2136
rect 1054 2113 1061 2116
rect 1054 2046 1057 2113
rect 1054 2043 1061 2046
rect 1034 1993 1037 2006
rect 1010 1983 1021 1986
rect 1010 1966 1013 1983
rect 1006 1963 1013 1966
rect 1006 1906 1009 1963
rect 1050 1956 1053 2026
rect 1018 1953 1053 1956
rect 1018 1933 1021 1953
rect 1034 1933 1037 1946
rect 1018 1923 1037 1926
rect 1018 1913 1021 1923
rect 1034 1913 1037 1923
rect 1006 1903 1013 1906
rect 986 1823 1005 1826
rect 986 1786 989 1816
rect 962 1703 973 1706
rect 982 1783 989 1786
rect 962 1613 965 1703
rect 954 1603 965 1606
rect 970 1603 973 1646
rect 982 1626 985 1783
rect 1010 1773 1013 1903
rect 1058 1896 1061 2043
rect 1066 1976 1069 2233
rect 1098 2223 1101 2343
rect 1106 2323 1109 2536
rect 1114 2513 1117 2526
rect 1126 2496 1129 2563
rect 1122 2493 1129 2496
rect 1122 2376 1125 2493
rect 1122 2373 1133 2376
rect 1130 2353 1133 2373
rect 1082 2196 1085 2216
rect 1074 2193 1085 2196
rect 1074 2133 1077 2193
rect 1082 2093 1085 2126
rect 1090 2016 1093 2136
rect 1098 2133 1101 2206
rect 1074 1993 1077 2016
rect 1090 2013 1097 2016
rect 1066 1973 1073 1976
rect 1050 1893 1061 1896
rect 1018 1766 1021 1836
rect 1050 1826 1053 1893
rect 1070 1886 1073 1973
rect 1082 1903 1085 2006
rect 1094 1896 1097 2013
rect 1114 1996 1117 2336
rect 1122 2333 1125 2346
rect 1138 2146 1141 2576
rect 1170 2533 1173 2586
rect 1194 2583 1205 2586
rect 1202 2563 1205 2583
rect 1218 2563 1221 2753
rect 1234 2733 1245 2736
rect 1274 2726 1277 2923
rect 1282 2816 1285 2826
rect 1290 2823 1293 2836
rect 1306 2816 1309 3040
rect 1386 3026 1389 3040
rect 1378 3023 1389 3026
rect 1378 2956 1381 3023
rect 1378 2953 1385 2956
rect 1314 2923 1317 2936
rect 1338 2906 1341 2926
rect 1346 2913 1349 2936
rect 1330 2903 1341 2906
rect 1330 2836 1333 2903
rect 1330 2833 1341 2836
rect 1282 2813 1293 2816
rect 1306 2813 1325 2816
rect 1306 2743 1309 2806
rect 1322 2756 1325 2813
rect 1338 2803 1341 2833
rect 1354 2816 1357 2936
rect 1362 2916 1365 2936
rect 1362 2913 1373 2916
rect 1370 2846 1373 2913
rect 1346 2813 1357 2816
rect 1362 2843 1373 2846
rect 1314 2753 1325 2756
rect 1234 2723 1253 2726
rect 1274 2723 1285 2726
rect 1234 2643 1237 2723
rect 1242 2636 1245 2716
rect 1250 2713 1269 2716
rect 1250 2703 1253 2713
rect 1258 2656 1261 2706
rect 1258 2653 1265 2656
rect 1226 2633 1245 2636
rect 1226 2613 1229 2633
rect 1234 2603 1237 2626
rect 1242 2543 1245 2616
rect 1250 2603 1253 2646
rect 1262 2606 1265 2653
rect 1282 2646 1285 2723
rect 1314 2656 1317 2753
rect 1322 2723 1325 2736
rect 1346 2706 1349 2813
rect 1354 2793 1357 2806
rect 1362 2803 1365 2843
rect 1382 2826 1385 2953
rect 1378 2823 1385 2826
rect 1362 2713 1365 2756
rect 1346 2703 1365 2706
rect 1370 2703 1373 2726
rect 1362 2656 1365 2703
rect 1314 2653 1333 2656
rect 1362 2653 1369 2656
rect 1258 2603 1265 2606
rect 1274 2643 1285 2646
rect 1258 2586 1261 2603
rect 1274 2596 1277 2643
rect 1274 2593 1281 2596
rect 1258 2583 1269 2586
rect 1258 2536 1261 2583
rect 1218 2523 1221 2536
rect 1242 2533 1261 2536
rect 1266 2533 1269 2566
rect 1242 2476 1245 2533
rect 1154 2333 1157 2406
rect 1162 2356 1165 2476
rect 1234 2473 1245 2476
rect 1186 2413 1189 2426
rect 1210 2423 1213 2436
rect 1170 2383 1173 2406
rect 1186 2403 1197 2406
rect 1234 2396 1237 2473
rect 1250 2403 1253 2526
rect 1258 2423 1261 2526
rect 1266 2413 1269 2526
rect 1278 2516 1281 2593
rect 1298 2556 1301 2606
rect 1298 2553 1325 2556
rect 1290 2533 1301 2536
rect 1306 2523 1309 2546
rect 1314 2523 1317 2536
rect 1278 2513 1285 2516
rect 1282 2426 1285 2513
rect 1322 2506 1325 2553
rect 1274 2423 1285 2426
rect 1314 2503 1325 2506
rect 1234 2393 1253 2396
rect 1162 2353 1181 2356
rect 1130 2143 1141 2146
rect 1130 2016 1133 2143
rect 1146 2123 1149 2136
rect 1154 2113 1157 2316
rect 1178 2226 1181 2353
rect 1170 2223 1181 2226
rect 1170 2106 1173 2223
rect 1202 2216 1205 2386
rect 1242 2333 1245 2356
rect 1242 2306 1245 2326
rect 1250 2323 1253 2393
rect 1274 2363 1277 2423
rect 1290 2383 1293 2406
rect 1314 2396 1317 2503
rect 1330 2403 1333 2653
rect 1346 2603 1349 2616
rect 1366 2566 1369 2653
rect 1362 2563 1369 2566
rect 1338 2516 1341 2556
rect 1362 2543 1365 2563
rect 1378 2536 1381 2823
rect 1394 2733 1397 2956
rect 1402 2916 1405 3026
rect 1418 2976 1421 3040
rect 1410 2973 1429 2976
rect 1410 2933 1413 2973
rect 1402 2913 1413 2916
rect 1410 2846 1413 2913
rect 1426 2906 1429 2973
rect 1434 2953 1437 3040
rect 1450 2966 1453 3040
rect 1466 3023 1469 3040
rect 1482 3003 1485 3040
rect 1506 2966 1509 3040
rect 1578 2976 1581 3040
rect 1530 2973 1581 2976
rect 1450 2963 1469 2966
rect 1506 2963 1513 2966
rect 1442 2933 1445 2946
rect 1426 2903 1445 2906
rect 1402 2843 1413 2846
rect 1354 2533 1381 2536
rect 1338 2513 1349 2516
rect 1346 2446 1349 2513
rect 1338 2443 1349 2446
rect 1338 2413 1341 2443
rect 1314 2393 1325 2396
rect 1234 2303 1245 2306
rect 1202 2213 1213 2216
rect 1186 2203 1197 2206
rect 1162 2103 1173 2106
rect 1130 2013 1137 2016
rect 1146 2013 1149 2096
rect 1162 2036 1165 2103
rect 1162 2033 1173 2036
rect 1114 1993 1125 1996
rect 1106 1933 1109 1986
rect 1122 1946 1125 1993
rect 1114 1943 1125 1946
rect 1134 1946 1137 2013
rect 1146 1953 1149 1986
rect 1134 1943 1141 1946
rect 1154 1943 1157 2026
rect 1034 1823 1053 1826
rect 1066 1883 1073 1886
rect 1090 1893 1097 1896
rect 1034 1786 1037 1823
rect 1058 1806 1061 1816
rect 1042 1803 1061 1806
rect 1034 1783 1045 1786
rect 994 1763 1021 1766
rect 982 1623 989 1626
rect 962 1596 965 1603
rect 978 1596 981 1606
rect 986 1603 989 1623
rect 962 1593 981 1596
rect 994 1566 997 1763
rect 986 1563 997 1566
rect 946 1523 949 1536
rect 986 1516 989 1563
rect 1002 1523 1005 1736
rect 1010 1573 1013 1746
rect 1018 1523 1021 1716
rect 1042 1706 1045 1783
rect 1066 1733 1069 1883
rect 1074 1706 1077 1816
rect 1090 1766 1093 1893
rect 1106 1823 1109 1856
rect 1114 1833 1117 1943
rect 1122 1903 1125 1926
rect 1138 1826 1141 1943
rect 1170 1936 1173 2033
rect 1186 2016 1189 2156
rect 1194 2143 1197 2203
rect 1210 2046 1213 2213
rect 1234 2196 1237 2303
rect 1258 2203 1261 2346
rect 1322 2246 1325 2393
rect 1338 2313 1341 2326
rect 1346 2256 1349 2426
rect 1362 2403 1365 2416
rect 1370 2413 1373 2436
rect 1354 2316 1357 2346
rect 1378 2323 1381 2533
rect 1386 2723 1397 2726
rect 1386 2523 1389 2723
rect 1394 2683 1397 2716
rect 1394 2613 1397 2636
rect 1394 2583 1397 2606
rect 1394 2533 1397 2566
rect 1386 2396 1389 2416
rect 1386 2393 1393 2396
rect 1390 2336 1393 2393
rect 1386 2333 1393 2336
rect 1386 2316 1389 2333
rect 1354 2313 1389 2316
rect 1346 2253 1397 2256
rect 1322 2243 1373 2246
rect 1266 2213 1269 2226
rect 1290 2196 1293 2216
rect 1234 2193 1245 2196
rect 1242 2133 1245 2193
rect 1282 2193 1293 2196
rect 1282 2136 1285 2193
rect 1306 2176 1309 2216
rect 1306 2173 1313 2176
rect 1282 2133 1301 2136
rect 1298 2123 1301 2133
rect 1130 1823 1141 1826
rect 1162 1933 1173 1936
rect 1182 2013 1189 2016
rect 1202 2043 1213 2046
rect 1106 1803 1109 1816
rect 1130 1766 1133 1823
rect 1146 1796 1149 1816
rect 1146 1793 1153 1796
rect 1090 1763 1117 1766
rect 1130 1763 1141 1766
rect 1082 1733 1085 1746
rect 1034 1703 1045 1706
rect 1066 1703 1077 1706
rect 1034 1666 1037 1703
rect 1034 1663 1045 1666
rect 1026 1603 1029 1616
rect 1034 1533 1037 1546
rect 962 1503 965 1516
rect 986 1513 997 1516
rect 938 1483 949 1486
rect 930 1473 941 1476
rect 898 1273 905 1276
rect 902 1216 905 1273
rect 902 1213 909 1216
rect 874 1133 893 1136
rect 898 1133 901 1196
rect 866 1123 885 1126
rect 890 1123 893 1133
rect 842 1073 849 1076
rect 842 923 845 1073
rect 850 1003 853 1056
rect 874 1013 877 1046
rect 882 1026 885 1116
rect 906 1093 909 1213
rect 914 1126 917 1456
rect 922 1203 925 1406
rect 930 1403 933 1473
rect 946 1346 949 1483
rect 938 1343 949 1346
rect 938 1336 941 1343
rect 930 1333 941 1336
rect 930 1296 933 1333
rect 938 1313 941 1326
rect 946 1316 949 1336
rect 954 1323 957 1346
rect 962 1333 965 1496
rect 994 1456 997 1513
rect 994 1453 1037 1456
rect 978 1423 997 1426
rect 970 1393 973 1416
rect 986 1386 989 1406
rect 982 1383 989 1386
rect 970 1316 973 1326
rect 946 1313 973 1316
rect 930 1293 941 1296
rect 938 1246 941 1293
rect 930 1243 941 1246
rect 930 1223 933 1243
rect 962 1213 965 1256
rect 982 1246 985 1383
rect 982 1243 989 1246
rect 970 1133 973 1216
rect 978 1126 981 1226
rect 914 1123 933 1126
rect 882 1023 909 1026
rect 866 996 869 1006
rect 882 1003 885 1023
rect 890 996 893 1006
rect 866 993 893 996
rect 898 976 901 1016
rect 906 993 909 1023
rect 874 973 901 976
rect 874 933 877 973
rect 906 956 909 976
rect 930 956 933 1123
rect 970 1123 981 1126
rect 890 953 909 956
rect 914 953 933 956
rect 882 903 885 926
rect 822 883 829 886
rect 818 813 821 836
rect 826 826 829 883
rect 826 823 837 826
rect 842 823 845 836
rect 826 806 829 816
rect 810 803 829 806
rect 738 716 741 746
rect 802 733 805 766
rect 826 753 829 803
rect 834 786 837 823
rect 842 803 845 816
rect 834 783 845 786
rect 802 723 813 726
rect 810 716 813 723
rect 818 716 821 736
rect 842 726 845 783
rect 882 726 885 756
rect 890 743 893 953
rect 898 923 901 936
rect 914 826 917 953
rect 954 926 957 1116
rect 970 1003 973 1123
rect 986 1106 989 1243
rect 994 1133 997 1423
rect 1002 1333 1005 1406
rect 1010 1403 1013 1416
rect 982 1103 989 1106
rect 982 1036 985 1103
rect 982 1033 989 1036
rect 970 933 973 946
rect 978 936 981 1016
rect 986 983 989 1033
rect 994 1023 997 1126
rect 978 933 989 936
rect 954 923 973 926
rect 914 823 933 826
rect 914 733 917 816
rect 930 766 933 823
rect 970 813 973 923
rect 994 886 997 926
rect 986 883 997 886
rect 986 836 989 883
rect 986 833 997 836
rect 994 813 997 833
rect 1002 796 1005 1306
rect 922 763 933 766
rect 986 793 1005 796
rect 1010 793 1013 1356
rect 1018 1096 1021 1436
rect 1034 1353 1037 1453
rect 1026 1326 1029 1346
rect 1026 1323 1033 1326
rect 1030 1236 1033 1323
rect 1026 1233 1033 1236
rect 1026 1123 1029 1233
rect 1042 1216 1045 1663
rect 1066 1636 1069 1703
rect 1066 1633 1077 1636
rect 1074 1613 1077 1633
rect 1090 1626 1093 1756
rect 1106 1716 1109 1736
rect 1102 1713 1109 1716
rect 1102 1646 1105 1713
rect 1102 1643 1109 1646
rect 1082 1623 1093 1626
rect 1082 1606 1085 1623
rect 1066 1603 1085 1606
rect 1090 1603 1093 1616
rect 1050 1533 1061 1536
rect 1066 1523 1069 1603
rect 1074 1543 1085 1546
rect 1058 1496 1061 1516
rect 1058 1493 1065 1496
rect 1050 1376 1053 1486
rect 1062 1386 1065 1493
rect 1082 1436 1085 1536
rect 1098 1503 1101 1626
rect 1106 1493 1109 1643
rect 1114 1533 1117 1763
rect 1122 1723 1125 1736
rect 1130 1723 1133 1746
rect 1138 1743 1141 1763
rect 1150 1736 1153 1793
rect 1146 1733 1153 1736
rect 1122 1586 1125 1646
rect 1146 1613 1149 1733
rect 1162 1646 1165 1933
rect 1182 1926 1185 2013
rect 1194 1933 1197 2006
rect 1182 1923 1189 1926
rect 1186 1866 1189 1923
rect 1178 1863 1189 1866
rect 1178 1786 1181 1863
rect 1178 1783 1189 1786
rect 1154 1643 1165 1646
rect 1154 1613 1165 1616
rect 1130 1603 1141 1606
rect 1154 1593 1157 1606
rect 1162 1603 1165 1613
rect 1170 1586 1173 1766
rect 1122 1583 1133 1586
rect 1130 1486 1133 1583
rect 1166 1583 1173 1586
rect 1154 1523 1157 1556
rect 1122 1483 1133 1486
rect 1082 1433 1089 1436
rect 1062 1383 1069 1386
rect 1050 1373 1057 1376
rect 1034 1213 1045 1216
rect 1018 1093 1025 1096
rect 1022 946 1025 1093
rect 1034 946 1037 1213
rect 1054 1206 1057 1373
rect 1042 1186 1045 1206
rect 1054 1203 1061 1206
rect 1042 1183 1049 1186
rect 1046 1106 1049 1183
rect 1042 1103 1049 1106
rect 1042 1083 1045 1103
rect 1058 1086 1061 1203
rect 1066 1176 1069 1383
rect 1074 1313 1077 1426
rect 1086 1356 1089 1433
rect 1098 1403 1101 1416
rect 1082 1353 1089 1356
rect 1074 1193 1077 1216
rect 1066 1173 1073 1176
rect 1054 1083 1061 1086
rect 1042 1003 1045 1016
rect 1054 956 1057 1083
rect 1070 1076 1073 1173
rect 1066 1073 1073 1076
rect 1054 953 1061 956
rect 1022 943 1029 946
rect 1034 943 1045 946
rect 1018 923 1021 936
rect 1026 836 1029 943
rect 1018 833 1029 836
rect 706 703 709 716
rect 738 713 749 716
rect 810 713 821 716
rect 826 723 845 726
rect 674 643 701 646
rect 618 613 621 626
rect 674 613 677 636
rect 658 563 661 606
rect 610 543 617 546
rect 594 533 605 536
rect 594 476 597 516
rect 586 473 597 476
rect 562 433 573 436
rect 530 423 557 426
rect 530 413 533 423
rect 538 346 541 416
rect 554 413 557 423
rect 554 383 557 406
rect 570 356 573 433
rect 586 396 589 473
rect 602 403 605 533
rect 614 456 617 543
rect 626 506 629 526
rect 642 523 645 536
rect 650 533 653 546
rect 674 516 677 606
rect 666 513 677 516
rect 626 503 637 506
rect 610 453 617 456
rect 610 416 613 453
rect 618 423 621 436
rect 610 413 621 416
rect 634 406 637 503
rect 666 426 669 513
rect 698 506 701 643
rect 730 623 733 706
rect 746 636 749 713
rect 826 706 829 723
rect 874 716 877 726
rect 882 723 909 726
rect 874 713 901 716
rect 738 633 749 636
rect 730 563 733 606
rect 738 603 741 633
rect 818 623 821 706
rect 826 703 845 706
rect 842 616 845 703
rect 906 633 909 723
rect 922 676 925 763
rect 986 746 989 793
rect 1018 763 1021 833
rect 1034 803 1037 816
rect 1042 786 1045 943
rect 1034 783 1045 786
rect 938 696 941 746
rect 962 733 965 746
rect 986 743 993 746
rect 990 696 993 743
rect 938 693 949 696
rect 914 673 925 676
rect 746 576 749 616
rect 826 613 845 616
rect 746 573 757 576
rect 722 533 741 536
rect 690 503 701 506
rect 666 423 677 426
rect 626 403 637 406
rect 586 393 597 396
rect 522 343 541 346
rect 562 353 573 356
rect 522 236 525 343
rect 562 336 565 353
rect 546 333 573 336
rect 522 233 541 236
rect 282 213 309 216
rect 314 203 317 233
rect 346 223 381 226
rect 362 213 381 216
rect 378 193 381 206
rect 274 113 277 126
rect 322 0 325 136
rect 354 113 357 126
rect 370 103 373 116
rect 378 103 381 116
rect 386 16 389 206
rect 434 173 437 206
rect 458 193 461 216
rect 514 183 517 216
rect 538 193 541 233
rect 546 203 549 326
rect 554 313 557 326
rect 570 323 573 333
rect 594 303 597 393
rect 570 166 573 206
rect 522 163 573 166
rect 418 123 429 126
rect 386 13 429 16
rect 426 0 429 13
rect 442 0 445 136
rect 474 133 477 146
rect 522 123 525 163
rect 578 156 581 236
rect 610 206 613 336
rect 626 326 629 403
rect 626 323 653 326
rect 650 303 653 316
rect 658 313 661 406
rect 674 403 677 423
rect 682 333 685 346
rect 690 323 693 503
rect 730 483 733 526
rect 754 476 757 573
rect 778 513 781 536
rect 786 533 789 556
rect 802 513 805 536
rect 826 496 829 613
rect 914 586 917 673
rect 922 646 925 666
rect 922 643 933 646
rect 910 583 917 586
rect 746 473 757 476
rect 818 493 829 496
rect 706 413 709 456
rect 698 343 725 346
rect 698 323 701 343
rect 714 326 717 336
rect 722 333 725 343
rect 706 323 717 326
rect 706 316 709 323
rect 690 313 709 316
rect 618 223 621 246
rect 610 203 621 206
rect 562 153 581 156
rect 562 123 565 153
rect 578 133 581 146
rect 626 123 629 156
rect 682 123 685 216
rect 690 203 693 313
rect 690 116 693 126
rect 698 123 701 196
rect 714 133 717 156
rect 722 116 725 326
rect 730 303 733 426
rect 746 323 749 473
rect 818 426 821 493
rect 794 406 797 426
rect 818 423 829 426
rect 762 383 765 406
rect 770 336 773 406
rect 790 403 797 406
rect 790 346 793 403
rect 802 393 805 406
rect 810 383 813 406
rect 762 333 773 336
rect 786 343 793 346
rect 786 303 789 343
rect 802 273 805 336
rect 810 333 813 346
rect 826 323 829 423
rect 842 336 845 536
rect 866 513 869 526
rect 910 516 913 583
rect 930 576 933 643
rect 922 573 933 576
rect 922 523 925 573
rect 946 556 949 693
rect 986 693 993 696
rect 970 613 973 626
rect 946 553 957 556
rect 930 533 933 546
rect 910 513 917 516
rect 858 403 861 486
rect 866 423 909 426
rect 834 333 845 336
rect 866 333 869 423
rect 898 396 901 416
rect 890 393 901 396
rect 890 346 893 393
rect 890 343 901 346
rect 754 223 773 226
rect 754 213 757 223
rect 762 213 773 216
rect 754 153 757 206
rect 786 193 789 216
rect 794 133 797 176
rect 834 173 837 333
rect 874 246 877 326
rect 882 256 885 326
rect 898 313 901 343
rect 882 253 893 256
rect 874 243 885 246
rect 890 236 893 253
rect 882 233 893 236
rect 842 213 845 226
rect 690 113 725 116
rect 746 113 749 126
rect 842 123 845 206
rect 874 63 877 156
rect 882 143 885 233
rect 898 203 909 206
rect 914 196 917 513
rect 930 493 933 526
rect 930 393 933 406
rect 954 376 957 553
rect 938 373 957 376
rect 922 333 925 346
rect 922 203 925 246
rect 906 193 917 196
rect 906 153 909 193
rect 938 143 941 373
rect 962 323 965 346
rect 978 236 981 636
rect 986 583 989 693
rect 1002 676 1005 726
rect 1002 673 1013 676
rect 1010 626 1013 673
rect 1034 656 1037 783
rect 1050 663 1053 936
rect 1058 823 1061 953
rect 1066 916 1069 1073
rect 1074 1023 1077 1046
rect 1082 996 1085 1353
rect 1090 1286 1093 1336
rect 1098 1313 1101 1326
rect 1090 1283 1101 1286
rect 1090 1193 1093 1216
rect 1098 1213 1101 1283
rect 1074 993 1085 996
rect 1074 933 1077 993
rect 1082 933 1085 976
rect 1066 913 1077 916
rect 1074 836 1077 913
rect 1066 833 1077 836
rect 1066 806 1069 833
rect 1090 816 1093 1126
rect 1106 1093 1109 1226
rect 1098 1003 1101 1086
rect 1106 996 1109 1016
rect 1098 993 1109 996
rect 1098 933 1101 993
rect 1106 903 1109 926
rect 1062 803 1069 806
rect 1082 813 1093 816
rect 1106 816 1109 896
rect 1106 813 1113 816
rect 1034 653 1045 656
rect 1002 623 1013 626
rect 1002 603 1005 623
rect 1002 513 1005 536
rect 1010 533 1021 536
rect 1026 513 1029 546
rect 1042 533 1045 653
rect 1062 646 1065 803
rect 1058 643 1065 646
rect 1058 596 1061 643
rect 1074 603 1077 796
rect 1082 756 1085 813
rect 1090 803 1101 806
rect 1082 753 1093 756
rect 1082 733 1085 746
rect 1090 646 1093 753
rect 1098 713 1101 803
rect 1110 766 1113 813
rect 1106 763 1113 766
rect 1122 766 1125 1483
rect 1166 1476 1169 1583
rect 1166 1473 1173 1476
rect 1170 1453 1173 1473
rect 1178 1426 1181 1736
rect 1186 1593 1189 1783
rect 1194 1483 1197 1856
rect 1202 1763 1205 2043
rect 1210 1906 1213 2026
rect 1226 2003 1229 2016
rect 1242 2003 1245 2116
rect 1310 2106 1313 2173
rect 1322 2123 1325 2136
rect 1330 2123 1341 2126
rect 1330 2116 1333 2123
rect 1322 2113 1333 2116
rect 1310 2103 1317 2106
rect 1242 1906 1245 1986
rect 1250 1923 1253 2026
rect 1314 2013 1317 2103
rect 1258 1913 1261 2006
rect 1210 1903 1221 1906
rect 1242 1903 1257 1906
rect 1218 1856 1221 1903
rect 1210 1853 1221 1856
rect 1210 1746 1213 1853
rect 1254 1846 1257 1903
rect 1282 1873 1285 2006
rect 1330 1926 1333 2006
rect 1314 1923 1333 1926
rect 1346 1903 1349 2206
rect 1370 2203 1373 2243
rect 1354 2113 1357 2126
rect 1386 2083 1389 2136
rect 1394 2023 1397 2253
rect 1378 1963 1381 2016
rect 1402 1993 1405 2843
rect 1410 2813 1413 2826
rect 1410 2716 1413 2736
rect 1410 2713 1417 2716
rect 1414 2576 1417 2713
rect 1426 2623 1429 2816
rect 1442 2813 1445 2903
rect 1434 2783 1437 2806
rect 1442 2703 1445 2806
rect 1450 2803 1453 2826
rect 1458 2803 1461 2816
rect 1466 2776 1469 2963
rect 1450 2773 1469 2776
rect 1450 2696 1453 2773
rect 1474 2766 1477 2946
rect 1482 2876 1485 2926
rect 1510 2886 1513 2963
rect 1530 2933 1533 2973
rect 1522 2903 1525 2926
rect 1506 2883 1513 2886
rect 1482 2873 1493 2876
rect 1466 2763 1477 2766
rect 1442 2693 1453 2696
rect 1442 2676 1445 2693
rect 1438 2673 1445 2676
rect 1438 2616 1441 2673
rect 1438 2613 1445 2616
rect 1442 2596 1445 2613
rect 1450 2603 1453 2646
rect 1458 2633 1461 2716
rect 1410 2573 1417 2576
rect 1410 2553 1413 2573
rect 1426 2533 1429 2596
rect 1442 2593 1453 2596
rect 1434 2506 1437 2546
rect 1426 2503 1437 2506
rect 1426 2426 1429 2503
rect 1450 2426 1453 2593
rect 1466 2583 1469 2763
rect 1490 2746 1493 2873
rect 1506 2823 1509 2883
rect 1530 2836 1533 2926
rect 1562 2886 1565 2946
rect 1522 2833 1533 2836
rect 1546 2883 1565 2886
rect 1522 2786 1525 2833
rect 1546 2803 1549 2883
rect 1594 2876 1597 3040
rect 1618 2966 1621 3040
rect 1762 2976 1765 3040
rect 1618 2963 1633 2966
rect 1586 2873 1597 2876
rect 1586 2826 1589 2873
rect 1610 2856 1613 2926
rect 1630 2916 1633 2963
rect 1642 2923 1645 2976
rect 1762 2973 1769 2976
rect 1630 2913 1637 2916
rect 1610 2853 1617 2856
rect 1578 2823 1589 2826
rect 1522 2783 1549 2786
rect 1490 2743 1541 2746
rect 1490 2706 1493 2736
rect 1538 2733 1541 2743
rect 1522 2723 1541 2726
rect 1506 2713 1517 2716
rect 1474 2703 1493 2706
rect 1538 2626 1541 2723
rect 1546 2716 1549 2783
rect 1546 2713 1557 2716
rect 1554 2656 1557 2713
rect 1570 2693 1573 2716
rect 1546 2653 1557 2656
rect 1546 2633 1549 2653
rect 1578 2626 1581 2823
rect 1594 2783 1597 2816
rect 1614 2776 1617 2853
rect 1626 2813 1629 2826
rect 1634 2796 1637 2913
rect 1610 2773 1617 2776
rect 1630 2793 1637 2796
rect 1610 2733 1613 2773
rect 1630 2726 1633 2793
rect 1642 2733 1645 2806
rect 1658 2796 1661 2936
rect 1706 2923 1709 2956
rect 1754 2933 1757 2966
rect 1766 2926 1769 2973
rect 1778 2963 1781 3040
rect 1762 2923 1769 2926
rect 1722 2886 1725 2916
rect 1714 2883 1725 2886
rect 1674 2813 1677 2826
rect 1654 2793 1661 2796
rect 1674 2793 1677 2806
rect 1654 2746 1657 2793
rect 1654 2743 1661 2746
rect 1586 2723 1605 2726
rect 1630 2723 1637 2726
rect 1618 2633 1621 2716
rect 1634 2653 1637 2723
rect 1538 2623 1557 2626
rect 1578 2623 1589 2626
rect 1514 2593 1517 2616
rect 1498 2503 1501 2526
rect 1514 2483 1517 2586
rect 1546 2553 1549 2616
rect 1554 2613 1557 2623
rect 1554 2523 1557 2606
rect 1562 2523 1565 2536
rect 1426 2423 1437 2426
rect 1410 2316 1413 2336
rect 1418 2333 1421 2406
rect 1410 2313 1417 2316
rect 1414 2236 1417 2313
rect 1434 2256 1437 2423
rect 1442 2423 1453 2426
rect 1442 2413 1445 2423
rect 1554 2416 1557 2466
rect 1450 2403 1453 2416
rect 1458 2383 1461 2406
rect 1466 2336 1469 2416
rect 1474 2403 1477 2416
rect 1482 2393 1485 2416
rect 1522 2413 1557 2416
rect 1506 2393 1509 2406
rect 1450 2303 1453 2326
rect 1434 2253 1441 2256
rect 1410 2233 1417 2236
rect 1410 2013 1413 2233
rect 1418 2173 1421 2216
rect 1438 2176 1441 2253
rect 1450 2203 1453 2216
rect 1434 2173 1441 2176
rect 1434 2133 1437 2173
rect 1450 2133 1453 2156
rect 1418 2096 1421 2116
rect 1418 2093 1429 2096
rect 1450 2093 1453 2126
rect 1426 2036 1429 2093
rect 1418 2033 1429 2036
rect 1354 1953 1413 1956
rect 1354 1933 1357 1953
rect 1254 1843 1261 1846
rect 1234 1813 1245 1816
rect 1258 1796 1261 1843
rect 1266 1813 1269 1856
rect 1274 1806 1277 1836
rect 1290 1806 1293 1816
rect 1274 1803 1293 1806
rect 1258 1793 1293 1796
rect 1210 1743 1229 1746
rect 1202 1623 1205 1716
rect 1210 1613 1213 1736
rect 1226 1606 1229 1743
rect 1258 1733 1261 1793
rect 1290 1773 1293 1793
rect 1338 1766 1341 1816
rect 1346 1803 1349 1886
rect 1322 1763 1341 1766
rect 1266 1733 1269 1746
rect 1314 1726 1317 1736
rect 1322 1733 1325 1763
rect 1354 1756 1357 1876
rect 1362 1846 1365 1936
rect 1410 1933 1413 1953
rect 1418 1923 1421 2033
rect 1442 2003 1445 2016
rect 1450 1986 1453 2006
rect 1442 1983 1453 1986
rect 1426 1933 1429 1946
rect 1362 1843 1373 1846
rect 1370 1766 1373 1843
rect 1402 1813 1405 1836
rect 1386 1803 1397 1806
rect 1370 1763 1397 1766
rect 1354 1753 1373 1756
rect 1258 1713 1269 1716
rect 1266 1706 1269 1713
rect 1290 1706 1293 1726
rect 1266 1703 1293 1706
rect 1314 1723 1365 1726
rect 1218 1603 1229 1606
rect 1162 1423 1181 1426
rect 1138 1333 1141 1346
rect 1146 1326 1149 1416
rect 1178 1413 1181 1423
rect 1218 1416 1221 1603
rect 1242 1596 1245 1666
rect 1238 1593 1245 1596
rect 1238 1546 1241 1593
rect 1250 1583 1261 1586
rect 1238 1543 1245 1546
rect 1234 1513 1237 1526
rect 1242 1523 1245 1543
rect 1250 1516 1253 1583
rect 1266 1533 1269 1596
rect 1274 1523 1277 1556
rect 1282 1533 1285 1546
rect 1290 1533 1293 1626
rect 1298 1603 1301 1626
rect 1290 1516 1293 1526
rect 1250 1513 1293 1516
rect 1298 1513 1301 1526
rect 1202 1413 1221 1416
rect 1242 1413 1245 1426
rect 1314 1416 1317 1723
rect 1362 1713 1365 1723
rect 1322 1603 1325 1616
rect 1354 1613 1357 1626
rect 1370 1596 1373 1753
rect 1378 1706 1381 1726
rect 1386 1723 1389 1736
rect 1378 1703 1385 1706
rect 1382 1636 1385 1703
rect 1378 1633 1385 1636
rect 1378 1603 1381 1633
rect 1370 1593 1381 1596
rect 1154 1396 1157 1406
rect 1162 1403 1173 1406
rect 1154 1393 1161 1396
rect 1138 1323 1149 1326
rect 1130 1183 1133 1206
rect 1138 1123 1141 1323
rect 1158 1306 1161 1393
rect 1170 1313 1173 1403
rect 1158 1303 1165 1306
rect 1162 1266 1165 1303
rect 1158 1263 1165 1266
rect 1146 1213 1149 1226
rect 1158 1156 1161 1263
rect 1170 1213 1173 1256
rect 1186 1213 1189 1336
rect 1202 1246 1205 1413
rect 1274 1403 1277 1416
rect 1298 1413 1317 1416
rect 1266 1333 1269 1396
rect 1306 1356 1309 1406
rect 1330 1393 1333 1416
rect 1306 1353 1325 1356
rect 1218 1306 1221 1326
rect 1218 1303 1229 1306
rect 1202 1243 1209 1246
rect 1194 1196 1197 1236
rect 1190 1193 1197 1196
rect 1158 1153 1165 1156
rect 1154 1126 1157 1136
rect 1146 1123 1157 1126
rect 1162 1123 1165 1153
rect 1170 1133 1173 1166
rect 1146 1106 1149 1123
rect 1138 1103 1149 1106
rect 1138 1026 1141 1103
rect 1138 1023 1149 1026
rect 1146 1006 1149 1023
rect 1138 1003 1149 1006
rect 1154 986 1157 1116
rect 1162 1023 1165 1046
rect 1150 983 1157 986
rect 1130 813 1133 826
rect 1122 763 1129 766
rect 1090 643 1101 646
rect 1082 623 1093 626
rect 1058 593 1069 596
rect 1066 496 1069 593
rect 1090 513 1093 526
rect 1018 323 1021 486
rect 1042 413 1045 496
rect 1058 493 1069 496
rect 1058 426 1061 493
rect 1098 483 1101 643
rect 1106 616 1109 763
rect 1114 733 1117 746
rect 1114 623 1117 726
rect 1106 613 1113 616
rect 1110 466 1113 613
rect 1126 566 1129 763
rect 1126 563 1133 566
rect 1050 423 1061 426
rect 1106 463 1113 466
rect 1050 406 1053 423
rect 1034 393 1037 406
rect 1042 403 1053 406
rect 1042 286 1045 403
rect 1066 323 1069 406
rect 1106 376 1109 463
rect 1122 386 1125 406
rect 1130 386 1133 563
rect 1138 413 1141 936
rect 1150 826 1153 983
rect 1150 823 1157 826
rect 1154 806 1157 823
rect 1162 813 1165 1016
rect 1178 1003 1181 1186
rect 1190 1116 1193 1193
rect 1206 1186 1209 1243
rect 1226 1236 1229 1303
rect 1298 1296 1301 1326
rect 1322 1306 1325 1353
rect 1218 1233 1229 1236
rect 1290 1293 1301 1296
rect 1314 1303 1325 1306
rect 1290 1236 1293 1293
rect 1290 1233 1301 1236
rect 1218 1203 1221 1233
rect 1206 1183 1213 1186
rect 1210 1136 1213 1183
rect 1226 1173 1229 1216
rect 1234 1213 1245 1216
rect 1234 1153 1237 1206
rect 1250 1193 1253 1216
rect 1266 1203 1269 1226
rect 1298 1213 1301 1233
rect 1202 1133 1213 1136
rect 1274 1133 1285 1136
rect 1190 1113 1197 1116
rect 1202 1113 1205 1133
rect 1274 1116 1277 1133
rect 1266 1113 1277 1116
rect 1194 1096 1197 1113
rect 1194 1093 1205 1096
rect 1202 996 1205 1093
rect 1194 993 1205 996
rect 1170 933 1173 946
rect 1178 873 1181 936
rect 1186 813 1189 826
rect 1194 816 1197 993
rect 1226 983 1237 986
rect 1202 923 1205 936
rect 1210 933 1221 936
rect 1226 933 1229 956
rect 1234 946 1237 983
rect 1242 963 1245 1096
rect 1266 1036 1269 1113
rect 1266 1033 1277 1036
rect 1234 943 1241 946
rect 1210 923 1221 926
rect 1202 823 1213 826
rect 1194 813 1205 816
rect 1218 813 1221 923
rect 1154 803 1181 806
rect 1154 626 1157 646
rect 1150 623 1157 626
rect 1150 556 1153 623
rect 1162 616 1165 726
rect 1178 713 1181 803
rect 1186 706 1189 726
rect 1178 703 1189 706
rect 1162 613 1173 616
rect 1162 583 1165 606
rect 1150 553 1157 556
rect 1146 523 1149 536
rect 1154 533 1157 553
rect 1146 393 1149 426
rect 1122 383 1149 386
rect 1106 373 1113 376
rect 1110 296 1113 373
rect 1110 293 1117 296
rect 1034 283 1045 286
rect 978 233 989 236
rect 954 223 981 226
rect 954 213 957 223
rect 986 216 989 233
rect 962 213 989 216
rect 882 103 885 136
rect 930 123 941 126
rect 962 123 965 213
rect 1018 176 1021 206
rect 1034 183 1037 283
rect 1058 176 1061 216
rect 1114 203 1117 293
rect 1122 253 1125 383
rect 1130 323 1133 336
rect 1170 323 1173 613
rect 1178 603 1181 703
rect 1202 626 1205 813
rect 1186 546 1189 626
rect 1194 623 1205 626
rect 1194 593 1197 623
rect 1178 543 1189 546
rect 1178 486 1181 543
rect 1202 513 1205 536
rect 1210 523 1221 526
rect 1218 486 1221 523
rect 1178 483 1221 486
rect 1178 333 1181 356
rect 1186 323 1189 483
rect 1226 466 1229 916
rect 1238 826 1241 943
rect 1234 823 1241 826
rect 1234 803 1237 823
rect 1250 733 1253 926
rect 1258 913 1261 1006
rect 1266 986 1269 1016
rect 1274 1003 1277 1033
rect 1290 1026 1293 1206
rect 1314 1203 1317 1303
rect 1338 1286 1341 1566
rect 1330 1283 1341 1286
rect 1330 1216 1333 1283
rect 1330 1213 1341 1216
rect 1338 1193 1341 1213
rect 1346 1186 1349 1396
rect 1370 1393 1373 1593
rect 1394 1563 1397 1763
rect 1410 1416 1413 1906
rect 1442 1856 1445 1983
rect 1442 1853 1453 1856
rect 1450 1833 1453 1853
rect 1458 1846 1461 2336
rect 1466 2333 1477 2336
rect 1474 2303 1477 2333
rect 1482 2303 1485 2316
rect 1482 2183 1485 2196
rect 1466 2133 1469 2176
rect 1474 2123 1477 2136
rect 1474 1993 1477 2016
rect 1466 1903 1469 1936
rect 1458 1843 1485 1846
rect 1418 1793 1421 1806
rect 1474 1766 1477 1816
rect 1482 1783 1485 1843
rect 1490 1776 1493 2386
rect 1498 2093 1501 2116
rect 1514 2036 1517 2366
rect 1522 2323 1525 2413
rect 1538 2393 1549 2396
rect 1554 2383 1557 2406
rect 1538 2303 1549 2306
rect 1554 2213 1557 2316
rect 1578 2226 1581 2566
rect 1586 2463 1589 2623
rect 1594 2593 1597 2606
rect 1602 2553 1605 2626
rect 1594 2493 1597 2526
rect 1602 2453 1605 2536
rect 1618 2446 1621 2616
rect 1642 2593 1645 2616
rect 1650 2586 1653 2726
rect 1658 2606 1661 2743
rect 1666 2733 1669 2786
rect 1674 2733 1677 2766
rect 1690 2753 1693 2816
rect 1698 2803 1709 2806
rect 1706 2733 1709 2803
rect 1714 2716 1717 2883
rect 1762 2876 1765 2923
rect 1786 2913 1789 2936
rect 1794 2906 1797 3040
rect 1802 2933 1805 2956
rect 1810 2923 1813 2966
rect 1818 2923 1821 2936
rect 1762 2873 1769 2876
rect 1754 2846 1757 2866
rect 1746 2843 1757 2846
rect 1746 2776 1749 2843
rect 1766 2816 1769 2873
rect 1766 2813 1781 2816
rect 1762 2793 1765 2806
rect 1746 2773 1757 2776
rect 1722 2753 1725 2766
rect 1754 2756 1757 2773
rect 1754 2753 1773 2756
rect 1666 2613 1669 2716
rect 1706 2713 1717 2716
rect 1722 2743 1765 2746
rect 1690 2636 1693 2656
rect 1686 2633 1693 2636
rect 1706 2636 1709 2713
rect 1706 2633 1717 2636
rect 1658 2603 1669 2606
rect 1602 2443 1621 2446
rect 1634 2583 1653 2586
rect 1634 2443 1637 2583
rect 1686 2546 1689 2633
rect 1698 2556 1701 2616
rect 1698 2553 1705 2556
rect 1642 2533 1653 2536
rect 1602 2406 1605 2443
rect 1642 2436 1645 2526
rect 1658 2503 1661 2516
rect 1666 2463 1669 2536
rect 1674 2526 1677 2546
rect 1686 2543 1693 2546
rect 1674 2523 1681 2526
rect 1678 2456 1681 2523
rect 1674 2453 1681 2456
rect 1618 2416 1621 2426
rect 1626 2423 1629 2436
rect 1634 2433 1645 2436
rect 1610 2413 1629 2416
rect 1602 2403 1613 2406
rect 1610 2356 1613 2403
rect 1594 2353 1613 2356
rect 1594 2253 1597 2353
rect 1610 2333 1613 2353
rect 1634 2346 1637 2433
rect 1650 2403 1653 2436
rect 1658 2393 1661 2406
rect 1674 2366 1677 2453
rect 1674 2363 1681 2366
rect 1634 2343 1645 2346
rect 1610 2236 1613 2316
rect 1642 2296 1645 2343
rect 1634 2293 1645 2296
rect 1634 2236 1637 2293
rect 1610 2233 1621 2236
rect 1578 2223 1605 2226
rect 1570 2213 1589 2216
rect 1538 2193 1541 2206
rect 1554 2196 1557 2206
rect 1554 2193 1565 2196
rect 1554 2116 1557 2186
rect 1538 2103 1541 2116
rect 1546 2113 1557 2116
rect 1506 2033 1517 2036
rect 1506 1966 1509 2033
rect 1522 2003 1525 2026
rect 1546 2023 1549 2113
rect 1530 1986 1533 2016
rect 1522 1983 1533 1986
rect 1506 1963 1517 1966
rect 1498 1923 1501 1936
rect 1506 1923 1509 1946
rect 1498 1803 1501 1826
rect 1514 1813 1517 1963
rect 1522 1923 1525 1983
rect 1538 1923 1541 1996
rect 1490 1773 1501 1776
rect 1474 1763 1493 1766
rect 1426 1716 1429 1736
rect 1422 1713 1429 1716
rect 1422 1516 1425 1713
rect 1422 1513 1429 1516
rect 1426 1436 1429 1513
rect 1434 1506 1437 1726
rect 1466 1723 1469 1756
rect 1474 1733 1477 1746
rect 1490 1743 1493 1763
rect 1498 1733 1501 1773
rect 1530 1736 1533 1816
rect 1522 1733 1533 1736
rect 1522 1686 1525 1733
rect 1522 1683 1533 1686
rect 1442 1583 1445 1616
rect 1450 1563 1453 1606
rect 1498 1583 1501 1606
rect 1442 1513 1445 1546
rect 1458 1533 1461 1556
rect 1458 1516 1461 1526
rect 1466 1523 1469 1546
rect 1458 1513 1485 1516
rect 1434 1503 1445 1506
rect 1442 1486 1445 1503
rect 1442 1483 1453 1486
rect 1450 1436 1453 1483
rect 1426 1433 1433 1436
rect 1394 1333 1397 1416
rect 1410 1413 1421 1416
rect 1402 1363 1405 1406
rect 1370 1223 1373 1326
rect 1402 1303 1405 1336
rect 1418 1296 1421 1413
rect 1410 1293 1421 1296
rect 1402 1216 1405 1226
rect 1370 1213 1405 1216
rect 1410 1216 1413 1293
rect 1430 1236 1433 1433
rect 1442 1433 1453 1436
rect 1442 1296 1445 1433
rect 1474 1413 1477 1426
rect 1466 1333 1477 1336
rect 1466 1313 1469 1326
rect 1442 1293 1453 1296
rect 1450 1246 1453 1293
rect 1442 1243 1453 1246
rect 1430 1233 1437 1236
rect 1410 1213 1429 1216
rect 1370 1203 1373 1213
rect 1346 1183 1357 1186
rect 1290 1023 1297 1026
rect 1306 1023 1309 1126
rect 1266 983 1273 986
rect 1270 906 1273 983
rect 1266 903 1273 906
rect 1266 813 1269 903
rect 1282 813 1285 1016
rect 1294 926 1297 1023
rect 1314 1003 1317 1136
rect 1330 1133 1333 1146
rect 1354 1126 1357 1183
rect 1378 1173 1381 1206
rect 1394 1156 1397 1206
rect 1402 1163 1405 1206
rect 1394 1153 1405 1156
rect 1402 1126 1405 1153
rect 1410 1133 1413 1206
rect 1426 1196 1429 1213
rect 1434 1206 1437 1233
rect 1442 1213 1445 1243
rect 1474 1226 1477 1333
rect 1490 1296 1493 1416
rect 1498 1403 1501 1566
rect 1506 1543 1509 1616
rect 1530 1603 1533 1683
rect 1546 1536 1549 1726
rect 1522 1516 1525 1536
rect 1514 1513 1525 1516
rect 1530 1533 1549 1536
rect 1514 1436 1517 1513
rect 1514 1433 1525 1436
rect 1506 1306 1509 1416
rect 1506 1303 1513 1306
rect 1490 1293 1501 1296
rect 1466 1223 1477 1226
rect 1434 1203 1453 1206
rect 1426 1193 1437 1196
rect 1322 1103 1325 1126
rect 1346 1123 1357 1126
rect 1290 923 1297 926
rect 1306 943 1325 946
rect 1290 903 1293 923
rect 1306 896 1309 943
rect 1298 893 1309 896
rect 1298 816 1301 893
rect 1290 813 1301 816
rect 1314 816 1317 936
rect 1322 923 1325 943
rect 1330 933 1333 1036
rect 1346 976 1349 1123
rect 1394 1053 1397 1126
rect 1402 1123 1409 1126
rect 1406 1056 1409 1123
rect 1418 1063 1421 1136
rect 1434 1133 1437 1193
rect 1434 1103 1437 1116
rect 1406 1053 1413 1056
rect 1410 1036 1413 1053
rect 1410 1033 1421 1036
rect 1378 1013 1397 1016
rect 1346 973 1357 976
rect 1338 933 1341 966
rect 1354 926 1357 973
rect 1346 923 1357 926
rect 1322 913 1333 916
rect 1314 813 1321 816
rect 1290 753 1293 806
rect 1306 793 1309 806
rect 1318 766 1321 813
rect 1314 763 1321 766
rect 1314 746 1317 763
rect 1266 743 1317 746
rect 1266 603 1269 743
rect 1298 636 1301 736
rect 1298 633 1309 636
rect 1274 613 1301 616
rect 1306 613 1309 633
rect 1210 463 1229 466
rect 1210 356 1213 463
rect 1210 353 1229 356
rect 1122 186 1125 216
rect 1162 203 1165 276
rect 1194 233 1197 336
rect 1018 173 1061 176
rect 1114 183 1125 186
rect 994 93 997 136
rect 1058 133 1061 146
rect 1114 136 1117 183
rect 1074 113 1077 136
rect 1114 133 1125 136
rect 1138 133 1141 186
rect 1090 93 1093 116
rect 1122 113 1125 133
rect 1162 123 1165 146
rect 1218 113 1221 126
rect 1226 6 1229 353
rect 1234 323 1237 526
rect 1242 483 1245 536
rect 1250 533 1253 546
rect 1298 533 1301 613
rect 1314 533 1317 716
rect 1322 613 1325 626
rect 1242 423 1269 426
rect 1242 403 1245 423
rect 1250 403 1253 416
rect 1258 306 1261 416
rect 1266 413 1269 423
rect 1306 406 1309 526
rect 1322 513 1325 526
rect 1290 403 1309 406
rect 1330 403 1333 913
rect 1346 846 1349 923
rect 1342 843 1349 846
rect 1342 796 1345 843
rect 1354 813 1357 836
rect 1342 793 1349 796
rect 1346 773 1349 793
rect 1370 766 1373 1006
rect 1386 993 1389 1006
rect 1394 976 1397 1013
rect 1386 973 1397 976
rect 1386 916 1389 973
rect 1402 923 1405 1026
rect 1418 966 1421 1033
rect 1410 963 1421 966
rect 1410 916 1413 963
rect 1418 923 1421 936
rect 1426 933 1429 946
rect 1386 913 1405 916
rect 1410 913 1429 916
rect 1386 803 1389 856
rect 1402 816 1405 913
rect 1426 826 1429 913
rect 1434 903 1437 1056
rect 1450 1046 1453 1203
rect 1446 1043 1453 1046
rect 1446 956 1449 1043
rect 1466 1036 1469 1223
rect 1482 1196 1485 1216
rect 1498 1213 1501 1293
rect 1510 1226 1513 1303
rect 1522 1293 1525 1433
rect 1530 1423 1533 1533
rect 1546 1333 1549 1456
rect 1554 1403 1557 2106
rect 1562 2033 1565 2193
rect 1570 2123 1573 2213
rect 1594 2206 1597 2216
rect 1578 2203 1597 2206
rect 1602 2153 1605 2223
rect 1618 2146 1621 2233
rect 1630 2233 1637 2236
rect 1630 2186 1633 2233
rect 1658 2226 1661 2326
rect 1678 2276 1681 2363
rect 1690 2296 1693 2543
rect 1702 2506 1705 2553
rect 1714 2533 1717 2633
rect 1722 2623 1725 2743
rect 1730 2606 1733 2636
rect 1738 2613 1741 2736
rect 1746 2703 1749 2726
rect 1762 2723 1765 2743
rect 1762 2666 1765 2686
rect 1754 2663 1765 2666
rect 1754 2616 1757 2663
rect 1754 2613 1765 2616
rect 1726 2603 1733 2606
rect 1726 2526 1729 2603
rect 1738 2536 1741 2596
rect 1762 2593 1765 2613
rect 1770 2576 1773 2753
rect 1766 2573 1773 2576
rect 1738 2533 1749 2536
rect 1726 2523 1733 2526
rect 1754 2523 1757 2546
rect 1698 2503 1705 2506
rect 1698 2463 1701 2503
rect 1706 2376 1709 2486
rect 1730 2426 1733 2523
rect 1766 2466 1769 2573
rect 1766 2463 1773 2466
rect 1730 2423 1741 2426
rect 1706 2373 1717 2376
rect 1714 2313 1717 2373
rect 1738 2346 1741 2423
rect 1754 2403 1757 2416
rect 1770 2363 1773 2463
rect 1778 2376 1781 2813
rect 1786 2703 1789 2906
rect 1794 2903 1805 2906
rect 1802 2836 1805 2903
rect 1798 2833 1805 2836
rect 1798 2706 1801 2833
rect 1826 2816 1829 2976
rect 1850 2966 1853 3040
rect 1866 2976 1869 3040
rect 1866 2973 1889 2976
rect 1850 2963 1877 2966
rect 1834 2906 1837 2936
rect 1850 2906 1853 2936
rect 1834 2903 1853 2906
rect 1874 2903 1877 2963
rect 1850 2893 1853 2903
rect 1886 2886 1889 2973
rect 1898 2893 1901 2926
rect 1886 2883 1893 2886
rect 1810 2813 1837 2816
rect 1810 2723 1813 2813
rect 1818 2773 1821 2796
rect 1826 2723 1829 2806
rect 1850 2803 1853 2826
rect 1866 2756 1869 2846
rect 1890 2816 1893 2883
rect 1866 2753 1877 2756
rect 1858 2736 1861 2746
rect 1834 2706 1837 2736
rect 1798 2703 1805 2706
rect 1802 2626 1805 2703
rect 1826 2703 1837 2706
rect 1826 2646 1829 2703
rect 1826 2643 1837 2646
rect 1802 2623 1813 2626
rect 1786 2613 1805 2616
rect 1810 2606 1813 2623
rect 1794 2603 1813 2606
rect 1794 2536 1797 2603
rect 1826 2593 1829 2606
rect 1834 2573 1837 2643
rect 1842 2613 1845 2736
rect 1850 2723 1853 2736
rect 1858 2733 1869 2736
rect 1866 2706 1869 2733
rect 1874 2723 1877 2753
rect 1882 2733 1885 2816
rect 1890 2813 1901 2816
rect 1914 2813 1917 3040
rect 1930 2953 1933 3040
rect 1946 3013 1949 3040
rect 1890 2773 1893 2806
rect 1898 2796 1901 2813
rect 1898 2793 1909 2796
rect 1890 2733 1893 2746
rect 1906 2726 1909 2793
rect 1890 2723 1909 2726
rect 1866 2703 1873 2706
rect 1790 2533 1797 2536
rect 1790 2436 1793 2533
rect 1790 2433 1797 2436
rect 1786 2393 1789 2416
rect 1778 2373 1785 2376
rect 1738 2343 1749 2346
rect 1746 2296 1749 2343
rect 1690 2293 1701 2296
rect 1674 2273 1681 2276
rect 1642 2196 1645 2226
rect 1658 2223 1669 2226
rect 1666 2203 1669 2223
rect 1674 2213 1677 2273
rect 1698 2216 1701 2293
rect 1730 2293 1749 2296
rect 1730 2246 1733 2293
rect 1682 2196 1685 2216
rect 1642 2193 1685 2196
rect 1690 2213 1701 2216
rect 1722 2243 1733 2246
rect 1690 2193 1693 2213
rect 1722 2186 1725 2243
rect 1738 2186 1741 2236
rect 1630 2183 1637 2186
rect 1722 2183 1733 2186
rect 1738 2183 1745 2186
rect 1762 2183 1765 2326
rect 1782 2306 1785 2373
rect 1778 2303 1785 2306
rect 1778 2233 1781 2303
rect 1786 2213 1789 2286
rect 1794 2206 1797 2433
rect 1802 2403 1805 2526
rect 1810 2523 1813 2556
rect 1818 2476 1821 2536
rect 1842 2523 1845 2536
rect 1850 2523 1853 2616
rect 1858 2613 1861 2696
rect 1870 2626 1873 2703
rect 1890 2656 1893 2723
rect 1922 2686 1925 2926
rect 1930 2903 1933 2926
rect 1962 2826 1965 3040
rect 1986 2913 1989 2936
rect 1994 2866 1997 3040
rect 2002 2893 2005 2936
rect 2010 2923 2013 2966
rect 1930 2823 1965 2826
rect 1970 2863 1997 2866
rect 1930 2803 1933 2823
rect 1946 2726 1949 2816
rect 1970 2763 1973 2863
rect 2018 2856 2021 2936
rect 1978 2853 2021 2856
rect 1978 2813 1981 2853
rect 1954 2733 1957 2756
rect 1994 2733 1997 2836
rect 1938 2693 1941 2726
rect 1946 2723 1957 2726
rect 1922 2683 1933 2686
rect 1866 2623 1873 2626
rect 1882 2653 1893 2656
rect 1866 2533 1869 2623
rect 1874 2573 1877 2606
rect 1842 2513 1861 2516
rect 1818 2473 1853 2476
rect 1826 2396 1829 2446
rect 1834 2403 1845 2406
rect 1850 2403 1853 2473
rect 1818 2393 1829 2396
rect 1818 2336 1821 2393
rect 1858 2376 1861 2513
rect 1866 2503 1869 2526
rect 1834 2373 1861 2376
rect 1818 2333 1829 2336
rect 1802 2233 1805 2326
rect 1810 2266 1813 2316
rect 1826 2283 1829 2333
rect 1834 2316 1837 2373
rect 1842 2333 1861 2336
rect 1866 2323 1869 2426
rect 1874 2316 1877 2516
rect 1882 2413 1885 2653
rect 1930 2636 1933 2683
rect 1890 2546 1893 2626
rect 1898 2613 1901 2636
rect 1930 2633 1957 2636
rect 1922 2583 1925 2606
rect 1938 2576 1941 2626
rect 1946 2603 1949 2626
rect 1954 2613 1957 2633
rect 1994 2623 1997 2696
rect 2026 2676 2029 3016
rect 2034 2833 2037 2946
rect 2050 2923 2053 2936
rect 2074 2843 2077 3040
rect 2098 2903 2101 2926
rect 2114 2923 2133 2926
rect 2114 2886 2117 2923
rect 2098 2883 2117 2886
rect 2058 2833 2077 2836
rect 2042 2743 2045 2816
rect 2058 2813 2061 2833
rect 2066 2786 2069 2826
rect 2074 2813 2077 2833
rect 2066 2783 2077 2786
rect 2018 2673 2029 2676
rect 1978 2613 1997 2616
rect 1922 2573 1941 2576
rect 1922 2546 1925 2573
rect 1890 2543 1925 2546
rect 1890 2513 1893 2543
rect 1882 2393 1893 2396
rect 1882 2336 1885 2393
rect 1882 2333 1893 2336
rect 1834 2313 1869 2316
rect 1874 2313 1881 2316
rect 1866 2296 1869 2313
rect 1858 2293 1869 2296
rect 1810 2263 1821 2266
rect 1786 2203 1797 2206
rect 1610 2143 1621 2146
rect 1578 2096 1581 2136
rect 1594 2113 1597 2126
rect 1578 2093 1589 2096
rect 1586 2026 1589 2093
rect 1578 2023 1589 2026
rect 1578 1976 1581 2023
rect 1570 1973 1581 1976
rect 1570 1926 1573 1973
rect 1586 1933 1589 1986
rect 1570 1923 1581 1926
rect 1570 1646 1573 1786
rect 1578 1706 1581 1923
rect 1610 1813 1613 2143
rect 1626 2113 1629 2126
rect 1634 2033 1637 2183
rect 1650 2133 1653 2166
rect 1698 2143 1701 2166
rect 1634 2003 1637 2016
rect 1658 2006 1661 2136
rect 1698 2126 1701 2136
rect 1674 2123 1701 2126
rect 1714 2086 1717 2166
rect 1730 2123 1733 2183
rect 1742 2116 1745 2183
rect 1738 2113 1745 2116
rect 1738 2093 1741 2113
rect 1698 2083 1717 2086
rect 1642 1933 1645 2006
rect 1650 2003 1661 2006
rect 1586 1743 1589 1806
rect 1602 1776 1605 1806
rect 1626 1793 1629 1816
rect 1650 1806 1653 2003
rect 1666 1983 1669 2006
rect 1674 1976 1677 2036
rect 1698 2016 1701 2083
rect 1754 2076 1757 2146
rect 1786 2136 1789 2203
rect 1802 2183 1805 2206
rect 1818 2176 1821 2263
rect 1858 2246 1861 2293
rect 1858 2243 1869 2246
rect 1866 2226 1869 2243
rect 1878 2236 1881 2313
rect 1878 2233 1885 2236
rect 1866 2223 1877 2226
rect 1858 2203 1877 2206
rect 1882 2186 1885 2233
rect 1762 2133 1789 2136
rect 1810 2173 1821 2176
rect 1878 2183 1885 2186
rect 1810 2133 1813 2173
rect 1762 2113 1765 2126
rect 1770 2116 1773 2133
rect 1858 2123 1861 2156
rect 1770 2113 1781 2116
rect 1714 2073 1757 2076
rect 1698 2013 1709 2016
rect 1714 2013 1717 2073
rect 1722 2013 1725 2046
rect 1738 2013 1741 2036
rect 1762 2013 1765 2096
rect 1778 2066 1781 2113
rect 1770 2063 1781 2066
rect 1770 2043 1773 2063
rect 1834 2023 1837 2036
rect 1858 2013 1861 2056
rect 1878 2046 1881 2183
rect 1890 2173 1893 2333
rect 1878 2043 1885 2046
rect 1890 2043 1893 2126
rect 1898 2096 1901 2416
rect 1906 2403 1909 2536
rect 1922 2503 1925 2543
rect 1930 2513 1933 2546
rect 1946 2533 1949 2576
rect 1970 2533 1973 2586
rect 1962 2506 1965 2526
rect 1954 2503 1965 2506
rect 1954 2436 1957 2503
rect 1954 2433 1965 2436
rect 1962 2416 1965 2433
rect 1922 2343 1925 2396
rect 1930 2376 1933 2416
rect 1954 2413 1965 2416
rect 1954 2376 1957 2413
rect 1970 2403 1973 2526
rect 1986 2523 1989 2613
rect 2018 2606 2021 2673
rect 2034 2613 2037 2676
rect 2042 2656 2045 2726
rect 2074 2723 2077 2783
rect 2082 2733 2085 2856
rect 2098 2826 2101 2883
rect 2138 2866 2141 2926
rect 2154 2923 2157 2936
rect 2090 2823 2101 2826
rect 2122 2863 2141 2866
rect 2090 2763 2093 2823
rect 2122 2813 2125 2863
rect 2130 2816 2133 2856
rect 2162 2836 2165 2956
rect 2170 2903 2173 2936
rect 2178 2923 2181 2966
rect 2186 2846 2189 2936
rect 2226 2933 2229 2946
rect 2258 2936 2261 3040
rect 2258 2933 2269 2936
rect 2322 2933 2325 2946
rect 2138 2823 2141 2836
rect 2130 2813 2141 2816
rect 2146 2813 2149 2836
rect 2158 2833 2165 2836
rect 2178 2843 2189 2846
rect 2158 2746 2161 2833
rect 2170 2796 2173 2826
rect 2178 2813 2181 2843
rect 2194 2803 2197 2846
rect 2234 2813 2237 2826
rect 2250 2803 2253 2926
rect 2170 2793 2181 2796
rect 2178 2746 2181 2793
rect 2258 2766 2261 2826
rect 2266 2803 2269 2933
rect 2402 2926 2405 3040
rect 2434 2933 2445 2936
rect 2450 2933 2453 2946
rect 2306 2853 2309 2926
rect 2250 2763 2261 2766
rect 2130 2733 2133 2746
rect 2082 2673 2085 2726
rect 2130 2696 2133 2716
rect 2146 2713 2149 2746
rect 2158 2743 2165 2746
rect 2154 2706 2157 2726
rect 2122 2693 2133 2696
rect 2146 2703 2157 2706
rect 2042 2653 2069 2656
rect 2066 2616 2069 2653
rect 2122 2646 2125 2693
rect 2122 2643 2133 2646
rect 2066 2613 2077 2616
rect 1994 2573 1997 2606
rect 2018 2603 2029 2606
rect 2074 2603 2077 2613
rect 2002 2536 2005 2546
rect 1994 2533 2005 2536
rect 1930 2373 1957 2376
rect 1906 2143 1909 2286
rect 1922 2216 1925 2326
rect 1914 2213 1925 2216
rect 1906 2113 1909 2136
rect 1898 2093 1905 2096
rect 1882 2026 1885 2043
rect 1902 2036 1905 2093
rect 1898 2033 1905 2036
rect 1882 2023 1889 2026
rect 1706 1996 1709 2013
rect 1658 1973 1677 1976
rect 1658 1933 1661 1973
rect 1698 1933 1701 1996
rect 1706 1993 1717 1996
rect 1746 1993 1749 2006
rect 1714 1946 1717 1993
rect 1706 1943 1717 1946
rect 1706 1923 1709 1943
rect 1754 1923 1757 2006
rect 1634 1783 1637 1806
rect 1646 1803 1653 1806
rect 1602 1773 1613 1776
rect 1586 1723 1589 1736
rect 1610 1726 1613 1773
rect 1646 1756 1649 1803
rect 1646 1753 1653 1756
rect 1602 1723 1613 1726
rect 1578 1703 1589 1706
rect 1602 1703 1605 1723
rect 1634 1706 1637 1726
rect 1626 1703 1637 1706
rect 1562 1643 1573 1646
rect 1562 1523 1565 1643
rect 1586 1636 1589 1703
rect 1578 1633 1589 1636
rect 1626 1636 1629 1703
rect 1626 1633 1637 1636
rect 1578 1576 1581 1633
rect 1602 1613 1613 1616
rect 1578 1573 1605 1576
rect 1602 1556 1605 1573
rect 1586 1553 1605 1556
rect 1586 1446 1589 1553
rect 1586 1443 1605 1446
rect 1578 1423 1589 1426
rect 1578 1266 1581 1336
rect 1586 1313 1589 1326
rect 1562 1263 1581 1266
rect 1506 1223 1513 1226
rect 1478 1193 1485 1196
rect 1478 1126 1481 1193
rect 1478 1123 1485 1126
rect 1482 1103 1485 1123
rect 1490 1106 1493 1206
rect 1498 1123 1501 1136
rect 1506 1123 1509 1223
rect 1522 1203 1525 1236
rect 1530 1213 1533 1226
rect 1490 1103 1501 1106
rect 1530 1103 1533 1116
rect 1458 1033 1469 1036
rect 1446 953 1453 956
rect 1450 933 1453 953
rect 1458 916 1461 1033
rect 1450 913 1461 916
rect 1426 823 1437 826
rect 1402 813 1413 816
rect 1354 763 1373 766
rect 1338 646 1341 666
rect 1338 643 1345 646
rect 1342 556 1345 643
rect 1338 553 1345 556
rect 1338 533 1341 553
rect 1250 303 1261 306
rect 1250 196 1253 303
rect 1266 296 1269 336
rect 1282 316 1285 336
rect 1290 323 1293 403
rect 1306 316 1309 326
rect 1282 313 1309 316
rect 1330 296 1333 336
rect 1354 333 1357 763
rect 1378 626 1381 756
rect 1402 646 1405 806
rect 1418 753 1421 806
rect 1434 756 1437 823
rect 1450 806 1453 913
rect 1466 813 1469 1016
rect 1482 1013 1485 1066
rect 1498 1036 1501 1103
rect 1490 1033 1501 1036
rect 1490 1013 1493 1033
rect 1474 893 1477 1006
rect 1490 946 1493 1006
rect 1482 943 1493 946
rect 1450 803 1461 806
rect 1482 803 1485 943
rect 1490 916 1493 936
rect 1490 913 1501 916
rect 1506 913 1509 936
rect 1498 816 1501 913
rect 1498 813 1509 816
rect 1522 813 1525 1016
rect 1530 993 1533 1016
rect 1546 976 1549 1156
rect 1562 1003 1565 1263
rect 1586 1213 1589 1236
rect 1586 1026 1589 1126
rect 1594 1116 1597 1396
rect 1602 1323 1605 1443
rect 1610 1413 1613 1606
rect 1618 1523 1621 1616
rect 1634 1613 1637 1633
rect 1626 1563 1629 1606
rect 1634 1533 1637 1546
rect 1642 1543 1645 1736
rect 1650 1626 1653 1753
rect 1658 1646 1661 1796
rect 1682 1723 1685 1816
rect 1690 1803 1693 1816
rect 1690 1723 1693 1736
rect 1706 1723 1709 1806
rect 1714 1753 1717 1816
rect 1722 1793 1725 1806
rect 1658 1643 1669 1646
rect 1650 1623 1657 1626
rect 1654 1566 1657 1623
rect 1650 1563 1657 1566
rect 1650 1453 1653 1563
rect 1666 1546 1669 1643
rect 1658 1543 1669 1546
rect 1610 1306 1613 1406
rect 1618 1323 1621 1336
rect 1650 1333 1653 1416
rect 1658 1333 1661 1543
rect 1682 1536 1685 1706
rect 1690 1673 1693 1716
rect 1730 1636 1733 1906
rect 1738 1803 1741 1846
rect 1762 1803 1765 1936
rect 1834 1933 1837 1946
rect 1794 1833 1797 1866
rect 1802 1823 1805 1926
rect 1826 1883 1829 1926
rect 1786 1743 1789 1796
rect 1810 1793 1813 1816
rect 1826 1813 1829 1826
rect 1834 1776 1837 1926
rect 1842 1886 1845 2006
rect 1874 1993 1877 2016
rect 1850 1923 1853 1966
rect 1886 1956 1889 2023
rect 1874 1933 1877 1956
rect 1882 1953 1889 1956
rect 1882 1916 1885 1953
rect 1898 1946 1901 2033
rect 1898 1943 1905 1946
rect 1874 1913 1885 1916
rect 1842 1883 1849 1886
rect 1846 1806 1849 1883
rect 1826 1773 1837 1776
rect 1842 1803 1849 1806
rect 1786 1716 1789 1736
rect 1770 1713 1781 1716
rect 1786 1713 1797 1716
rect 1746 1636 1749 1656
rect 1730 1633 1749 1636
rect 1706 1613 1709 1626
rect 1714 1603 1717 1616
rect 1682 1533 1693 1536
rect 1666 1506 1669 1526
rect 1666 1503 1677 1506
rect 1674 1446 1677 1503
rect 1670 1443 1677 1446
rect 1670 1376 1673 1443
rect 1690 1426 1693 1533
rect 1714 1513 1717 1526
rect 1722 1496 1725 1616
rect 1730 1603 1733 1633
rect 1738 1523 1741 1626
rect 1746 1543 1749 1633
rect 1770 1626 1773 1713
rect 1794 1646 1797 1713
rect 1826 1706 1829 1773
rect 1842 1743 1845 1803
rect 1850 1713 1853 1786
rect 1826 1703 1837 1706
rect 1858 1703 1861 1896
rect 1866 1766 1869 1806
rect 1874 1776 1877 1913
rect 1890 1893 1893 1936
rect 1902 1886 1905 1943
rect 1898 1883 1905 1886
rect 1898 1846 1901 1883
rect 1890 1843 1901 1846
rect 1890 1833 1893 1843
rect 1906 1836 1909 1866
rect 1898 1833 1909 1836
rect 1882 1783 1885 1826
rect 1890 1816 1893 1826
rect 1914 1823 1917 2213
rect 1930 2206 1933 2236
rect 1946 2213 1949 2226
rect 1922 2203 1933 2206
rect 1922 2133 1925 2203
rect 1962 2186 1965 2396
rect 1994 2336 1997 2533
rect 2002 2523 2021 2526
rect 2026 2506 2029 2603
rect 2018 2503 2029 2506
rect 2018 2416 2021 2503
rect 2018 2413 2029 2416
rect 2002 2393 2013 2396
rect 2026 2376 2029 2413
rect 2018 2373 2029 2376
rect 1994 2333 2005 2336
rect 1978 2283 1981 2326
rect 2002 2276 2005 2333
rect 2018 2286 2021 2373
rect 2018 2283 2029 2286
rect 1994 2273 2005 2276
rect 1994 2216 1997 2273
rect 2026 2263 2029 2283
rect 2034 2246 2037 2506
rect 2030 2243 2037 2246
rect 1978 2206 1981 2216
rect 1994 2213 2013 2216
rect 2018 2213 2021 2226
rect 1978 2203 2005 2206
rect 1962 2183 1973 2186
rect 1994 2183 1997 2203
rect 1946 2133 1949 2156
rect 1954 2086 1957 2176
rect 1930 2083 1957 2086
rect 1930 1993 1933 2083
rect 1970 2076 1973 2183
rect 2010 2143 2013 2213
rect 2030 2176 2033 2243
rect 2018 2173 2033 2176
rect 1986 2133 2005 2136
rect 2018 2126 2021 2173
rect 2042 2166 2045 2416
rect 2058 2403 2061 2536
rect 2082 2523 2085 2626
rect 2122 2616 2125 2626
rect 2098 2613 2125 2616
rect 2130 2613 2133 2643
rect 2090 2533 2093 2556
rect 2074 2503 2077 2516
rect 2090 2423 2093 2526
rect 2098 2513 2101 2613
rect 2106 2556 2109 2606
rect 2106 2553 2117 2556
rect 2114 2533 2117 2553
rect 2122 2506 2125 2526
rect 2106 2503 2125 2506
rect 2146 2506 2149 2703
rect 2162 2686 2165 2743
rect 2170 2743 2181 2746
rect 2170 2723 2173 2743
rect 2158 2683 2165 2686
rect 2158 2566 2161 2683
rect 2158 2563 2165 2566
rect 2154 2533 2157 2546
rect 2146 2503 2153 2506
rect 2106 2486 2109 2503
rect 2102 2483 2109 2486
rect 2122 2493 2141 2496
rect 2102 2426 2105 2483
rect 2102 2423 2109 2426
rect 2066 2403 2069 2416
rect 2106 2403 2109 2423
rect 2114 2413 2117 2456
rect 2122 2433 2125 2493
rect 2130 2366 2133 2426
rect 2138 2403 2141 2493
rect 2150 2396 2153 2503
rect 2146 2393 2153 2396
rect 2146 2373 2149 2393
rect 2126 2363 2133 2366
rect 2050 2243 2053 2336
rect 2066 2306 2069 2326
rect 2066 2303 2077 2306
rect 2058 2266 2061 2286
rect 2058 2263 2065 2266
rect 2038 2163 2045 2166
rect 1962 2073 1973 2076
rect 2002 2123 2021 2126
rect 1962 2036 1965 2073
rect 2002 2036 2005 2123
rect 2026 2106 2029 2146
rect 2018 2103 2029 2106
rect 2018 2046 2021 2103
rect 2038 2096 2041 2163
rect 2050 2106 2053 2216
rect 2062 2206 2065 2263
rect 2074 2223 2077 2303
rect 2082 2293 2085 2336
rect 2062 2203 2069 2206
rect 2066 2146 2069 2203
rect 2058 2143 2069 2146
rect 2058 2123 2061 2143
rect 2090 2133 2093 2266
rect 2098 2216 2101 2236
rect 2098 2213 2105 2216
rect 2114 2213 2117 2326
rect 2126 2286 2129 2363
rect 2162 2306 2165 2563
rect 2170 2486 2173 2716
rect 2178 2616 2181 2696
rect 2194 2616 2197 2736
rect 2210 2623 2213 2736
rect 2234 2723 2237 2746
rect 2250 2686 2253 2763
rect 2290 2713 2293 2806
rect 2298 2733 2301 2816
rect 2306 2803 2309 2816
rect 2314 2723 2317 2826
rect 2354 2816 2357 2826
rect 2346 2813 2357 2816
rect 2330 2733 2333 2746
rect 2298 2713 2333 2716
rect 2250 2683 2261 2686
rect 2258 2646 2261 2683
rect 2242 2643 2261 2646
rect 2178 2613 2189 2616
rect 2194 2613 2213 2616
rect 2242 2613 2245 2643
rect 2266 2626 2269 2636
rect 2250 2623 2269 2626
rect 2298 2613 2301 2713
rect 2346 2696 2349 2813
rect 2362 2803 2365 2926
rect 2386 2923 2405 2926
rect 2370 2813 2373 2826
rect 2386 2806 2389 2923
rect 2386 2803 2413 2806
rect 2338 2693 2349 2696
rect 2338 2636 2341 2693
rect 2178 2543 2181 2606
rect 2178 2503 2181 2526
rect 2170 2483 2177 2486
rect 2174 2416 2177 2483
rect 2170 2413 2177 2416
rect 2170 2393 2173 2413
rect 2170 2333 2173 2346
rect 2146 2303 2165 2306
rect 2126 2283 2133 2286
rect 2130 2226 2133 2283
rect 2130 2223 2137 2226
rect 2102 2126 2105 2213
rect 2114 2163 2117 2206
rect 2122 2183 2125 2216
rect 2122 2146 2125 2176
rect 2134 2156 2137 2223
rect 2146 2163 2149 2303
rect 2154 2206 2157 2296
rect 2186 2266 2189 2613
rect 2194 2543 2197 2556
rect 2210 2373 2213 2613
rect 2314 2606 2317 2636
rect 2338 2633 2349 2636
rect 2346 2613 2349 2633
rect 2362 2613 2365 2736
rect 2378 2723 2381 2796
rect 2386 2713 2389 2736
rect 2394 2703 2397 2726
rect 2410 2723 2413 2803
rect 2426 2766 2429 2836
rect 2434 2823 2437 2926
rect 2458 2913 2461 2966
rect 2474 2946 2477 3040
rect 2562 2966 2565 3040
rect 2546 2963 2589 2966
rect 2474 2943 2485 2946
rect 2450 2786 2453 2856
rect 2466 2823 2469 2936
rect 2482 2846 2485 2943
rect 2506 2933 2509 2956
rect 2530 2923 2533 2946
rect 2546 2886 2549 2963
rect 2586 2923 2589 2963
rect 2602 2933 2605 2956
rect 2618 2946 2621 3040
rect 2618 2943 2629 2946
rect 2546 2883 2557 2886
rect 2474 2843 2485 2846
rect 2474 2816 2477 2843
rect 2490 2823 2501 2826
rect 2458 2813 2477 2816
rect 2458 2793 2461 2813
rect 2426 2763 2433 2766
rect 2418 2723 2421 2756
rect 2430 2716 2433 2763
rect 2426 2713 2433 2716
rect 2426 2693 2429 2713
rect 2394 2653 2437 2656
rect 2226 2533 2229 2606
rect 2234 2466 2237 2526
rect 2226 2463 2237 2466
rect 2226 2426 2229 2463
rect 2266 2436 2269 2606
rect 2298 2546 2301 2606
rect 2314 2603 2325 2606
rect 2322 2556 2325 2603
rect 2354 2563 2357 2606
rect 2314 2553 2325 2556
rect 2298 2543 2309 2546
rect 2282 2523 2285 2536
rect 2266 2433 2277 2436
rect 2226 2423 2269 2426
rect 2218 2323 2221 2356
rect 2186 2263 2221 2266
rect 2162 2213 2189 2216
rect 2194 2213 2205 2216
rect 2154 2203 2181 2206
rect 2118 2143 2125 2146
rect 2130 2153 2137 2156
rect 2102 2123 2109 2126
rect 2050 2103 2061 2106
rect 2034 2093 2041 2096
rect 2018 2043 2029 2046
rect 1954 2033 1965 2036
rect 1938 1903 1941 2006
rect 1954 1946 1957 2033
rect 1970 1956 1973 2026
rect 1970 1953 1977 1956
rect 1954 1943 1965 1946
rect 1962 1923 1965 1943
rect 1890 1813 1917 1816
rect 1874 1773 1885 1776
rect 1866 1763 1877 1766
rect 1766 1623 1773 1626
rect 1786 1643 1797 1646
rect 1754 1603 1757 1616
rect 1766 1546 1769 1623
rect 1786 1616 1789 1643
rect 1778 1613 1789 1616
rect 1802 1613 1805 1626
rect 1778 1596 1781 1613
rect 1834 1606 1837 1703
rect 1874 1606 1877 1763
rect 1890 1746 1893 1813
rect 1914 1783 1917 1813
rect 1886 1743 1893 1746
rect 1886 1686 1889 1743
rect 1898 1723 1901 1736
rect 1914 1723 1917 1776
rect 1922 1733 1925 1856
rect 1898 1696 1901 1716
rect 1898 1693 1909 1696
rect 1886 1683 1893 1686
rect 1826 1603 1845 1606
rect 1866 1603 1877 1606
rect 1778 1593 1789 1596
rect 1826 1593 1829 1603
rect 1762 1543 1769 1546
rect 1762 1526 1765 1543
rect 1754 1523 1765 1526
rect 1730 1503 1733 1516
rect 1722 1493 1741 1496
rect 1682 1423 1693 1426
rect 1682 1393 1685 1423
rect 1722 1413 1725 1426
rect 1698 1393 1701 1406
rect 1670 1373 1677 1376
rect 1674 1326 1677 1373
rect 1706 1343 1733 1346
rect 1610 1303 1621 1306
rect 1602 1213 1605 1246
rect 1618 1236 1621 1303
rect 1610 1233 1621 1236
rect 1602 1123 1605 1206
rect 1610 1133 1613 1233
rect 1618 1203 1621 1216
rect 1642 1203 1645 1326
rect 1666 1323 1677 1326
rect 1618 1123 1629 1126
rect 1594 1113 1605 1116
rect 1578 1023 1589 1026
rect 1538 973 1549 976
rect 1538 916 1541 973
rect 1554 923 1557 976
rect 1538 913 1549 916
rect 1426 753 1437 756
rect 1426 733 1429 753
rect 1458 736 1461 803
rect 1490 783 1493 806
rect 1514 793 1517 806
rect 1546 796 1549 913
rect 1562 906 1565 926
rect 1538 793 1549 796
rect 1558 903 1565 906
rect 1558 796 1561 903
rect 1570 803 1573 936
rect 1578 913 1581 926
rect 1558 793 1565 796
rect 1450 733 1461 736
rect 1450 666 1453 733
rect 1474 676 1477 776
rect 1474 673 1485 676
rect 1450 663 1461 666
rect 1370 623 1381 626
rect 1398 643 1405 646
rect 1458 643 1461 663
rect 1370 556 1373 623
rect 1370 553 1381 556
rect 1378 533 1381 553
rect 1386 516 1389 616
rect 1398 586 1401 643
rect 1410 633 1453 636
rect 1410 596 1413 633
rect 1418 613 1421 626
rect 1450 613 1453 633
rect 1482 626 1485 673
rect 1466 613 1469 626
rect 1474 623 1485 626
rect 1410 593 1421 596
rect 1398 583 1405 586
rect 1378 513 1389 516
rect 1378 446 1381 513
rect 1378 443 1389 446
rect 1386 366 1389 443
rect 1402 396 1405 583
rect 1418 553 1421 593
rect 1474 573 1477 623
rect 1410 513 1413 536
rect 1426 413 1429 536
rect 1458 526 1461 546
rect 1450 523 1461 526
rect 1402 393 1413 396
rect 1378 363 1389 366
rect 1378 316 1381 363
rect 1386 323 1389 356
rect 1410 316 1413 393
rect 1450 356 1453 523
rect 1466 506 1469 526
rect 1462 503 1469 506
rect 1462 416 1465 503
rect 1462 413 1469 416
rect 1466 393 1469 413
rect 1474 376 1477 496
rect 1490 413 1493 606
rect 1482 393 1485 406
rect 1474 373 1485 376
rect 1450 353 1461 356
rect 1378 313 1389 316
rect 1402 313 1413 316
rect 1266 293 1277 296
rect 1274 226 1277 293
rect 1322 293 1333 296
rect 1322 236 1325 293
rect 1322 233 1333 236
rect 1266 223 1277 226
rect 1266 203 1269 223
rect 1250 193 1261 196
rect 1258 123 1261 193
rect 1274 123 1277 136
rect 1298 113 1301 216
rect 1322 133 1325 216
rect 1330 196 1333 233
rect 1338 213 1341 306
rect 1402 296 1405 313
rect 1434 303 1437 336
rect 1442 296 1445 336
rect 1402 293 1445 296
rect 1346 213 1349 226
rect 1330 193 1341 196
rect 1338 126 1341 193
rect 1370 133 1389 136
rect 1330 123 1341 126
rect 1386 126 1389 133
rect 1386 123 1397 126
rect 1330 63 1333 123
rect 1402 113 1405 136
rect 1418 133 1421 146
rect 1426 133 1429 236
rect 1442 213 1445 226
rect 1458 156 1461 353
rect 1482 246 1485 373
rect 1506 313 1509 536
rect 1514 486 1517 736
rect 1538 616 1541 793
rect 1554 743 1557 756
rect 1562 626 1565 793
rect 1586 766 1589 1023
rect 1594 996 1597 1016
rect 1602 1003 1605 1113
rect 1626 1043 1629 1123
rect 1634 1106 1637 1126
rect 1634 1103 1645 1106
rect 1642 1036 1645 1103
rect 1634 1033 1645 1036
rect 1610 996 1613 1006
rect 1594 993 1613 996
rect 1594 923 1597 956
rect 1618 876 1621 1016
rect 1634 976 1637 1033
rect 1630 973 1637 976
rect 1630 926 1633 973
rect 1642 946 1645 966
rect 1642 943 1649 946
rect 1630 923 1637 926
rect 1634 903 1637 923
rect 1646 896 1649 943
rect 1642 893 1649 896
rect 1618 873 1629 876
rect 1602 793 1605 806
rect 1610 776 1613 866
rect 1578 763 1589 766
rect 1602 773 1613 776
rect 1570 723 1573 736
rect 1578 733 1581 763
rect 1602 726 1605 773
rect 1618 733 1621 816
rect 1626 803 1629 873
rect 1642 836 1645 893
rect 1658 873 1661 1266
rect 1666 1213 1669 1323
rect 1690 1246 1693 1326
rect 1706 1323 1709 1343
rect 1714 1323 1717 1336
rect 1722 1323 1725 1336
rect 1730 1323 1733 1343
rect 1690 1243 1709 1246
rect 1690 1223 1693 1236
rect 1698 1196 1701 1226
rect 1690 1193 1701 1196
rect 1690 1146 1693 1193
rect 1690 1143 1701 1146
rect 1698 1123 1701 1143
rect 1706 1133 1709 1243
rect 1730 1196 1733 1246
rect 1738 1216 1741 1493
rect 1754 1436 1757 1523
rect 1770 1443 1773 1536
rect 1786 1526 1789 1593
rect 1786 1523 1797 1526
rect 1754 1433 1765 1436
rect 1738 1213 1757 1216
rect 1738 1203 1741 1213
rect 1762 1196 1765 1433
rect 1778 1416 1781 1506
rect 1778 1413 1789 1416
rect 1794 1396 1797 1523
rect 1810 1513 1813 1536
rect 1818 1533 1829 1536
rect 1834 1533 1837 1546
rect 1818 1493 1821 1526
rect 1866 1446 1869 1603
rect 1890 1586 1893 1683
rect 1882 1583 1893 1586
rect 1882 1506 1885 1583
rect 1906 1576 1909 1693
rect 1930 1656 1933 1846
rect 1946 1836 1949 1906
rect 1938 1833 1949 1836
rect 1938 1816 1941 1833
rect 1938 1813 1949 1816
rect 1946 1736 1949 1813
rect 1962 1803 1965 1916
rect 1974 1856 1977 1953
rect 1986 1923 1989 2036
rect 1998 2033 2005 2036
rect 1998 1946 2001 2033
rect 1998 1943 2005 1946
rect 1994 1913 1997 1926
rect 1970 1853 1977 1856
rect 1938 1733 1949 1736
rect 1938 1713 1941 1733
rect 1962 1686 1965 1706
rect 1898 1573 1909 1576
rect 1922 1653 1933 1656
rect 1954 1683 1965 1686
rect 1898 1513 1901 1573
rect 1922 1526 1925 1653
rect 1954 1546 1957 1683
rect 1954 1543 1965 1546
rect 1882 1503 1893 1506
rect 1802 1423 1805 1446
rect 1866 1443 1877 1446
rect 1810 1403 1813 1426
rect 1850 1423 1869 1426
rect 1850 1413 1853 1423
rect 1794 1393 1805 1396
rect 1858 1393 1861 1416
rect 1866 1413 1869 1423
rect 1770 1326 1773 1346
rect 1802 1326 1805 1393
rect 1874 1376 1877 1443
rect 1890 1416 1893 1503
rect 1890 1413 1901 1416
rect 1858 1373 1877 1376
rect 1770 1323 1781 1326
rect 1802 1323 1813 1326
rect 1778 1236 1781 1323
rect 1810 1313 1813 1323
rect 1858 1256 1861 1373
rect 1882 1356 1885 1406
rect 1874 1353 1885 1356
rect 1874 1276 1877 1353
rect 1898 1346 1901 1413
rect 1890 1343 1901 1346
rect 1874 1273 1885 1276
rect 1858 1253 1877 1256
rect 1874 1236 1877 1253
rect 1730 1193 1741 1196
rect 1714 1106 1717 1136
rect 1722 1133 1733 1136
rect 1706 1103 1717 1106
rect 1706 1046 1709 1103
rect 1722 1063 1725 1126
rect 1674 1013 1677 1046
rect 1706 1043 1717 1046
rect 1674 916 1677 996
rect 1714 973 1717 1043
rect 1722 1013 1725 1026
rect 1738 1003 1741 1193
rect 1754 1193 1765 1196
rect 1774 1233 1781 1236
rect 1834 1233 1877 1236
rect 1754 1046 1757 1193
rect 1774 1186 1777 1233
rect 1834 1223 1837 1233
rect 1786 1203 1789 1216
rect 1750 1043 1757 1046
rect 1770 1183 1777 1186
rect 1750 986 1753 1043
rect 1770 1036 1773 1183
rect 1762 1033 1773 1036
rect 1750 983 1757 986
rect 1754 963 1757 983
rect 1682 943 1701 946
rect 1682 923 1685 943
rect 1690 916 1693 936
rect 1698 933 1701 943
rect 1674 913 1693 916
rect 1638 833 1645 836
rect 1638 786 1641 833
rect 1634 783 1641 786
rect 1602 723 1613 726
rect 1562 623 1573 626
rect 1538 613 1549 616
rect 1522 506 1525 526
rect 1538 523 1541 596
rect 1546 533 1549 613
rect 1562 603 1565 616
rect 1554 523 1557 566
rect 1570 546 1573 623
rect 1594 613 1597 636
rect 1610 603 1613 723
rect 1634 706 1637 783
rect 1650 733 1653 826
rect 1690 806 1693 913
rect 1698 883 1701 926
rect 1706 913 1709 926
rect 1714 806 1717 816
rect 1690 803 1709 806
rect 1714 803 1733 806
rect 1690 793 1709 796
rect 1690 756 1693 793
rect 1682 753 1693 756
rect 1626 703 1637 706
rect 1626 646 1629 703
rect 1642 696 1645 716
rect 1682 706 1685 753
rect 1730 746 1733 803
rect 1762 793 1765 1033
rect 1794 1026 1797 1216
rect 1802 1203 1805 1216
rect 1826 1186 1829 1216
rect 1818 1183 1829 1186
rect 1818 1036 1821 1183
rect 1834 1146 1837 1206
rect 1834 1143 1845 1146
rect 1834 1116 1837 1136
rect 1830 1113 1837 1116
rect 1830 1056 1833 1113
rect 1830 1053 1837 1056
rect 1818 1033 1829 1036
rect 1794 1023 1801 1026
rect 1770 926 1773 996
rect 1770 923 1781 926
rect 1786 816 1789 1016
rect 1798 966 1801 1023
rect 1794 963 1801 966
rect 1810 1013 1821 1016
rect 1794 943 1797 963
rect 1810 923 1813 1013
rect 1826 946 1829 1033
rect 1818 943 1829 946
rect 1818 826 1821 943
rect 1834 936 1837 1053
rect 1826 933 1837 936
rect 1818 823 1829 826
rect 1778 813 1789 816
rect 1730 743 1737 746
rect 1706 713 1709 736
rect 1682 703 1709 706
rect 1642 693 1653 696
rect 1650 646 1653 693
rect 1626 643 1633 646
rect 1618 613 1621 626
rect 1630 586 1633 643
rect 1642 643 1653 646
rect 1642 596 1645 643
rect 1650 603 1653 616
rect 1682 613 1685 636
rect 1642 593 1653 596
rect 1630 583 1637 586
rect 1562 543 1573 546
rect 1578 543 1581 576
rect 1522 503 1541 506
rect 1514 483 1525 486
rect 1522 426 1525 483
rect 1514 423 1525 426
rect 1474 243 1485 246
rect 1474 223 1477 243
rect 1450 153 1461 156
rect 1450 106 1453 153
rect 1474 113 1477 136
rect 1498 123 1501 146
rect 1506 133 1509 216
rect 1450 103 1461 106
rect 1458 16 1461 103
rect 1514 86 1517 423
rect 1538 346 1541 503
rect 1562 436 1565 543
rect 1570 516 1573 536
rect 1634 533 1637 583
rect 1570 513 1581 516
rect 1522 343 1541 346
rect 1554 433 1565 436
rect 1522 323 1525 343
rect 1538 303 1541 316
rect 1554 306 1557 433
rect 1578 426 1581 513
rect 1570 423 1581 426
rect 1570 353 1573 423
rect 1578 333 1581 396
rect 1650 393 1653 593
rect 1674 446 1677 576
rect 1698 556 1701 606
rect 1690 553 1701 556
rect 1690 523 1693 553
rect 1706 533 1709 703
rect 1734 696 1737 743
rect 1778 733 1781 813
rect 1794 806 1797 816
rect 1786 803 1797 806
rect 1730 693 1737 696
rect 1674 443 1685 446
rect 1682 396 1685 443
rect 1698 413 1701 526
rect 1714 426 1717 616
rect 1730 603 1733 693
rect 1738 436 1741 616
rect 1746 606 1749 726
rect 1786 723 1789 803
rect 1810 786 1813 816
rect 1802 783 1813 786
rect 1802 706 1805 783
rect 1826 776 1829 823
rect 1842 803 1845 1143
rect 1850 1123 1853 1216
rect 1858 1213 1861 1226
rect 1850 923 1853 1026
rect 1858 1013 1861 1206
rect 1866 1123 1869 1166
rect 1858 963 1861 1006
rect 1874 906 1877 1233
rect 1882 1216 1885 1273
rect 1890 1223 1893 1343
rect 1898 1306 1901 1326
rect 1898 1303 1905 1306
rect 1902 1236 1905 1303
rect 1898 1233 1905 1236
rect 1882 1213 1893 1216
rect 1898 1213 1901 1233
rect 1890 1016 1893 1213
rect 1914 1196 1917 1526
rect 1922 1523 1933 1526
rect 1930 1403 1933 1523
rect 1946 1506 1949 1526
rect 1942 1503 1949 1506
rect 1942 1436 1945 1503
rect 1942 1433 1949 1436
rect 1938 1366 1941 1416
rect 1946 1393 1949 1433
rect 1954 1413 1957 1516
rect 1962 1406 1965 1543
rect 1970 1476 1973 1853
rect 1978 1833 1997 1836
rect 1978 1823 1981 1833
rect 1986 1783 1989 1826
rect 1994 1823 1997 1833
rect 2002 1783 2005 1943
rect 2010 1833 2013 2026
rect 2026 2016 2029 2043
rect 2018 2013 2029 2016
rect 2026 1923 2029 1976
rect 2034 1913 2037 2093
rect 2042 2016 2045 2036
rect 2042 2013 2049 2016
rect 2046 1946 2049 2013
rect 2042 1943 2049 1946
rect 2042 1923 2045 1943
rect 2058 1906 2061 2103
rect 2082 1933 2085 2016
rect 2098 1933 2101 1946
rect 2106 1906 2109 2123
rect 2118 2046 2121 2143
rect 2130 2056 2133 2153
rect 2138 2133 2149 2136
rect 2130 2053 2137 2056
rect 2118 2043 2125 2046
rect 2122 2023 2125 2043
rect 2134 1996 2137 2053
rect 2146 2003 2149 2133
rect 2162 2113 2165 2136
rect 2178 2133 2181 2186
rect 2170 2093 2173 2126
rect 2186 2076 2189 2166
rect 2202 2156 2205 2213
rect 2210 2203 2213 2256
rect 2218 2163 2221 2263
rect 2226 2173 2229 2423
rect 2234 2163 2237 2346
rect 2242 2173 2245 2416
rect 2250 2196 2253 2326
rect 2258 2306 2261 2416
rect 2266 2393 2269 2423
rect 2274 2326 2277 2433
rect 2298 2403 2301 2536
rect 2306 2496 2309 2543
rect 2314 2516 2317 2553
rect 2378 2536 2381 2626
rect 2394 2613 2397 2653
rect 2410 2603 2413 2616
rect 2434 2613 2437 2653
rect 2442 2606 2445 2786
rect 2450 2783 2461 2786
rect 2450 2723 2453 2736
rect 2458 2733 2461 2783
rect 2482 2656 2485 2736
rect 2490 2703 2493 2716
rect 2478 2653 2485 2656
rect 2434 2603 2445 2606
rect 2322 2533 2341 2536
rect 2370 2533 2381 2536
rect 2322 2523 2325 2533
rect 2370 2523 2373 2533
rect 2314 2513 2341 2516
rect 2370 2513 2389 2516
rect 2394 2513 2397 2566
rect 2418 2523 2421 2556
rect 2434 2523 2437 2603
rect 2458 2526 2461 2616
rect 2478 2596 2481 2653
rect 2490 2606 2493 2646
rect 2498 2613 2501 2806
rect 2506 2676 2509 2846
rect 2514 2813 2517 2836
rect 2554 2806 2557 2883
rect 2570 2823 2573 2836
rect 2586 2833 2613 2836
rect 2578 2813 2581 2826
rect 2530 2803 2565 2806
rect 2514 2713 2517 2736
rect 2530 2696 2533 2796
rect 2546 2703 2549 2726
rect 2554 2723 2557 2736
rect 2562 2723 2565 2803
rect 2594 2743 2597 2826
rect 2610 2786 2613 2833
rect 2626 2793 2629 2943
rect 2650 2923 2653 2956
rect 2714 2933 2725 2936
rect 2762 2933 2765 2956
rect 2682 2903 2685 2926
rect 2714 2836 2717 2933
rect 2770 2896 2773 2926
rect 2778 2916 2781 2936
rect 2778 2913 2789 2916
rect 2762 2893 2773 2896
rect 2762 2846 2765 2893
rect 2786 2866 2789 2913
rect 2778 2863 2789 2866
rect 2762 2843 2773 2846
rect 2778 2843 2781 2863
rect 2610 2783 2621 2786
rect 2554 2696 2557 2716
rect 2530 2693 2541 2696
rect 2554 2693 2565 2696
rect 2506 2673 2517 2676
rect 2490 2603 2501 2606
rect 2478 2593 2485 2596
rect 2458 2523 2469 2526
rect 2306 2493 2317 2496
rect 2314 2426 2317 2493
rect 2306 2423 2317 2426
rect 2378 2426 2381 2513
rect 2378 2423 2397 2426
rect 2306 2403 2309 2423
rect 2314 2386 2317 2406
rect 2290 2383 2317 2386
rect 2290 2333 2293 2383
rect 2298 2333 2301 2376
rect 2314 2333 2333 2336
rect 2314 2326 2317 2333
rect 2274 2323 2285 2326
rect 2306 2323 2317 2326
rect 2258 2303 2269 2306
rect 2266 2246 2269 2303
rect 2258 2243 2269 2246
rect 2258 2213 2261 2243
rect 2282 2226 2285 2323
rect 2338 2313 2341 2416
rect 2394 2406 2397 2423
rect 2410 2413 2413 2506
rect 2386 2403 2397 2406
rect 2346 2343 2349 2386
rect 2386 2326 2389 2403
rect 2410 2376 2413 2396
rect 2406 2373 2413 2376
rect 2306 2233 2309 2246
rect 2266 2203 2269 2226
rect 2282 2223 2317 2226
rect 2314 2213 2317 2223
rect 2250 2193 2257 2196
rect 2290 2193 2293 2206
rect 2198 2153 2205 2156
rect 2198 2106 2201 2153
rect 2218 2133 2221 2156
rect 2242 2113 2245 2126
rect 2198 2103 2205 2106
rect 2178 2073 2189 2076
rect 2130 1993 2137 1996
rect 2146 1993 2157 1996
rect 2130 1973 2133 1993
rect 2178 1976 2181 2073
rect 2178 1973 2189 1976
rect 2114 1916 2117 1936
rect 2114 1913 2125 1916
rect 2050 1903 2061 1906
rect 2098 1903 2109 1906
rect 2050 1856 2053 1903
rect 2042 1853 2053 1856
rect 2026 1803 2029 1816
rect 1978 1713 1981 1726
rect 1986 1716 1989 1736
rect 1986 1713 1997 1716
rect 1994 1626 1997 1713
rect 1986 1623 1997 1626
rect 1986 1603 1989 1623
rect 2018 1613 2021 1716
rect 2034 1603 2037 1616
rect 2042 1613 2045 1853
rect 2058 1796 2061 1816
rect 2054 1793 2061 1796
rect 2054 1686 2057 1793
rect 2066 1696 2069 1886
rect 2074 1823 2077 1846
rect 2098 1816 2101 1903
rect 2122 1866 2125 1913
rect 2162 1873 2165 1936
rect 2114 1863 2125 1866
rect 2098 1813 2109 1816
rect 2114 1813 2117 1863
rect 2138 1813 2141 1846
rect 2082 1736 2085 1786
rect 2098 1773 2101 1796
rect 2106 1746 2109 1813
rect 2106 1743 2125 1746
rect 2082 1733 2117 1736
rect 2082 1713 2085 1733
rect 2066 1693 2077 1696
rect 2054 1683 2061 1686
rect 2058 1613 2061 1683
rect 2058 1596 2061 1606
rect 2034 1593 2061 1596
rect 1986 1523 1989 1536
rect 2034 1523 2037 1593
rect 2074 1586 2077 1693
rect 2090 1623 2093 1726
rect 2098 1723 2109 1726
rect 2098 1586 2101 1616
rect 2066 1583 2077 1586
rect 2090 1583 2101 1586
rect 2066 1523 2069 1583
rect 1970 1473 1981 1476
rect 1954 1403 1965 1406
rect 1938 1363 1949 1366
rect 1922 1203 1925 1256
rect 1930 1213 1933 1346
rect 1938 1316 1941 1336
rect 1946 1323 1949 1363
rect 1954 1333 1957 1403
rect 1978 1376 1981 1473
rect 2090 1446 2093 1583
rect 2106 1556 2109 1723
rect 2122 1703 2125 1743
rect 2138 1733 2141 1806
rect 2162 1646 2165 1726
rect 2170 1713 2173 1816
rect 2186 1813 2189 1973
rect 2194 1923 2197 1946
rect 2202 1916 2205 2103
rect 2254 2096 2257 2193
rect 2314 2166 2317 2186
rect 2250 2093 2257 2096
rect 2250 2076 2253 2093
rect 2242 2073 2253 2076
rect 2218 1966 2221 2016
rect 2242 1976 2245 2073
rect 2258 1993 2261 2016
rect 2242 1973 2253 1976
rect 2198 1913 2205 1916
rect 2210 1963 2221 1966
rect 2198 1836 2201 1913
rect 2210 1843 2213 1963
rect 2242 1923 2245 1956
rect 2250 1943 2253 1973
rect 2194 1833 2201 1836
rect 2178 1803 2189 1806
rect 2162 1643 2173 1646
rect 2114 1603 2117 1626
rect 2170 1623 2173 1643
rect 2122 1603 2125 1616
rect 2146 1576 2149 1606
rect 2178 1603 2181 1726
rect 2194 1616 2197 1833
rect 2218 1666 2221 1876
rect 2266 1813 2269 2166
rect 2310 2163 2317 2166
rect 2298 2123 2301 2146
rect 2310 2106 2313 2163
rect 2306 2103 2313 2106
rect 2306 2036 2309 2103
rect 2322 2053 2325 2206
rect 2306 2033 2317 2036
rect 2314 2016 2317 2033
rect 2282 2013 2309 2016
rect 2314 2013 2321 2016
rect 2274 1956 2277 2006
rect 2290 1993 2293 2006
rect 2298 1956 2301 2006
rect 2274 1953 2301 1956
rect 2306 1923 2309 2013
rect 2318 1926 2321 2013
rect 2314 1923 2321 1926
rect 2314 1906 2317 1923
rect 2306 1903 2317 1906
rect 2306 1856 2309 1903
rect 2306 1853 2317 1856
rect 2314 1836 2317 1853
rect 2314 1833 2325 1836
rect 2306 1823 2317 1826
rect 2306 1803 2309 1823
rect 2322 1816 2325 1833
rect 2314 1813 2325 1816
rect 2226 1783 2229 1796
rect 2306 1733 2309 1786
rect 2298 1706 2301 1726
rect 2314 1716 2317 1813
rect 2186 1613 2197 1616
rect 2210 1663 2221 1666
rect 2290 1703 2301 1706
rect 2310 1713 2317 1716
rect 2146 1573 2181 1576
rect 2106 1553 2117 1556
rect 2090 1443 2101 1446
rect 2042 1423 2089 1426
rect 2042 1413 2045 1423
rect 1970 1373 1981 1376
rect 1970 1343 1973 1373
rect 2034 1356 2037 1406
rect 2050 1403 2053 1416
rect 2058 1363 2061 1416
rect 1994 1353 2069 1356
rect 1962 1316 1965 1336
rect 1938 1313 1965 1316
rect 1954 1226 1957 1296
rect 1954 1223 1965 1226
rect 1938 1196 1941 1206
rect 1914 1193 1941 1196
rect 1914 1133 1917 1146
rect 1930 1133 1933 1176
rect 1946 1163 1949 1216
rect 1962 1176 1965 1223
rect 1994 1216 1997 1353
rect 2018 1306 2021 1346
rect 2066 1333 2069 1353
rect 2074 1323 2077 1406
rect 2086 1366 2089 1423
rect 2086 1363 2093 1366
rect 2018 1303 2037 1306
rect 1994 1213 2001 1216
rect 2018 1213 2021 1296
rect 2034 1286 2037 1303
rect 2034 1283 2045 1286
rect 2042 1226 2045 1283
rect 2034 1223 2045 1226
rect 1954 1173 1965 1176
rect 1954 1156 1957 1173
rect 1946 1153 1957 1156
rect 1938 1106 1941 1126
rect 1930 1103 1941 1106
rect 1890 1013 1901 1016
rect 1882 1003 1893 1006
rect 1898 946 1901 1013
rect 1906 1003 1909 1066
rect 1930 1016 1933 1103
rect 1930 1013 1941 1016
rect 1858 903 1877 906
rect 1882 943 1909 946
rect 1858 836 1861 903
rect 1882 896 1885 943
rect 1890 916 1893 936
rect 1906 923 1909 943
rect 1938 926 1941 1013
rect 1946 973 1949 1153
rect 1954 1116 1957 1136
rect 1954 1113 1965 1116
rect 1962 1046 1965 1113
rect 1954 1043 1965 1046
rect 1954 963 1957 1043
rect 1978 1013 1981 1146
rect 1986 1113 1989 1206
rect 1998 1166 2001 1213
rect 2010 1193 2013 1206
rect 2034 1196 2037 1223
rect 2082 1213 2085 1346
rect 2090 1323 2093 1363
rect 2098 1343 2101 1443
rect 2098 1313 2101 1336
rect 2106 1263 2109 1546
rect 2114 1376 2117 1553
rect 2122 1523 2125 1536
rect 2178 1526 2181 1573
rect 2186 1533 2189 1613
rect 2194 1576 2197 1606
rect 2210 1603 2213 1663
rect 2290 1646 2293 1703
rect 2290 1643 2301 1646
rect 2234 1576 2237 1616
rect 2290 1596 2293 1616
rect 2194 1573 2237 1576
rect 2274 1593 2293 1596
rect 2274 1536 2277 1593
rect 2218 1533 2277 1536
rect 2282 1533 2285 1586
rect 2290 1573 2293 1593
rect 2298 1526 2301 1643
rect 2310 1626 2313 1713
rect 2322 1633 2325 1726
rect 2310 1623 2317 1626
rect 2314 1543 2317 1623
rect 2162 1463 2165 1526
rect 2178 1523 2189 1526
rect 2282 1523 2301 1526
rect 2298 1513 2301 1523
rect 2330 1513 2333 2226
rect 2338 2193 2341 2206
rect 2338 2013 2341 2146
rect 2346 2106 2349 2326
rect 2362 2223 2365 2326
rect 2386 2323 2397 2326
rect 2354 2123 2357 2166
rect 2346 2103 2357 2106
rect 2354 2016 2357 2103
rect 2378 2053 2381 2306
rect 2394 2116 2397 2323
rect 2406 2156 2409 2373
rect 2418 2196 2421 2416
rect 2434 2403 2437 2506
rect 2442 2413 2445 2426
rect 2426 2323 2437 2326
rect 2434 2313 2437 2323
rect 2442 2313 2445 2326
rect 2426 2213 2429 2226
rect 2442 2213 2445 2306
rect 2450 2266 2453 2516
rect 2466 2456 2469 2523
rect 2462 2453 2469 2456
rect 2462 2336 2465 2453
rect 2474 2403 2477 2436
rect 2482 2413 2485 2593
rect 2498 2533 2501 2603
rect 2514 2596 2517 2673
rect 2538 2636 2541 2693
rect 2538 2633 2549 2636
rect 2538 2603 2541 2616
rect 2546 2613 2549 2633
rect 2562 2626 2565 2693
rect 2618 2636 2621 2783
rect 2634 2746 2637 2836
rect 2642 2823 2653 2826
rect 2658 2823 2661 2836
rect 2706 2833 2717 2836
rect 2650 2816 2653 2823
rect 2642 2753 2645 2816
rect 2650 2813 2669 2816
rect 2634 2743 2653 2746
rect 2618 2633 2629 2636
rect 2554 2623 2565 2626
rect 2506 2593 2517 2596
rect 2506 2563 2509 2593
rect 2514 2543 2517 2576
rect 2554 2556 2557 2623
rect 2594 2603 2597 2616
rect 2610 2596 2613 2616
rect 2626 2613 2629 2633
rect 2642 2626 2645 2736
rect 2650 2733 2653 2743
rect 2650 2716 2653 2726
rect 2658 2723 2661 2813
rect 2706 2803 2709 2833
rect 2714 2823 2749 2826
rect 2714 2813 2717 2823
rect 2730 2813 2741 2816
rect 2746 2813 2749 2823
rect 2722 2793 2725 2806
rect 2738 2753 2741 2806
rect 2674 2726 2677 2736
rect 2666 2723 2677 2726
rect 2666 2716 2669 2723
rect 2650 2713 2669 2716
rect 2674 2703 2677 2716
rect 2722 2656 2725 2736
rect 2770 2733 2773 2843
rect 2802 2836 2805 3006
rect 2798 2833 2805 2836
rect 2786 2803 2789 2816
rect 2798 2786 2801 2833
rect 2842 2826 2845 3040
rect 2842 2823 2853 2826
rect 2798 2783 2805 2786
rect 2818 2783 2821 2806
rect 2842 2793 2845 2816
rect 2850 2813 2853 2823
rect 2722 2653 2733 2656
rect 2642 2623 2653 2626
rect 2634 2613 2645 2616
rect 2606 2593 2613 2596
rect 2554 2553 2565 2556
rect 2538 2543 2557 2546
rect 2506 2396 2509 2536
rect 2522 2433 2525 2526
rect 2538 2433 2541 2526
rect 2554 2523 2557 2536
rect 2458 2333 2465 2336
rect 2498 2393 2509 2396
rect 2458 2286 2461 2333
rect 2498 2326 2501 2393
rect 2522 2326 2525 2426
rect 2546 2336 2549 2426
rect 2538 2333 2549 2336
rect 2498 2323 2509 2326
rect 2466 2303 2469 2316
rect 2506 2303 2509 2323
rect 2522 2323 2533 2326
rect 2458 2283 2469 2286
rect 2522 2283 2525 2323
rect 2450 2263 2457 2266
rect 2454 2206 2457 2263
rect 2426 2203 2437 2206
rect 2450 2203 2457 2206
rect 2418 2193 2445 2196
rect 2450 2183 2453 2203
rect 2466 2176 2469 2283
rect 2490 2203 2493 2216
rect 2514 2193 2517 2206
rect 2522 2193 2525 2266
rect 2530 2216 2533 2316
rect 2538 2263 2541 2333
rect 2554 2316 2557 2346
rect 2546 2313 2557 2316
rect 2562 2273 2565 2553
rect 2594 2516 2597 2536
rect 2586 2513 2597 2516
rect 2586 2456 2589 2513
rect 2586 2453 2597 2456
rect 2578 2333 2581 2436
rect 2594 2423 2597 2453
rect 2606 2446 2609 2593
rect 2606 2443 2613 2446
rect 2618 2443 2621 2606
rect 2626 2603 2637 2606
rect 2650 2556 2653 2623
rect 2666 2596 2669 2626
rect 2666 2593 2677 2596
rect 2634 2553 2653 2556
rect 2634 2446 2637 2553
rect 2674 2546 2677 2593
rect 2650 2523 2653 2546
rect 2666 2543 2677 2546
rect 2634 2443 2641 2446
rect 2610 2426 2613 2443
rect 2610 2423 2621 2426
rect 2602 2413 2613 2416
rect 2610 2403 2613 2413
rect 2618 2356 2621 2423
rect 2610 2353 2621 2356
rect 2570 2303 2573 2326
rect 2578 2256 2581 2326
rect 2610 2303 2613 2353
rect 2618 2333 2621 2346
rect 2626 2316 2629 2436
rect 2638 2376 2641 2443
rect 2634 2373 2641 2376
rect 2634 2326 2637 2373
rect 2642 2333 2645 2356
rect 2650 2326 2653 2426
rect 2658 2423 2661 2526
rect 2666 2373 2669 2543
rect 2682 2503 2685 2516
rect 2666 2333 2669 2346
rect 2634 2323 2645 2326
rect 2650 2323 2661 2326
rect 2626 2313 2637 2316
rect 2642 2296 2645 2323
rect 2546 2253 2581 2256
rect 2634 2293 2645 2296
rect 2546 2223 2549 2253
rect 2554 2243 2581 2246
rect 2530 2213 2549 2216
rect 2554 2213 2557 2243
rect 2406 2153 2413 2156
rect 2410 2133 2413 2153
rect 2394 2113 2413 2116
rect 2394 2026 2397 2113
rect 2418 2106 2421 2176
rect 2458 2173 2469 2176
rect 2458 2133 2461 2173
rect 2530 2146 2533 2206
rect 2526 2143 2533 2146
rect 2546 2186 2549 2213
rect 2562 2193 2565 2236
rect 2578 2226 2581 2243
rect 2578 2223 2597 2226
rect 2578 2186 2581 2216
rect 2602 2203 2605 2246
rect 2634 2216 2637 2293
rect 2634 2213 2645 2216
rect 2658 2213 2661 2323
rect 2642 2196 2645 2213
rect 2674 2203 2677 2436
rect 2682 2383 2685 2426
rect 2690 2413 2693 2436
rect 2698 2423 2701 2606
rect 2722 2573 2725 2626
rect 2714 2513 2717 2536
rect 2730 2533 2733 2653
rect 2746 2603 2749 2726
rect 2802 2646 2805 2783
rect 2858 2733 2861 2826
rect 2890 2813 2901 2816
rect 2922 2783 2925 2806
rect 2946 2766 2949 2816
rect 2898 2763 2949 2766
rect 2834 2713 2837 2726
rect 2802 2643 2809 2646
rect 2770 2633 2797 2636
rect 2762 2623 2789 2626
rect 2762 2593 2765 2616
rect 2786 2613 2789 2623
rect 2754 2513 2757 2526
rect 2794 2476 2797 2633
rect 2806 2546 2809 2643
rect 2842 2633 2845 2726
rect 2850 2706 2853 2726
rect 2850 2703 2861 2706
rect 2858 2646 2861 2703
rect 2850 2643 2861 2646
rect 2850 2626 2853 2643
rect 2802 2543 2809 2546
rect 2802 2503 2805 2543
rect 2818 2526 2821 2626
rect 2834 2623 2853 2626
rect 2834 2613 2837 2623
rect 2850 2613 2869 2616
rect 2842 2543 2845 2606
rect 2786 2473 2797 2476
rect 2706 2426 2709 2446
rect 2706 2423 2717 2426
rect 2690 2356 2693 2376
rect 2714 2366 2717 2423
rect 2738 2376 2741 2456
rect 2746 2403 2757 2406
rect 2762 2383 2765 2396
rect 2786 2386 2789 2473
rect 2786 2383 2797 2386
rect 2738 2373 2757 2376
rect 2686 2353 2693 2356
rect 2706 2363 2717 2366
rect 2686 2246 2689 2353
rect 2686 2243 2693 2246
rect 2690 2226 2693 2243
rect 2698 2233 2701 2326
rect 2690 2223 2701 2226
rect 2546 2183 2581 2186
rect 2410 2103 2421 2106
rect 2410 2046 2413 2103
rect 2434 2096 2437 2126
rect 2434 2093 2453 2096
rect 2350 2013 2357 2016
rect 2378 2023 2397 2026
rect 2402 2043 2413 2046
rect 2338 1723 2341 1976
rect 2350 1916 2353 2013
rect 2362 1933 2365 1996
rect 2350 1913 2357 1916
rect 2378 1913 2381 2023
rect 2354 1846 2357 1913
rect 2394 1893 2397 1926
rect 2402 1903 2405 2043
rect 2418 2013 2421 2026
rect 2426 2023 2445 2026
rect 2450 2023 2453 2093
rect 2482 2076 2485 2126
rect 2474 2073 2485 2076
rect 2474 2026 2477 2073
rect 2474 2023 2485 2026
rect 2426 2003 2429 2023
rect 2442 2016 2445 2023
rect 2346 1843 2357 1846
rect 2346 1636 2349 1843
rect 2354 1823 2381 1826
rect 2354 1813 2357 1823
rect 2362 1813 2373 1816
rect 2410 1813 2413 1946
rect 2426 1913 2429 1926
rect 2434 1823 2437 2016
rect 2442 2013 2453 2016
rect 2482 2003 2485 2023
rect 2498 2003 2501 2136
rect 2526 2076 2529 2143
rect 2538 2086 2541 2136
rect 2546 2123 2549 2183
rect 2538 2083 2549 2086
rect 2526 2073 2533 2076
rect 2530 2026 2533 2073
rect 2526 2023 2533 2026
rect 2514 1996 2517 2006
rect 2498 1993 2517 1996
rect 2442 1846 2445 1966
rect 2490 1933 2493 1966
rect 2498 1923 2501 1993
rect 2526 1976 2529 2023
rect 2522 1973 2529 1976
rect 2506 1923 2509 1936
rect 2442 1843 2453 1846
rect 2354 1766 2357 1806
rect 2362 1783 2365 1813
rect 2394 1776 2397 1806
rect 2410 1783 2413 1806
rect 2434 1776 2437 1816
rect 2394 1773 2437 1776
rect 2450 1766 2453 1843
rect 2354 1763 2373 1766
rect 2370 1666 2373 1763
rect 2442 1763 2453 1766
rect 2474 1813 2493 1816
rect 2394 1733 2397 1746
rect 2394 1723 2413 1726
rect 2354 1663 2373 1666
rect 2354 1643 2357 1663
rect 2346 1633 2365 1636
rect 2418 1633 2421 1736
rect 2442 1636 2445 1763
rect 2474 1716 2477 1813
rect 2466 1713 2477 1716
rect 2482 1713 2485 1726
rect 2466 1656 2469 1713
rect 2466 1653 2477 1656
rect 2442 1633 2453 1636
rect 2338 1613 2341 1626
rect 2338 1523 2357 1526
rect 2178 1413 2181 1436
rect 2186 1433 2245 1436
rect 2114 1373 2125 1376
rect 2122 1326 2125 1373
rect 2162 1363 2165 1406
rect 2186 1403 2189 1433
rect 2218 1413 2221 1426
rect 2234 1403 2237 1416
rect 2242 1413 2245 1433
rect 2242 1396 2245 1406
rect 2234 1393 2245 1396
rect 2114 1323 2125 1326
rect 2114 1303 2117 1323
rect 2114 1213 2117 1236
rect 2146 1213 2149 1336
rect 2194 1333 2197 1346
rect 2234 1336 2237 1393
rect 2226 1333 2237 1336
rect 2170 1236 2173 1256
rect 2170 1233 2177 1236
rect 2034 1193 2045 1196
rect 1994 1163 2001 1166
rect 1994 1096 1997 1163
rect 2042 1133 2045 1193
rect 2050 1133 2053 1206
rect 2098 1133 2101 1146
rect 2026 1113 2029 1126
rect 1994 1093 2053 1096
rect 2002 993 2005 1006
rect 2034 963 2037 1016
rect 1954 953 2013 956
rect 1954 933 1957 953
rect 1962 926 1965 936
rect 2010 933 2013 953
rect 2042 943 2045 1006
rect 1938 923 1965 926
rect 1890 913 1925 916
rect 1882 893 1893 896
rect 1858 833 1877 836
rect 1874 813 1877 833
rect 1890 816 1893 893
rect 1962 863 1965 923
rect 2026 903 2029 926
rect 2034 916 2037 926
rect 2050 916 2053 1093
rect 2082 1086 2085 1126
rect 2106 1123 2109 1206
rect 2114 1176 2117 1206
rect 2162 1186 2165 1206
rect 2138 1183 2165 1186
rect 2114 1173 2125 1176
rect 2122 1116 2125 1173
rect 2138 1133 2141 1183
rect 2174 1156 2177 1233
rect 2170 1153 2177 1156
rect 2114 1113 2125 1116
rect 2082 1083 2093 1086
rect 2114 1083 2117 1113
rect 2058 923 2061 996
rect 2034 913 2053 916
rect 1890 813 1901 816
rect 1866 803 1885 806
rect 1818 773 1829 776
rect 1818 713 1821 773
rect 1826 723 1829 736
rect 1802 703 1813 706
rect 1746 603 1757 606
rect 1762 546 1765 616
rect 1754 543 1765 546
rect 1754 523 1757 543
rect 1770 523 1773 536
rect 1738 433 1749 436
rect 1714 423 1741 426
rect 1678 393 1685 396
rect 1602 313 1605 326
rect 1554 303 1565 306
rect 1522 236 1525 256
rect 1562 236 1565 303
rect 1658 286 1661 356
rect 1666 333 1669 346
rect 1678 306 1681 393
rect 1714 376 1717 423
rect 1730 403 1733 416
rect 1738 413 1741 423
rect 1698 373 1717 376
rect 1698 323 1701 373
rect 1746 346 1749 433
rect 1742 343 1749 346
rect 1714 313 1717 336
rect 1678 303 1685 306
rect 1626 283 1661 286
rect 1522 233 1529 236
rect 1562 233 1581 236
rect 1526 176 1529 233
rect 1554 213 1557 226
rect 1562 206 1565 226
rect 1538 203 1565 206
rect 1562 193 1565 203
rect 1482 83 1517 86
rect 1522 173 1529 176
rect 1522 86 1525 173
rect 1554 123 1557 166
rect 1578 156 1581 233
rect 1626 166 1629 283
rect 1650 233 1661 236
rect 1682 226 1685 303
rect 1730 296 1733 316
rect 1722 293 1733 296
rect 1722 236 1725 293
rect 1722 233 1733 236
rect 1650 223 1661 226
rect 1674 223 1685 226
rect 1626 163 1637 166
rect 1574 153 1581 156
rect 1562 113 1565 146
rect 1562 86 1565 106
rect 1574 96 1577 153
rect 1602 143 1613 146
rect 1586 133 1605 136
rect 1610 116 1613 143
rect 1634 126 1637 163
rect 1650 133 1653 223
rect 1674 126 1677 223
rect 1730 213 1733 233
rect 1698 133 1701 206
rect 1742 146 1745 343
rect 1754 156 1757 336
rect 1770 323 1773 516
rect 1794 426 1797 626
rect 1810 603 1813 703
rect 1858 696 1861 716
rect 1850 693 1861 696
rect 1850 646 1853 693
rect 1850 643 1861 646
rect 1842 593 1845 606
rect 1850 456 1853 626
rect 1858 573 1861 643
rect 1874 613 1877 803
rect 1898 726 1901 813
rect 1898 723 1909 726
rect 1914 723 1917 736
rect 1874 563 1877 606
rect 1898 593 1901 616
rect 1906 543 1909 723
rect 1922 656 1925 736
rect 1946 733 1949 816
rect 1946 713 1949 726
rect 1962 713 1965 726
rect 1918 653 1925 656
rect 1918 596 1921 653
rect 1946 613 1957 616
rect 1914 593 1921 596
rect 1914 526 1917 593
rect 1970 583 1973 736
rect 2058 716 2061 736
rect 2074 723 2077 836
rect 2082 803 2085 1076
rect 2090 1003 2093 1083
rect 2146 1013 2149 1126
rect 2162 1123 2165 1136
rect 2170 1096 2173 1153
rect 2178 1113 2181 1126
rect 2170 1093 2181 1096
rect 2170 1066 2173 1086
rect 2162 1063 2173 1066
rect 2162 996 2165 1063
rect 2178 1003 2181 1093
rect 2186 1073 2189 1306
rect 2194 1196 2197 1206
rect 2202 1203 2205 1316
rect 2226 1246 2229 1333
rect 2234 1306 2237 1326
rect 2258 1313 2261 1326
rect 2266 1306 2269 1326
rect 2234 1303 2269 1306
rect 2282 1286 2285 1426
rect 2290 1406 2293 1436
rect 2290 1403 2301 1406
rect 2298 1356 2301 1403
rect 2290 1353 2301 1356
rect 2290 1333 2293 1353
rect 2330 1333 2333 1416
rect 2338 1403 2341 1496
rect 2370 1403 2373 1626
rect 2402 1606 2405 1626
rect 2394 1603 2405 1606
rect 2394 1536 2397 1603
rect 2394 1533 2405 1536
rect 2402 1513 2405 1533
rect 2410 1523 2413 1616
rect 2426 1526 2429 1626
rect 2434 1613 2437 1626
rect 2450 1586 2453 1633
rect 2474 1603 2477 1653
rect 2450 1583 2461 1586
rect 2418 1523 2429 1526
rect 2378 1326 2381 1416
rect 2394 1333 2397 1416
rect 2418 1343 2421 1523
rect 2426 1493 2429 1516
rect 2434 1373 2437 1536
rect 2458 1426 2461 1583
rect 2482 1523 2485 1706
rect 2490 1533 2493 1736
rect 2498 1723 2501 1856
rect 2522 1826 2525 1973
rect 2538 1923 2541 2016
rect 2546 1993 2549 2083
rect 2554 2036 2557 2056
rect 2554 2033 2561 2036
rect 2558 1956 2561 2033
rect 2554 1953 2561 1956
rect 2506 1813 2509 1826
rect 2522 1823 2533 1826
rect 2538 1823 2541 1896
rect 2546 1886 2549 1946
rect 2554 1933 2557 1953
rect 2570 1936 2573 2136
rect 2610 2086 2613 2106
rect 2602 2083 2613 2086
rect 2602 2036 2605 2083
rect 2618 2036 2621 2076
rect 2626 2043 2629 2116
rect 2634 2096 2637 2196
rect 2642 2193 2649 2196
rect 2646 2136 2649 2193
rect 2698 2186 2701 2223
rect 2642 2133 2649 2136
rect 2690 2183 2701 2186
rect 2642 2103 2645 2133
rect 2650 2096 2653 2116
rect 2634 2093 2653 2096
rect 2690 2096 2693 2183
rect 2706 2103 2709 2363
rect 2730 2333 2733 2346
rect 2738 2333 2749 2336
rect 2714 2313 2725 2316
rect 2738 2313 2741 2326
rect 2754 2323 2757 2373
rect 2794 2366 2797 2383
rect 2786 2363 2797 2366
rect 2762 2333 2765 2346
rect 2802 2323 2805 2446
rect 2810 2413 2813 2526
rect 2818 2523 2845 2526
rect 2858 2523 2861 2606
rect 2866 2533 2869 2606
rect 2818 2333 2821 2516
rect 2842 2446 2845 2523
rect 2866 2496 2869 2516
rect 2862 2493 2869 2496
rect 2842 2443 2853 2446
rect 2826 2423 2845 2426
rect 2850 2423 2853 2443
rect 2862 2426 2865 2493
rect 2862 2423 2869 2426
rect 2826 2413 2829 2423
rect 2842 2416 2845 2423
rect 2834 2333 2837 2416
rect 2842 2413 2853 2416
rect 2850 2403 2853 2413
rect 2714 2213 2717 2226
rect 2714 2133 2717 2146
rect 2730 2123 2733 2286
rect 2842 2266 2845 2396
rect 2858 2356 2861 2406
rect 2850 2353 2861 2356
rect 2866 2366 2869 2423
rect 2874 2413 2877 2526
rect 2882 2393 2885 2736
rect 2898 2733 2901 2763
rect 2890 2716 2893 2726
rect 2906 2723 2909 2736
rect 2922 2716 2925 2726
rect 2890 2713 2925 2716
rect 2930 2633 2933 2736
rect 2890 2593 2893 2606
rect 2898 2523 2901 2616
rect 2930 2576 2933 2606
rect 2954 2576 2957 2786
rect 2978 2733 2981 2776
rect 3002 2773 3005 2816
rect 3010 2756 3013 2806
rect 3002 2753 3013 2756
rect 3002 2666 3005 2753
rect 3002 2663 3009 2666
rect 2930 2573 2957 2576
rect 2890 2433 2893 2516
rect 2906 2383 2909 2406
rect 2866 2363 2901 2366
rect 2850 2333 2853 2353
rect 2858 2333 2861 2346
rect 2850 2316 2853 2326
rect 2866 2323 2869 2363
rect 2874 2336 2877 2356
rect 2874 2333 2893 2336
rect 2882 2316 2885 2326
rect 2850 2313 2885 2316
rect 2842 2263 2869 2266
rect 2746 2176 2749 2206
rect 2762 2183 2765 2206
rect 2786 2176 2789 2216
rect 2842 2213 2845 2236
rect 2746 2173 2789 2176
rect 2690 2093 2717 2096
rect 2602 2033 2613 2036
rect 2618 2033 2629 2036
rect 2578 1993 2581 2006
rect 2562 1906 2565 1936
rect 2570 1933 2589 1936
rect 2594 1926 2597 2016
rect 2610 1966 2613 2033
rect 2626 2003 2629 2033
rect 2602 1933 2605 1966
rect 2610 1963 2621 1966
rect 2578 1923 2597 1926
rect 2562 1903 2569 1906
rect 2546 1883 2557 1886
rect 2554 1826 2557 1883
rect 2546 1823 2557 1826
rect 2566 1826 2569 1903
rect 2566 1823 2573 1826
rect 2514 1783 2517 1806
rect 2530 1766 2533 1823
rect 2526 1763 2533 1766
rect 2506 1656 2509 1736
rect 2514 1723 2517 1736
rect 2526 1696 2529 1763
rect 2546 1756 2549 1823
rect 2562 1776 2565 1806
rect 2570 1803 2573 1823
rect 2578 1813 2581 1923
rect 2618 1916 2621 1963
rect 2650 1933 2653 2016
rect 2706 1993 2709 2016
rect 2666 1933 2669 1956
rect 2586 1853 2589 1916
rect 2610 1913 2621 1916
rect 2586 1793 2605 1796
rect 2586 1776 2589 1793
rect 2610 1786 2613 1913
rect 2618 1813 2621 1826
rect 2626 1813 2645 1816
rect 2626 1803 2629 1813
rect 2634 1786 2637 1806
rect 2610 1783 2637 1786
rect 2538 1753 2549 1756
rect 2538 1706 2541 1753
rect 2554 1733 2557 1776
rect 2562 1773 2581 1776
rect 2586 1773 2597 1776
rect 2578 1723 2581 1773
rect 2594 1716 2597 1773
rect 2586 1713 2597 1716
rect 2634 1716 2637 1726
rect 2642 1723 2645 1786
rect 2650 1716 2653 1746
rect 2634 1713 2653 1716
rect 2538 1703 2549 1706
rect 2526 1693 2533 1696
rect 2498 1653 2509 1656
rect 2498 1543 2501 1653
rect 2530 1626 2533 1693
rect 2514 1623 2533 1626
rect 2514 1606 2517 1623
rect 2522 1613 2541 1616
rect 2514 1603 2525 1606
rect 2546 1603 2549 1703
rect 2570 1623 2573 1636
rect 2522 1546 2525 1603
rect 2522 1543 2533 1546
rect 2498 1533 2509 1536
rect 2498 1506 2501 1526
rect 2490 1503 2501 1506
rect 2490 1436 2493 1503
rect 2490 1433 2501 1436
rect 2442 1423 2461 1426
rect 2442 1403 2445 1423
rect 2346 1323 2357 1326
rect 2362 1313 2365 1326
rect 2378 1323 2389 1326
rect 2258 1283 2285 1286
rect 2226 1243 2237 1246
rect 2210 1213 2213 1226
rect 2226 1213 2229 1236
rect 2234 1206 2237 1243
rect 2218 1196 2221 1206
rect 2194 1193 2221 1196
rect 2226 1203 2237 1206
rect 2194 1103 2197 1136
rect 2210 1006 2213 1193
rect 2226 1106 2229 1203
rect 2242 1193 2245 1206
rect 2258 1183 2261 1283
rect 2314 1203 2317 1236
rect 2322 1213 2325 1226
rect 2322 1183 2325 1206
rect 2258 1106 2261 1126
rect 2226 1103 2261 1106
rect 2274 1076 2277 1136
rect 2282 1133 2285 1176
rect 2338 1133 2341 1146
rect 2370 1133 2373 1206
rect 2378 1203 2381 1226
rect 2386 1206 2389 1323
rect 2434 1316 2437 1336
rect 2426 1313 2437 1316
rect 2426 1246 2429 1313
rect 2426 1243 2437 1246
rect 2394 1223 2429 1226
rect 2394 1213 2397 1223
rect 2386 1203 2413 1206
rect 2418 1136 2421 1216
rect 2426 1203 2429 1223
rect 2434 1213 2437 1243
rect 2442 1203 2445 1326
rect 2450 1213 2453 1326
rect 2458 1316 2461 1336
rect 2490 1333 2493 1416
rect 2498 1343 2501 1433
rect 2506 1316 2509 1516
rect 2530 1446 2533 1543
rect 2562 1523 2565 1546
rect 2578 1516 2581 1606
rect 2586 1533 2589 1713
rect 2658 1696 2661 1926
rect 2674 1783 2677 1826
rect 2682 1823 2685 1926
rect 2714 1923 2717 2093
rect 2738 2016 2741 2146
rect 2754 2023 2765 2026
rect 2690 1833 2709 1836
rect 2682 1806 2685 1816
rect 2698 1813 2701 1826
rect 2706 1813 2709 1833
rect 2682 1803 2709 1806
rect 2650 1693 2661 1696
rect 2594 1643 2621 1646
rect 2594 1523 2597 1643
rect 2610 1616 2613 1636
rect 2602 1613 2613 1616
rect 2618 1613 2621 1643
rect 2602 1533 2605 1613
rect 2626 1583 2629 1626
rect 2650 1606 2653 1693
rect 2666 1613 2669 1726
rect 2682 1723 2685 1803
rect 2714 1786 2717 1856
rect 2706 1783 2717 1786
rect 2706 1736 2709 1783
rect 2706 1733 2717 1736
rect 2714 1713 2717 1733
rect 2722 1703 2725 1936
rect 2730 1853 2733 2016
rect 2738 2013 2757 2016
rect 2754 1956 2757 2013
rect 2754 1953 2765 1956
rect 2738 1933 2749 1936
rect 2738 1913 2749 1916
rect 2762 1896 2765 1953
rect 2754 1893 2765 1896
rect 2754 1826 2757 1893
rect 2754 1823 2765 1826
rect 2762 1803 2765 1823
rect 2770 1803 2773 1836
rect 2778 1816 2781 2156
rect 2802 2003 2805 2126
rect 2810 2003 2813 2046
rect 2842 2003 2845 2106
rect 2850 2073 2853 2156
rect 2858 2093 2861 2146
rect 2866 2116 2869 2263
rect 2890 2213 2893 2333
rect 2898 2316 2901 2363
rect 2906 2323 2909 2336
rect 2898 2313 2909 2316
rect 2906 2236 2909 2313
rect 2930 2306 2933 2573
rect 2962 2533 2965 2616
rect 3006 2606 3009 2663
rect 3018 2613 3021 2626
rect 3006 2603 3013 2606
rect 2970 2513 2973 2526
rect 2970 2426 2973 2436
rect 2978 2433 2981 2446
rect 2986 2433 2989 2536
rect 2962 2403 2965 2426
rect 2970 2423 2989 2426
rect 2970 2353 2973 2416
rect 2954 2323 2957 2346
rect 2902 2233 2909 2236
rect 2922 2303 2933 2306
rect 2902 2186 2905 2233
rect 2902 2183 2909 2186
rect 2906 2126 2909 2183
rect 2922 2153 2925 2303
rect 2994 2216 2997 2306
rect 2946 2146 2949 2216
rect 2914 2143 2949 2146
rect 2994 2213 3005 2216
rect 2914 2133 2917 2143
rect 2922 2133 2949 2136
rect 2922 2126 2925 2133
rect 2898 2116 2901 2126
rect 2906 2123 2925 2126
rect 2938 2116 2941 2126
rect 2866 2113 2877 2116
rect 2874 2066 2877 2113
rect 2898 2113 2941 2116
rect 2898 2096 2901 2113
rect 2866 2063 2877 2066
rect 2890 2093 2901 2096
rect 2866 2046 2869 2063
rect 2862 2043 2869 2046
rect 2802 1986 2805 1996
rect 2802 1983 2813 1986
rect 2802 1923 2805 1936
rect 2778 1813 2789 1816
rect 2738 1723 2741 1786
rect 2778 1763 2781 1806
rect 2786 1773 2789 1813
rect 2810 1766 2813 1966
rect 2826 1803 2829 1836
rect 2842 1803 2845 1816
rect 2850 1803 2853 2016
rect 2862 1986 2865 2043
rect 2890 2036 2893 2093
rect 2906 2056 2909 2076
rect 2906 2053 2913 2056
rect 2890 2033 2901 2036
rect 2874 2013 2893 2016
rect 2862 1983 2869 1986
rect 2890 1983 2893 2006
rect 2898 2003 2901 2033
rect 2910 1996 2913 2053
rect 2930 2046 2933 2066
rect 2930 2043 2937 2046
rect 2906 1993 2913 1996
rect 2866 1946 2869 1983
rect 2866 1943 2885 1946
rect 2874 1923 2877 1936
rect 2882 1926 2885 1943
rect 2882 1923 2889 1926
rect 2874 1896 2877 1916
rect 2866 1893 2877 1896
rect 2866 1846 2869 1893
rect 2866 1843 2877 1846
rect 2786 1763 2813 1766
rect 2682 1623 2685 1636
rect 2650 1603 2685 1606
rect 2690 1603 2693 1616
rect 2730 1606 2733 1716
rect 2714 1603 2733 1606
rect 2658 1533 2661 1566
rect 2674 1533 2677 1546
rect 2682 1526 2685 1603
rect 2690 1533 2693 1586
rect 2738 1563 2741 1606
rect 2786 1603 2789 1763
rect 2810 1673 2813 1736
rect 2818 1703 2821 1726
rect 2826 1713 2829 1736
rect 2858 1733 2861 1816
rect 2866 1803 2869 1826
rect 2874 1803 2877 1843
rect 2886 1826 2889 1923
rect 2882 1823 2889 1826
rect 2882 1803 2885 1823
rect 2898 1763 2901 1906
rect 2874 1683 2877 1736
rect 2906 1686 2909 1993
rect 2922 1913 2925 2026
rect 2934 1926 2937 2043
rect 2930 1923 2937 1926
rect 2914 1833 2917 1906
rect 2930 1826 2933 1923
rect 2922 1823 2933 1826
rect 2906 1683 2913 1686
rect 2794 1613 2805 1616
rect 2610 1516 2613 1526
rect 2578 1513 2613 1516
rect 2666 1516 2669 1526
rect 2674 1523 2685 1526
rect 2698 1516 2701 1526
rect 2666 1513 2701 1516
rect 2730 1513 2733 1536
rect 2522 1443 2533 1446
rect 2458 1313 2469 1316
rect 2466 1236 2469 1313
rect 2458 1233 2469 1236
rect 2498 1313 2509 1316
rect 2514 1313 2517 1326
rect 2498 1236 2501 1313
rect 2522 1306 2525 1443
rect 2538 1403 2541 1426
rect 2514 1303 2525 1306
rect 2498 1233 2509 1236
rect 2458 1146 2461 1233
rect 2378 1133 2421 1136
rect 2434 1143 2461 1146
rect 2482 1143 2485 1216
rect 2506 1213 2509 1233
rect 2514 1186 2517 1303
rect 2530 1226 2533 1376
rect 2538 1336 2541 1346
rect 2538 1333 2549 1336
rect 2554 1333 2557 1426
rect 2570 1336 2573 1416
rect 2594 1413 2597 1426
rect 2634 1413 2653 1416
rect 2634 1336 2637 1413
rect 2570 1333 2589 1336
rect 2602 1333 2637 1336
rect 2658 1396 2661 1416
rect 2682 1403 2685 1416
rect 2690 1413 2693 1456
rect 2770 1436 2773 1536
rect 2794 1523 2797 1546
rect 2802 1533 2805 1606
rect 2810 1593 2813 1616
rect 2818 1603 2821 1626
rect 2858 1596 2861 1616
rect 2898 1613 2901 1676
rect 2850 1593 2861 1596
rect 2850 1546 2853 1593
rect 2874 1556 2877 1606
rect 2910 1586 2913 1683
rect 2906 1583 2913 1586
rect 2906 1566 2909 1583
rect 2866 1553 2877 1556
rect 2898 1563 2909 1566
rect 2850 1543 2861 1546
rect 2850 1513 2853 1526
rect 2858 1523 2861 1543
rect 2762 1433 2773 1436
rect 2762 1413 2765 1433
rect 2770 1423 2813 1426
rect 2770 1413 2773 1423
rect 2706 1396 2709 1406
rect 2658 1393 2709 1396
rect 2538 1313 2541 1326
rect 2546 1316 2549 1333
rect 2546 1313 2557 1316
rect 2554 1236 2557 1313
rect 2546 1233 2557 1236
rect 2530 1223 2537 1226
rect 2506 1183 2517 1186
rect 2346 1096 2349 1116
rect 2266 1073 2277 1076
rect 2218 1023 2245 1026
rect 2218 1013 2221 1023
rect 2202 1003 2213 1006
rect 2162 993 2173 996
rect 2170 956 2173 993
rect 2162 953 2173 956
rect 2114 913 2117 936
rect 2130 933 2133 946
rect 2138 926 2141 936
rect 2122 923 2141 926
rect 2122 903 2125 923
rect 2162 906 2165 953
rect 2226 933 2229 966
rect 2242 956 2245 1023
rect 2266 1013 2269 1073
rect 2234 953 2245 956
rect 2234 933 2237 953
rect 2162 903 2173 906
rect 2130 823 2133 836
rect 2114 716 2117 816
rect 2170 813 2173 903
rect 2202 806 2205 926
rect 2258 876 2261 936
rect 2266 926 2269 1006
rect 2322 986 2325 1026
rect 2338 1013 2341 1096
rect 2346 1093 2357 1096
rect 2354 1036 2357 1093
rect 2346 1033 2357 1036
rect 2346 1013 2349 1033
rect 2322 983 2333 986
rect 2290 953 2317 956
rect 2290 933 2293 953
rect 2306 926 2309 936
rect 2314 933 2317 953
rect 2330 926 2333 983
rect 2354 956 2357 1006
rect 2378 993 2381 1126
rect 2394 1113 2397 1126
rect 2418 1096 2421 1126
rect 2434 1123 2437 1143
rect 2506 1136 2509 1183
rect 2402 1093 2421 1096
rect 2402 966 2405 1093
rect 2426 976 2429 1116
rect 2442 1093 2445 1136
rect 2506 1133 2517 1136
rect 2482 1106 2485 1126
rect 2514 1113 2517 1133
rect 2466 1036 2469 1106
rect 2482 1103 2493 1106
rect 2522 1103 2525 1216
rect 2534 1136 2537 1223
rect 2530 1133 2537 1136
rect 2530 1103 2533 1133
rect 2546 1123 2549 1233
rect 2570 1173 2573 1216
rect 2586 1203 2589 1333
rect 2618 1186 2621 1326
rect 2658 1323 2661 1393
rect 2602 1183 2621 1186
rect 2602 1176 2605 1183
rect 2586 1173 2605 1176
rect 2490 1046 2493 1103
rect 2482 1043 2493 1046
rect 2466 1033 2473 1036
rect 2450 1016 2453 1026
rect 2434 1013 2453 1016
rect 2450 983 2453 1006
rect 2426 973 2433 976
rect 2402 963 2417 966
rect 2266 923 2301 926
rect 2306 923 2333 926
rect 2346 953 2357 956
rect 2258 873 2277 876
rect 2194 803 2205 806
rect 2274 803 2277 873
rect 2298 856 2301 923
rect 2346 906 2349 953
rect 2378 906 2381 926
rect 2402 913 2405 936
rect 2346 903 2381 906
rect 2414 896 2417 963
rect 2430 916 2433 973
rect 2442 933 2445 946
rect 2458 923 2461 1026
rect 2470 986 2473 1033
rect 2482 1003 2485 1043
rect 2506 993 2509 1026
rect 2522 1003 2525 1036
rect 2538 1023 2541 1116
rect 2586 1056 2589 1173
rect 2602 1133 2605 1156
rect 2618 1143 2621 1176
rect 2634 1133 2637 1216
rect 2666 1153 2669 1216
rect 2682 1096 2685 1326
rect 2698 1153 2709 1156
rect 2706 1136 2709 1153
rect 2578 1053 2589 1056
rect 2674 1093 2685 1096
rect 2698 1133 2709 1136
rect 2562 1013 2565 1036
rect 2470 983 2477 986
rect 2430 913 2437 916
rect 2410 893 2417 896
rect 2290 853 2301 856
rect 2290 813 2293 853
rect 2314 813 2333 816
rect 2386 813 2389 886
rect 2314 746 2317 813
rect 2410 806 2413 893
rect 2434 836 2437 913
rect 2458 886 2461 916
rect 2426 833 2437 836
rect 2450 883 2461 886
rect 2450 836 2453 883
rect 2474 836 2477 983
rect 2498 933 2501 966
rect 2522 923 2525 986
rect 2538 836 2541 1006
rect 2578 976 2581 1053
rect 2674 1036 2677 1093
rect 2698 1066 2701 1133
rect 2698 1063 2705 1066
rect 2714 1063 2717 1406
rect 2786 1403 2789 1416
rect 2810 1413 2813 1423
rect 2866 1413 2869 1553
rect 2874 1533 2877 1546
rect 2898 1446 2901 1563
rect 2898 1443 2909 1446
rect 2898 1413 2901 1426
rect 2738 1303 2741 1326
rect 2754 1323 2765 1326
rect 2794 1266 2797 1406
rect 2810 1333 2813 1346
rect 2818 1323 2821 1406
rect 2874 1403 2885 1406
rect 2906 1373 2909 1443
rect 2922 1403 2925 1823
rect 2946 1813 2949 2133
rect 2954 2116 2957 2136
rect 2994 2133 2997 2213
rect 3010 2116 3013 2603
rect 3018 2323 3021 2336
rect 2954 2113 2965 2116
rect 2962 2046 2965 2113
rect 3002 2113 3013 2116
rect 2954 2043 2965 2046
rect 2954 2013 2957 2043
rect 2978 2003 2981 2086
rect 2954 1933 2965 1936
rect 2954 1906 2957 1926
rect 2970 1923 2973 1946
rect 2954 1903 2965 1906
rect 2962 1836 2965 1903
rect 2954 1833 2965 1836
rect 2938 1746 2941 1806
rect 2954 1763 2957 1833
rect 3002 1826 3005 2113
rect 3002 1823 3013 1826
rect 2978 1803 2981 1816
rect 2938 1743 2949 1746
rect 2946 1723 2949 1743
rect 2986 1726 2989 1806
rect 2986 1723 3005 1726
rect 2954 1613 2957 1676
rect 3010 1663 3013 1823
rect 2946 1523 2949 1536
rect 3002 1523 3005 1546
rect 2946 1413 2949 1426
rect 3002 1383 3005 1416
rect 2898 1353 2933 1356
rect 2882 1323 2885 1336
rect 2778 1263 2797 1266
rect 2730 1213 2733 1226
rect 2762 1183 2765 1216
rect 2770 1213 2773 1226
rect 2778 1186 2781 1263
rect 2834 1213 2837 1236
rect 2842 1226 2845 1316
rect 2874 1303 2877 1316
rect 2898 1276 2901 1353
rect 2930 1333 2933 1353
rect 2914 1286 2917 1326
rect 2954 1286 2957 1326
rect 3010 1323 3013 1336
rect 2914 1283 2957 1286
rect 2898 1273 2909 1276
rect 2842 1223 2877 1226
rect 2786 1193 2789 1206
rect 2794 1203 2805 1206
rect 2850 1193 2853 1216
rect 2874 1213 2877 1223
rect 2858 1186 2861 1206
rect 2778 1183 2861 1186
rect 2866 1183 2869 1206
rect 2730 1123 2741 1126
rect 2746 1123 2749 1146
rect 2670 1033 2677 1036
rect 2578 973 2589 976
rect 2578 923 2581 946
rect 2586 883 2589 973
rect 2602 923 2605 996
rect 2618 933 2621 1016
rect 2634 963 2637 1006
rect 2670 986 2673 1033
rect 2682 1013 2685 1026
rect 2702 1006 2705 1063
rect 2714 1013 2717 1046
rect 2730 1013 2733 1026
rect 2702 1003 2709 1006
rect 2670 983 2677 986
rect 2674 963 2677 983
rect 2634 903 2637 916
rect 2602 853 2645 856
rect 2450 833 2461 836
rect 2426 813 2429 833
rect 2458 813 2461 833
rect 2466 833 2477 836
rect 2514 833 2557 836
rect 2466 813 2469 833
rect 2490 813 2493 826
rect 2322 803 2357 806
rect 2410 803 2421 806
rect 2314 743 2325 746
rect 2050 713 2061 716
rect 2050 666 2053 713
rect 2050 663 2061 666
rect 1906 523 1917 526
rect 1906 466 1909 523
rect 1922 496 1925 576
rect 1978 546 1981 566
rect 1970 543 1981 546
rect 1930 503 1933 536
rect 1938 523 1957 526
rect 1922 493 1941 496
rect 1906 463 1917 466
rect 1850 453 1893 456
rect 1794 423 1805 426
rect 1778 403 1781 416
rect 1770 223 1773 316
rect 1778 213 1781 336
rect 1786 323 1789 416
rect 1802 336 1805 423
rect 1826 406 1829 426
rect 1794 333 1805 336
rect 1818 403 1829 406
rect 1818 336 1821 403
rect 1834 376 1837 406
rect 1850 393 1853 406
rect 1874 376 1877 416
rect 1834 373 1877 376
rect 1818 333 1837 336
rect 1794 213 1797 333
rect 1754 153 1761 156
rect 1714 133 1717 146
rect 1742 143 1749 146
rect 1522 83 1533 86
rect 1458 13 1469 16
rect 1226 3 1245 6
rect 1242 0 1269 3
rect 1466 0 1469 13
rect 1482 0 1485 83
rect 1530 0 1533 83
rect 1554 83 1565 86
rect 1570 93 1577 96
rect 1594 113 1613 116
rect 1618 123 1637 126
rect 1650 123 1677 126
rect 1554 16 1557 83
rect 1570 63 1573 93
rect 1594 76 1597 113
rect 1578 73 1597 76
rect 1554 13 1565 16
rect 1562 0 1565 13
rect 1578 0 1581 73
rect 1594 0 1597 66
rect 1618 0 1621 123
rect 1650 0 1653 123
rect 1682 113 1685 126
rect 1690 113 1693 126
rect 1714 16 1717 126
rect 1738 113 1741 126
rect 1746 106 1749 143
rect 1738 103 1749 106
rect 1714 13 1725 16
rect 1722 0 1725 13
rect 1738 0 1741 103
rect 1758 76 1761 153
rect 1786 116 1789 206
rect 1802 123 1805 236
rect 1810 223 1813 316
rect 1818 213 1821 226
rect 1786 113 1797 116
rect 1794 76 1797 113
rect 1758 73 1765 76
rect 1762 16 1765 73
rect 1754 13 1765 16
rect 1786 73 1797 76
rect 1786 16 1789 73
rect 1786 13 1797 16
rect 1754 0 1757 13
rect 1794 0 1797 13
rect 1810 0 1813 206
rect 1818 76 1821 136
rect 1834 123 1837 333
rect 1850 323 1853 336
rect 1858 146 1861 326
rect 1866 303 1869 316
rect 1858 143 1885 146
rect 1858 113 1861 143
rect 1818 73 1837 76
rect 1834 16 1837 73
rect 1826 13 1837 16
rect 1826 0 1829 13
rect 1874 0 1877 136
rect 1882 116 1885 143
rect 1890 123 1893 453
rect 1914 413 1917 463
rect 1922 406 1925 476
rect 1938 436 1941 493
rect 1970 476 1973 543
rect 1986 486 1989 606
rect 2010 533 2013 616
rect 2058 613 2061 663
rect 2066 536 2069 616
rect 2018 533 2069 536
rect 2074 526 2077 716
rect 2114 713 2125 716
rect 2098 616 2101 706
rect 2122 636 2125 713
rect 2090 613 2101 616
rect 2114 633 2125 636
rect 2114 616 2117 633
rect 2146 626 2149 726
rect 2170 636 2173 736
rect 2210 713 2213 736
rect 2234 716 2237 736
rect 2298 726 2301 736
rect 2282 723 2301 726
rect 2170 633 2197 636
rect 2146 623 2157 626
rect 2114 613 2133 616
rect 2082 563 2085 606
rect 2090 596 2093 613
rect 2090 593 2101 596
rect 2098 556 2101 593
rect 2122 556 2125 606
rect 2098 553 2125 556
rect 2066 523 2077 526
rect 2018 513 2029 516
rect 2066 506 2069 523
rect 2018 503 2029 506
rect 1986 483 2005 486
rect 1970 473 1981 476
rect 1930 433 1941 436
rect 1930 413 1933 433
rect 1914 403 1925 406
rect 1914 313 1917 403
rect 1938 346 1941 416
rect 1962 346 1965 406
rect 1978 393 1981 473
rect 1930 343 1941 346
rect 1954 343 1965 346
rect 1922 246 1925 326
rect 1914 243 1925 246
rect 1930 243 1933 343
rect 1938 313 1941 326
rect 1954 266 1957 343
rect 1954 263 1965 266
rect 1914 213 1917 243
rect 1938 133 1941 206
rect 1962 193 1965 263
rect 1970 213 1973 336
rect 1978 323 1981 346
rect 2002 316 2005 483
rect 2026 413 2029 503
rect 2058 503 2069 506
rect 2074 503 2077 516
rect 2058 446 2061 503
rect 2058 443 2069 446
rect 2066 423 2069 443
rect 2082 416 2085 536
rect 2090 513 2093 526
rect 2082 413 2089 416
rect 2074 366 2077 406
rect 2086 366 2089 413
rect 2066 363 2077 366
rect 2082 363 2089 366
rect 2050 333 2053 346
rect 2066 323 2069 363
rect 1994 313 2005 316
rect 2074 313 2077 326
rect 1994 266 1997 313
rect 2066 286 2069 306
rect 1986 263 1997 266
rect 2058 283 2069 286
rect 1986 246 1989 263
rect 1982 243 1989 246
rect 1982 166 1985 243
rect 2018 206 2021 246
rect 2058 236 2061 283
rect 2082 263 2085 363
rect 2090 303 2093 346
rect 2058 233 2069 236
rect 2010 203 2021 206
rect 2010 186 2013 203
rect 2006 183 2013 186
rect 1982 163 1989 166
rect 1986 143 1989 163
rect 1882 113 1893 116
rect 1962 113 1965 126
rect 2006 116 2009 183
rect 2018 123 2021 196
rect 2050 133 2053 216
rect 2066 203 2069 233
rect 2074 123 2077 156
rect 2006 113 2013 116
rect 2010 3 2013 113
rect 2082 106 2085 236
rect 2074 103 2085 106
rect 2074 16 2077 103
rect 2074 13 2085 16
rect 1978 0 2013 3
rect 2082 0 2085 13
rect 2098 0 2101 553
rect 2106 503 2109 526
rect 2130 473 2133 613
rect 2138 513 2141 616
rect 2146 606 2149 616
rect 2154 613 2157 623
rect 2170 606 2173 633
rect 2202 623 2205 636
rect 2146 603 2173 606
rect 2178 603 2181 616
rect 2226 613 2229 716
rect 2234 713 2245 716
rect 2242 656 2245 713
rect 2234 653 2245 656
rect 2234 623 2237 653
rect 2250 606 2253 636
rect 2298 626 2301 716
rect 2322 646 2325 743
rect 2386 736 2389 796
rect 2378 716 2381 736
rect 2386 733 2397 736
rect 2418 733 2421 803
rect 2370 713 2381 716
rect 2370 666 2373 713
rect 2370 663 2381 666
rect 2314 643 2325 646
rect 2314 626 2317 643
rect 2290 623 2301 626
rect 2306 623 2317 626
rect 2306 606 2309 623
rect 2322 613 2325 626
rect 2378 613 2381 663
rect 2394 636 2397 733
rect 2390 633 2397 636
rect 2226 546 2229 606
rect 2250 603 2269 606
rect 2282 603 2309 606
rect 2226 543 2233 546
rect 2154 523 2197 526
rect 2106 313 2109 406
rect 2122 356 2125 426
rect 2154 393 2157 523
rect 2118 353 2125 356
rect 2118 296 2121 353
rect 2130 343 2141 346
rect 2178 333 2181 506
rect 2194 413 2197 516
rect 2202 393 2205 416
rect 2218 346 2221 536
rect 2230 496 2233 543
rect 2242 513 2277 516
rect 2282 496 2285 603
rect 2290 576 2293 596
rect 2290 573 2297 576
rect 2230 493 2237 496
rect 2234 366 2237 493
rect 2274 493 2285 496
rect 2202 343 2221 346
rect 2226 363 2237 366
rect 2202 316 2205 343
rect 2130 303 2133 316
rect 2194 313 2205 316
rect 2118 293 2125 296
rect 2114 183 2117 216
rect 2106 113 2109 136
rect 2122 123 2125 293
rect 2194 266 2197 313
rect 2210 296 2213 326
rect 2218 323 2221 336
rect 2226 316 2229 363
rect 2258 346 2261 436
rect 2242 343 2261 346
rect 2242 333 2245 343
rect 2226 313 2237 316
rect 2258 313 2261 336
rect 2210 293 2217 296
rect 2162 216 2165 266
rect 2194 263 2205 266
rect 2202 226 2205 263
rect 2194 223 2205 226
rect 2162 213 2173 216
rect 2138 123 2141 206
rect 2154 203 2165 206
rect 2154 123 2157 203
rect 2162 183 2165 196
rect 2170 126 2173 213
rect 2194 176 2197 223
rect 2194 173 2205 176
rect 2178 133 2181 156
rect 2170 123 2181 126
rect 2146 103 2149 116
rect 2178 113 2181 123
rect 2186 103 2189 126
rect 2202 113 2205 173
rect 2214 126 2217 293
rect 2234 236 2237 313
rect 2274 296 2277 493
rect 2294 486 2297 573
rect 2306 563 2349 566
rect 2306 533 2309 563
rect 2322 533 2325 556
rect 2346 523 2349 563
rect 2354 553 2357 606
rect 2390 586 2393 633
rect 2390 583 2397 586
rect 2394 563 2397 583
rect 2402 523 2405 626
rect 2434 613 2437 736
rect 2450 693 2453 736
rect 2466 733 2469 806
rect 2474 733 2493 736
rect 2514 716 2517 833
rect 2538 793 2541 816
rect 2554 803 2557 833
rect 2602 813 2605 853
rect 2634 813 2637 826
rect 2642 813 2645 853
rect 2690 813 2693 836
rect 2658 796 2661 806
rect 2698 803 2701 936
rect 2706 906 2709 1003
rect 2722 993 2725 1006
rect 2738 916 2741 946
rect 2746 933 2749 1066
rect 2754 1013 2757 1036
rect 2770 993 2773 1016
rect 2778 1006 2781 1183
rect 2810 1113 2813 1126
rect 2818 1123 2821 1166
rect 2906 1156 2909 1273
rect 2946 1163 2949 1226
rect 2978 1223 2981 1236
rect 2906 1153 2933 1156
rect 2882 1133 2885 1146
rect 2906 1136 2909 1153
rect 2898 1133 2909 1136
rect 2930 1133 2933 1153
rect 2786 1016 2789 1046
rect 2834 1026 2837 1116
rect 2874 1113 2877 1126
rect 2826 1023 2837 1026
rect 2786 1013 2797 1016
rect 2826 1013 2829 1023
rect 2778 1003 2789 1006
rect 2738 913 2745 916
rect 2706 903 2733 906
rect 2706 796 2709 816
rect 2722 813 2725 826
rect 2658 793 2709 796
rect 2714 793 2717 806
rect 2538 743 2565 746
rect 2658 743 2677 746
rect 2538 723 2541 743
rect 2514 713 2533 716
rect 2506 613 2509 686
rect 2530 656 2533 713
rect 2554 683 2557 736
rect 2562 723 2565 743
rect 2570 716 2573 736
rect 2562 713 2573 716
rect 2578 713 2581 736
rect 2530 653 2541 656
rect 2458 556 2461 606
rect 2538 576 2541 653
rect 2562 613 2565 713
rect 2650 696 2653 736
rect 2730 726 2733 903
rect 2742 766 2745 913
rect 2754 803 2757 926
rect 2770 813 2773 956
rect 2786 923 2789 1003
rect 2850 953 2853 1026
rect 2882 1023 2885 1036
rect 2898 1026 2901 1133
rect 2914 1086 2917 1126
rect 2954 1086 2957 1126
rect 3002 1123 3013 1126
rect 2914 1083 2957 1086
rect 2914 1053 2957 1056
rect 2898 1023 2909 1026
rect 2882 1003 2893 1006
rect 2850 916 2853 936
rect 2842 913 2853 916
rect 2842 856 2845 913
rect 2794 823 2797 856
rect 2842 853 2853 856
rect 2826 823 2829 836
rect 2850 803 2853 853
rect 2858 806 2861 966
rect 2866 913 2869 926
rect 2882 923 2885 1003
rect 2906 986 2909 1023
rect 2914 1013 2917 1053
rect 2954 1013 2957 1053
rect 3002 1013 3013 1016
rect 2930 986 2933 1006
rect 2906 983 2933 986
rect 2930 963 2933 983
rect 2866 813 2869 836
rect 2858 803 2869 806
rect 2738 763 2745 766
rect 2738 743 2741 763
rect 2818 733 2821 756
rect 2866 733 2869 803
rect 2882 753 2885 816
rect 2890 793 2893 936
rect 2938 923 2941 956
rect 3002 933 3005 1013
rect 2906 813 2909 856
rect 2954 823 2957 926
rect 2978 913 2981 926
rect 2994 823 2997 836
rect 2930 726 2933 806
rect 2722 723 2733 726
rect 2642 693 2653 696
rect 2570 613 2581 616
rect 2594 606 2597 616
rect 2642 613 2645 693
rect 2658 613 2669 616
rect 2570 593 2573 606
rect 2586 603 2597 606
rect 2586 596 2589 603
rect 2578 593 2589 596
rect 2530 573 2541 576
rect 2458 553 2469 556
rect 2434 523 2437 536
rect 2290 483 2297 486
rect 2290 303 2293 483
rect 2466 476 2469 553
rect 2482 523 2485 556
rect 2458 473 2469 476
rect 2298 423 2309 426
rect 2314 423 2317 436
rect 2298 403 2301 416
rect 2306 366 2309 423
rect 2394 373 2397 406
rect 2402 403 2405 416
rect 2410 396 2413 416
rect 2458 406 2461 473
rect 2402 393 2413 396
rect 2306 363 2317 366
rect 2314 333 2317 363
rect 2394 333 2397 356
rect 2402 343 2405 393
rect 2418 386 2421 406
rect 2458 403 2469 406
rect 2482 403 2485 516
rect 2466 386 2469 403
rect 2418 383 2429 386
rect 2274 293 2285 296
rect 2226 233 2237 236
rect 2226 176 2229 233
rect 2242 196 2245 206
rect 2250 203 2253 216
rect 2282 213 2285 293
rect 2322 213 2325 226
rect 2330 213 2333 326
rect 2354 226 2357 306
rect 2354 223 2365 226
rect 2338 213 2357 216
rect 2322 196 2325 206
rect 2346 203 2357 206
rect 2242 193 2261 196
rect 2322 193 2349 196
rect 2226 173 2237 176
rect 2210 123 2217 126
rect 2210 103 2213 123
rect 2234 96 2237 173
rect 2258 123 2261 193
rect 2322 133 2325 146
rect 2346 123 2349 193
rect 2362 166 2365 223
rect 2378 213 2381 326
rect 2410 236 2413 346
rect 2426 336 2429 383
rect 2458 383 2477 386
rect 2418 333 2429 336
rect 2418 313 2421 333
rect 2442 323 2445 376
rect 2458 316 2461 383
rect 2474 333 2477 383
rect 2498 323 2501 356
rect 2514 316 2517 526
rect 2530 523 2533 573
rect 2578 523 2581 593
rect 2594 556 2597 596
rect 2594 553 2605 556
rect 2602 486 2605 553
rect 2618 533 2621 556
rect 2634 536 2637 606
rect 2674 596 2677 636
rect 2682 623 2685 646
rect 2730 633 2733 723
rect 2658 593 2677 596
rect 2706 593 2741 596
rect 2642 543 2645 576
rect 2658 536 2661 593
rect 2634 533 2661 536
rect 2594 483 2605 486
rect 2530 413 2533 426
rect 2562 353 2565 416
rect 2578 403 2581 426
rect 2594 393 2597 483
rect 2442 313 2461 316
rect 2410 233 2429 236
rect 2362 163 2405 166
rect 2362 126 2365 163
rect 2354 123 2365 126
rect 2402 123 2405 163
rect 2442 133 2445 313
rect 2474 256 2477 316
rect 2506 313 2517 316
rect 2554 313 2557 326
rect 2570 256 2573 336
rect 2594 323 2597 376
rect 2610 296 2613 316
rect 2466 253 2477 256
rect 2538 253 2573 256
rect 2606 293 2613 296
rect 2466 206 2469 253
rect 2482 233 2485 246
rect 2490 213 2493 226
rect 2466 203 2477 206
rect 2474 123 2477 203
rect 2538 143 2541 253
rect 2554 243 2565 246
rect 2562 213 2565 243
rect 2606 176 2609 293
rect 2618 243 2621 526
rect 2634 516 2637 533
rect 2634 513 2645 516
rect 2698 513 2701 526
rect 2642 446 2645 513
rect 2634 443 2645 446
rect 2634 406 2637 443
rect 2682 423 2709 426
rect 2682 413 2685 423
rect 2706 413 2709 423
rect 2634 403 2645 406
rect 2642 346 2645 403
rect 2638 343 2645 346
rect 2638 286 2641 343
rect 2634 283 2641 286
rect 2606 173 2613 176
rect 2274 103 2277 116
rect 2226 93 2237 96
rect 2226 0 2229 93
rect 2354 0 2357 123
rect 2546 43 2549 146
rect 2554 113 2557 126
rect 2578 106 2581 126
rect 2610 113 2613 173
rect 2618 106 2621 216
rect 2634 213 2637 283
rect 2626 113 2629 126
rect 2634 116 2637 206
rect 2634 113 2645 116
rect 2578 103 2621 106
rect 2618 73 2621 103
rect 2650 43 2653 326
rect 2674 123 2677 406
rect 2698 346 2701 406
rect 2714 403 2717 566
rect 2730 513 2733 526
rect 2722 413 2725 426
rect 2690 343 2701 346
rect 2690 326 2693 343
rect 2698 333 2717 336
rect 2690 323 2701 326
rect 2698 316 2701 323
rect 2698 313 2717 316
rect 2698 163 2701 206
rect 2706 203 2709 216
rect 2722 193 2725 326
rect 2738 213 2741 593
rect 2754 563 2757 726
rect 2850 686 2853 726
rect 2890 686 2893 726
rect 2930 723 2949 726
rect 2986 723 2997 726
rect 2850 683 2893 686
rect 2786 613 2789 646
rect 2810 623 2813 636
rect 2834 626 2837 646
rect 2826 623 2837 626
rect 2778 563 2781 606
rect 2802 593 2805 616
rect 2826 576 2829 623
rect 2850 616 2853 626
rect 2842 613 2853 616
rect 2858 616 2861 636
rect 2866 623 2869 646
rect 2858 613 2877 616
rect 2930 613 2933 626
rect 2826 573 2837 576
rect 2754 423 2757 546
rect 2770 523 2773 536
rect 2818 513 2821 526
rect 2770 466 2773 486
rect 2770 463 2781 466
rect 2778 416 2781 463
rect 2770 413 2781 416
rect 2690 113 2693 136
rect 2706 133 2709 156
rect 2746 103 2749 126
rect 2754 0 2757 406
rect 2770 336 2773 413
rect 2802 396 2805 416
rect 2826 403 2829 426
rect 2834 423 2837 573
rect 2842 483 2845 613
rect 2914 596 2917 606
rect 2962 603 2965 636
rect 2914 593 2981 596
rect 2858 533 2861 566
rect 2946 543 2949 576
rect 2930 533 2949 536
rect 2978 526 2981 593
rect 2986 533 2989 596
rect 3002 573 3005 736
rect 2850 506 2853 526
rect 2906 506 2909 526
rect 2850 503 2861 506
rect 2858 396 2861 503
rect 2898 503 2909 506
rect 2898 446 2901 503
rect 2898 443 2909 446
rect 2906 426 2909 443
rect 2906 423 2917 426
rect 2794 393 2805 396
rect 2850 393 2861 396
rect 2766 333 2773 336
rect 2766 256 2769 333
rect 2766 253 2773 256
rect 2770 233 2773 253
rect 2778 206 2781 326
rect 2786 316 2789 336
rect 2794 323 2797 393
rect 2850 376 2853 393
rect 2834 373 2853 376
rect 2810 343 2837 346
rect 2810 323 2813 343
rect 2818 316 2821 326
rect 2786 313 2821 316
rect 2794 233 2805 236
rect 2810 213 2813 226
rect 2778 203 2821 206
rect 2778 133 2781 203
rect 2762 113 2765 126
rect 2770 0 2773 86
rect 2786 0 2789 126
rect 2802 86 2805 156
rect 2826 103 2829 336
rect 2834 326 2837 343
rect 2890 333 2893 346
rect 2834 323 2853 326
rect 2850 156 2853 323
rect 2898 316 2901 416
rect 2906 333 2909 406
rect 2914 396 2917 423
rect 2922 416 2925 526
rect 2946 513 2949 526
rect 2978 523 2989 526
rect 2922 413 2933 416
rect 2914 393 2933 396
rect 2890 313 2901 316
rect 2890 246 2893 313
rect 2914 256 2917 326
rect 2962 313 2965 336
rect 2970 313 2973 326
rect 2986 313 2989 523
rect 2914 253 2925 256
rect 2890 243 2901 246
rect 2898 223 2901 243
rect 2838 153 2853 156
rect 2838 96 2841 153
rect 2834 93 2841 96
rect 2802 83 2813 86
rect 2810 16 2813 83
rect 2834 73 2837 93
rect 2802 13 2813 16
rect 2802 0 2805 13
rect 2850 0 2853 136
rect 2874 133 2877 166
rect 2898 153 2901 216
rect 2922 156 2925 253
rect 2914 153 2925 156
rect 2914 123 2917 153
rect 2946 143 2949 206
rect 2954 196 2957 216
rect 2970 213 2973 226
rect 2954 193 2965 196
rect 2962 136 2965 193
rect 2874 103 2877 116
rect 2922 83 2925 136
rect 2954 133 2965 136
rect 2978 133 2981 306
rect 2954 73 2957 133
rect 2986 83 2989 126
rect 3030 37 3050 3003
rect 3054 13 3074 3027
<< metal3 >>
rect 1401 3022 1470 3027
rect 1945 3012 2030 3017
rect 1201 3002 1390 3007
rect 1385 2997 1390 3002
rect 1457 3002 1934 3007
rect 1457 2997 1462 3002
rect 1385 2992 1462 2997
rect 1929 2997 1934 3002
rect 2041 3002 2806 3007
rect 2041 2997 2046 3002
rect 1929 2992 2046 2997
rect 513 2982 670 2987
rect 513 2977 518 2982
rect 489 2972 518 2977
rect 665 2977 670 2982
rect 665 2972 814 2977
rect 1153 2972 1238 2977
rect 1577 2972 1646 2977
rect 1793 2972 1830 2977
rect 1849 2972 1990 2977
rect 1153 2967 1158 2972
rect 1057 2962 1158 2967
rect 1233 2967 1238 2972
rect 1793 2967 1798 2972
rect 1849 2967 1854 2972
rect 1233 2962 1262 2967
rect 1753 2962 1798 2967
rect 1809 2962 1854 2967
rect 1985 2967 1990 2972
rect 2033 2972 2158 2977
rect 2033 2967 2038 2972
rect 1985 2962 2038 2967
rect 2153 2967 2158 2972
rect 2201 2972 2438 2977
rect 2201 2967 2206 2972
rect 2153 2962 2206 2967
rect 2433 2967 2438 2972
rect 2433 2962 2462 2967
rect 193 2952 286 2957
rect 505 2952 654 2957
rect 1393 2952 1438 2957
rect 1705 2952 1806 2957
rect 1929 2952 2166 2957
rect 2417 2952 2606 2957
rect 2649 2952 2766 2957
rect 2417 2947 2422 2952
rect 673 2942 758 2947
rect 1121 2942 1238 2947
rect 1265 2942 1334 2947
rect 1441 2942 2326 2947
rect 2337 2942 2422 2947
rect 2449 2942 2534 2947
rect 673 2937 678 2942
rect 313 2932 406 2937
rect 465 2932 526 2937
rect 313 2927 318 2932
rect 81 2922 166 2927
rect 289 2922 318 2927
rect 401 2927 406 2932
rect 521 2927 526 2932
rect 593 2932 678 2937
rect 753 2937 758 2942
rect 1265 2937 1270 2942
rect 753 2932 958 2937
rect 1241 2932 1270 2937
rect 1329 2937 1334 2942
rect 1329 2932 1430 2937
rect 1785 2932 1814 2937
rect 1833 2932 2198 2937
rect 593 2927 598 2932
rect 1425 2927 1430 2932
rect 1697 2927 1790 2932
rect 401 2922 502 2927
rect 521 2922 598 2927
rect 641 2922 750 2927
rect 977 2922 1078 2927
rect 1217 2922 1318 2927
rect 1425 2922 1702 2927
rect 1817 2922 1926 2927
rect 2049 2922 2054 2932
rect 2065 2922 2158 2927
rect 2065 2917 2070 2922
rect 721 2912 822 2917
rect 1025 2912 1206 2917
rect 1201 2907 1206 2912
rect 1321 2912 1350 2917
rect 1721 2912 2070 2917
rect 2193 2917 2198 2932
rect 2337 2917 2342 2942
rect 2441 2932 2470 2937
rect 2545 2932 2718 2937
rect 2465 2927 2550 2932
rect 2625 2917 2702 2922
rect 2193 2912 2342 2917
rect 2457 2912 2486 2917
rect 1321 2907 1326 2912
rect 2481 2907 2486 2912
rect 2601 2912 2630 2917
rect 2697 2912 2774 2917
rect 2601 2907 2606 2912
rect 321 2902 390 2907
rect 809 2902 910 2907
rect 1201 2902 1326 2907
rect 1441 2902 1526 2907
rect 1785 2902 1934 2907
rect 2097 2902 2174 2907
rect 2481 2902 2606 2907
rect 2625 2902 2686 2907
rect 1657 2892 1854 2897
rect 1897 2892 2006 2897
rect 249 2882 310 2887
rect 305 2877 310 2882
rect 401 2882 454 2887
rect 401 2877 406 2882
rect 305 2872 406 2877
rect 2025 2872 2326 2877
rect 2025 2867 2030 2872
rect 1753 2862 2030 2867
rect 2321 2867 2326 2872
rect 2321 2862 2454 2867
rect 2017 2852 2134 2857
rect 2273 2852 2310 2857
rect 2449 2852 2454 2862
rect 2529 2862 2678 2867
rect 2273 2847 2278 2852
rect 2529 2847 2534 2862
rect 2673 2857 2678 2862
rect 2673 2852 2758 2857
rect 1865 2842 2278 2847
rect 2505 2842 2534 2847
rect 2753 2847 2758 2852
rect 2753 2842 2782 2847
rect 145 2832 214 2837
rect 313 2832 414 2837
rect 1257 2832 1294 2837
rect 1529 2832 1606 2837
rect 1529 2827 1534 2832
rect 321 2822 422 2827
rect 665 2822 982 2827
rect 1185 2822 1254 2827
rect 1265 2822 1286 2827
rect 1409 2822 1534 2827
rect 1601 2827 1606 2832
rect 1745 2832 1830 2837
rect 1993 2832 2038 2837
rect 2137 2832 2182 2837
rect 2433 2832 2518 2837
rect 2569 2832 2662 2837
rect 1745 2827 1750 2832
rect 1601 2822 1630 2827
rect 1673 2822 1750 2827
rect 1825 2827 1830 2832
rect 2729 2827 2838 2832
rect 1825 2822 1854 2827
rect 1961 2822 2070 2827
rect 2233 2822 2318 2827
rect 2369 2822 2470 2827
rect 2497 2822 2582 2827
rect 2705 2822 2734 2827
rect 2833 2822 2862 2827
rect 1249 2817 1254 2822
rect 2369 2817 2374 2822
rect 121 2812 214 2817
rect 505 2812 598 2817
rect 1249 2812 1462 2817
rect 1457 2807 1462 2812
rect 1841 2812 2062 2817
rect 2145 2812 2374 2817
rect 2737 2812 2774 2817
rect 2785 2812 2894 2817
rect 1841 2807 1846 2812
rect 2393 2807 2478 2812
rect 2513 2807 2646 2812
rect 1361 2802 1446 2807
rect 1457 2802 1646 2807
rect 1761 2802 1846 2807
rect 2073 2802 2142 2807
rect 2353 2802 2398 2807
rect 2473 2802 2518 2807
rect 2641 2802 3014 2807
rect 1169 2797 1254 2802
rect 1857 2797 2078 2802
rect 2137 2797 2142 2802
rect 2249 2797 2358 2802
rect 241 2792 318 2797
rect 441 2792 518 2797
rect 577 2792 702 2797
rect 737 2792 822 2797
rect 865 2792 942 2797
rect 1097 2792 1174 2797
rect 1249 2792 1358 2797
rect 1673 2792 1862 2797
rect 2137 2792 2254 2797
rect 2377 2792 2462 2797
rect 2529 2792 2630 2797
rect 2721 2792 2846 2797
rect 929 2782 1094 2787
rect 929 2777 934 2782
rect 65 2772 446 2777
rect 441 2767 446 2772
rect 649 2772 934 2777
rect 1089 2777 1094 2782
rect 1185 2782 1238 2787
rect 1369 2782 1438 2787
rect 1593 2782 1670 2787
rect 1793 2782 2118 2787
rect 1185 2777 1190 2782
rect 1233 2777 1374 2782
rect 1681 2777 1798 2782
rect 2113 2777 2118 2782
rect 2273 2782 2446 2787
rect 2817 2782 2958 2787
rect 2273 2777 2278 2782
rect 1089 2772 1190 2777
rect 1457 2772 1574 2777
rect 1641 2772 1686 2777
rect 1817 2772 1894 2777
rect 2113 2772 2278 2777
rect 2977 2772 3088 2777
rect 649 2767 654 2772
rect 1457 2767 1462 2772
rect 441 2762 654 2767
rect 1273 2762 1462 2767
rect 1569 2767 1574 2772
rect 1569 2762 1750 2767
rect 1881 2762 2094 2767
rect 2465 2762 2622 2767
rect 1745 2757 1750 2762
rect 2465 2757 2470 2762
rect 65 2752 118 2757
rect 673 2752 734 2757
rect 817 2752 854 2757
rect 1361 2752 1390 2757
rect 1385 2747 1390 2752
rect 1529 2752 1558 2757
rect 1529 2747 1534 2752
rect 89 2742 214 2747
rect 225 2742 302 2747
rect 353 2742 422 2747
rect 761 2742 886 2747
rect 1385 2742 1534 2747
rect 1553 2747 1558 2752
rect 1665 2752 1694 2757
rect 1745 2752 1958 2757
rect 2297 2752 2470 2757
rect 2617 2757 2622 2762
rect 2617 2752 2742 2757
rect 1665 2747 1670 2752
rect 1553 2742 1670 2747
rect 1857 2742 1894 2747
rect 2041 2742 2134 2747
rect 2233 2742 2334 2747
rect 2457 2742 2654 2747
rect 2817 2742 2886 2747
rect 2817 2737 2822 2742
rect 465 2732 494 2737
rect 1241 2732 1326 2737
rect 1737 2732 1854 2737
rect 2313 2732 2366 2737
rect 2769 2732 2822 2737
rect 2881 2737 2886 2742
rect 2881 2732 2910 2737
rect 289 2722 382 2727
rect 465 2707 470 2732
rect 2177 2727 2294 2732
rect 505 2722 614 2727
rect 609 2712 614 2722
rect 1553 2722 1718 2727
rect 1921 2722 2014 2727
rect 2153 2722 2182 2727
rect 2289 2722 2558 2727
rect 2913 2722 3088 2727
rect 1553 2717 1558 2722
rect 1713 2717 1806 2722
rect 1921 2717 1926 2722
rect 1513 2712 1558 2717
rect 1801 2712 1926 2717
rect 2009 2717 2014 2722
rect 2913 2717 2918 2722
rect 2009 2712 2150 2717
rect 2169 2712 2294 2717
rect 2385 2712 2558 2717
rect 2833 2712 2918 2717
rect 145 2702 214 2707
rect 337 2702 470 2707
rect 889 2702 974 2707
rect 1105 2702 1374 2707
rect 1609 2702 1694 2707
rect 1745 2702 1790 2707
rect 2393 2702 2494 2707
rect 2545 2702 2678 2707
rect 1609 2697 1614 2702
rect 1569 2692 1614 2697
rect 1689 2697 1694 2702
rect 1689 2692 1862 2697
rect 1937 2692 1998 2697
rect 2177 2692 2206 2697
rect 2201 2687 2206 2692
rect 2305 2692 2430 2697
rect 2305 2687 2310 2692
rect 1393 2682 1558 2687
rect 1553 2677 1558 2682
rect 1625 2682 1766 2687
rect 2201 2682 2310 2687
rect 1625 2677 1630 2682
rect 1553 2672 1630 2677
rect 1649 2672 1678 2677
rect 1777 2672 2086 2677
rect 1673 2667 1782 2672
rect 641 2662 726 2667
rect 641 2657 646 2662
rect 617 2652 646 2657
rect 721 2657 726 2662
rect 721 2652 982 2657
rect 1473 2652 1566 2657
rect 1633 2652 1694 2657
rect 1713 2652 1918 2657
rect 1473 2647 1478 2652
rect 625 2642 710 2647
rect 1233 2642 1286 2647
rect 1449 2642 1478 2647
rect 1561 2647 1566 2652
rect 1713 2647 1718 2652
rect 1561 2642 1718 2647
rect 1913 2647 1918 2652
rect 2193 2652 2470 2657
rect 2193 2647 2198 2652
rect 1913 2642 2198 2647
rect 2465 2647 2470 2652
rect 2465 2642 2494 2647
rect 2513 2642 2646 2647
rect 1281 2637 1286 2642
rect 89 2632 206 2637
rect 1281 2632 1550 2637
rect 1617 2632 1646 2637
rect 1729 2632 1902 2637
rect 2265 2632 2318 2637
rect 1641 2627 1734 2632
rect 2513 2627 2518 2642
rect 97 2592 102 2627
rect 417 2617 422 2627
rect 601 2622 654 2627
rect 817 2622 854 2627
rect 961 2622 1054 2627
rect 1105 2622 1238 2627
rect 1841 2622 1950 2627
rect 2209 2622 2278 2627
rect 2361 2622 2518 2627
rect 2641 2627 2646 2642
rect 2817 2632 2934 2637
rect 2641 2622 2670 2627
rect 2273 2617 2278 2622
rect 113 2592 118 2617
rect 281 2612 422 2617
rect 1329 2612 1654 2617
rect 1665 2612 1854 2617
rect 2273 2612 2462 2617
rect 2537 2612 2638 2617
rect 1329 2597 1334 2612
rect 1649 2607 1654 2612
rect 1345 2602 1382 2607
rect 1649 2602 1670 2607
rect 1857 2602 2270 2607
rect 2593 2602 2630 2607
rect 201 2592 278 2597
rect 417 2592 510 2597
rect 681 2592 742 2597
rect 1249 2592 1334 2597
rect 1377 2597 1382 2602
rect 1857 2597 1862 2602
rect 2817 2597 2822 2632
rect 3017 2617 3022 2627
rect 3009 2612 3022 2617
rect 3009 2607 3014 2612
rect 3009 2602 3088 2607
rect 3009 2597 3014 2602
rect 1377 2592 1430 2597
rect 1513 2592 1598 2597
rect 1641 2592 1742 2597
rect 1825 2592 1862 2597
rect 2697 2592 2822 2597
rect 2889 2592 3014 2597
rect 1249 2587 1254 2592
rect 1065 2582 1254 2587
rect 1265 2582 1398 2587
rect 1465 2582 1518 2587
rect 1921 2582 1974 2587
rect 2337 2582 2438 2587
rect 2457 2582 2734 2587
rect 1537 2577 1734 2582
rect 2337 2577 2342 2582
rect 1137 2572 1542 2577
rect 1729 2572 1838 2577
rect 1873 2572 1950 2577
rect 1993 2572 2342 2577
rect 2433 2577 2438 2582
rect 2433 2572 2518 2577
rect 2721 2567 2726 2577
rect 953 2562 1054 2567
rect 1049 2557 1054 2562
rect 1177 2562 1206 2567
rect 1217 2562 1718 2567
rect 2353 2562 2510 2567
rect 2641 2562 2726 2567
rect 1177 2557 1182 2562
rect 2641 2557 2646 2562
rect 1049 2552 1182 2557
rect 1337 2552 1550 2557
rect 1601 2552 1814 2557
rect 2089 2552 2198 2557
rect 2417 2552 2446 2557
rect 2521 2552 2646 2557
rect 2441 2547 2526 2552
rect 241 2542 342 2547
rect 849 2542 910 2547
rect 1241 2542 1758 2547
rect 2649 2542 2846 2547
rect 1217 2532 1294 2537
rect 1561 2532 1646 2537
rect 1769 2532 1870 2537
rect 2001 2532 2094 2537
rect 2113 2532 2286 2537
rect 2497 2532 2558 2537
rect 1769 2527 1774 2532
rect 753 2522 822 2527
rect 841 2522 934 2527
rect 1265 2522 1558 2527
rect 1641 2522 1774 2527
rect 1841 2522 1974 2527
rect 1985 2522 2094 2527
rect 2113 2517 2118 2532
rect 457 2512 542 2517
rect 593 2512 630 2517
rect 977 2512 1118 2517
rect 1873 2512 2118 2517
rect 2713 2512 2758 2517
rect 2865 2512 2974 2517
rect 961 2502 1038 2507
rect 1497 2502 1606 2507
rect 1657 2502 1870 2507
rect 1921 2502 1950 2507
rect 1945 2497 1950 2502
rect 2009 2502 2078 2507
rect 2121 2502 2182 2507
rect 2409 2502 2686 2507
rect 2801 2502 2822 2507
rect 2009 2497 2014 2502
rect 1449 2492 1598 2497
rect 1945 2492 2014 2497
rect 1513 2482 1542 2487
rect 1609 2482 1710 2487
rect 1537 2477 1614 2482
rect 993 2472 1166 2477
rect 1553 2462 1702 2467
rect 1729 2462 2094 2467
rect 1729 2457 1734 2462
rect 1601 2452 1734 2457
rect 2089 2457 2094 2462
rect 2089 2452 2118 2457
rect 2177 2452 2454 2457
rect 2737 2452 2814 2457
rect 2833 2452 2958 2457
rect 337 2442 438 2447
rect 337 2437 342 2442
rect 313 2432 342 2437
rect 433 2437 438 2442
rect 1393 2442 1494 2447
rect 1633 2442 1830 2447
rect 1393 2437 1398 2442
rect 433 2432 478 2437
rect 273 2417 278 2427
rect 0 2412 278 2417
rect 321 2412 422 2417
rect 705 2407 710 2437
rect 721 2432 774 2437
rect 945 2432 1094 2437
rect 1369 2432 1398 2437
rect 1489 2437 1494 2442
rect 2177 2437 2182 2452
rect 1489 2432 1630 2437
rect 1649 2432 2182 2437
rect 2449 2437 2454 2452
rect 2833 2447 2838 2452
rect 2617 2442 2710 2447
rect 2801 2442 2838 2447
rect 2953 2447 2958 2452
rect 2953 2442 2982 2447
rect 2449 2432 2526 2437
rect 2657 2432 2990 2437
rect 769 2427 774 2432
rect 769 2422 798 2427
rect 865 2422 974 2427
rect 1185 2422 1214 2427
rect 1617 2422 1646 2427
rect 1641 2417 1646 2422
rect 1729 2422 1806 2427
rect 2193 2422 2446 2427
rect 2625 2422 2702 2427
rect 1729 2417 1734 2422
rect 2025 2417 2126 2422
rect 2193 2417 2198 2422
rect 2833 2417 2982 2422
rect 937 2412 966 2417
rect 1361 2412 1478 2417
rect 1641 2412 1734 2417
rect 1857 2412 2030 2417
rect 2121 2412 2198 2417
rect 2417 2412 2486 2417
rect 2809 2412 2838 2417
rect 2977 2412 3088 2417
rect 537 2402 582 2407
rect 705 2402 742 2407
rect 785 2402 822 2407
rect 577 2397 582 2402
rect 961 2397 966 2412
rect 993 2402 1166 2407
rect 1193 2402 1438 2407
rect 1449 2402 1510 2407
rect 1753 2402 1838 2407
rect 993 2397 998 2402
rect 577 2392 694 2397
rect 689 2387 694 2392
rect 777 2392 806 2397
rect 961 2392 998 2397
rect 1161 2397 1166 2402
rect 1433 2397 1438 2402
rect 1161 2392 1422 2397
rect 1433 2392 1486 2397
rect 1505 2392 1510 2402
rect 1857 2397 1862 2412
rect 2041 2402 2110 2407
rect 2609 2402 2750 2407
rect 2833 2402 2966 2407
rect 1545 2392 1862 2397
rect 1889 2392 2030 2397
rect 2121 2392 2262 2397
rect 2841 2392 2886 2397
rect 777 2387 782 2392
rect 2025 2387 2126 2392
rect 689 2382 782 2387
rect 985 2382 1294 2387
rect 1457 2382 1558 2387
rect 2345 2382 2686 2387
rect 2761 2382 2910 2387
rect 521 2372 622 2377
rect 1161 2372 1798 2377
rect 1033 2367 1142 2372
rect 1793 2367 1798 2372
rect 2089 2372 2150 2377
rect 2209 2372 2302 2377
rect 2665 2372 2694 2377
rect 2089 2367 2094 2372
rect 873 2362 966 2367
rect 1009 2362 1038 2367
rect 1137 2362 1278 2367
rect 1513 2362 1542 2367
rect 873 2357 878 2362
rect 73 2352 158 2357
rect 529 2352 646 2357
rect 849 2352 878 2357
rect 961 2357 966 2362
rect 1537 2357 1542 2362
rect 1745 2362 1774 2367
rect 1793 2362 2094 2367
rect 2657 2362 2790 2367
rect 1745 2357 1750 2362
rect 2657 2357 2662 2362
rect 961 2352 1158 2357
rect 1153 2347 1158 2352
rect 1217 2352 1246 2357
rect 1537 2352 1750 2357
rect 2217 2352 2662 2357
rect 2673 2352 2974 2357
rect 1217 2347 1222 2352
rect 545 2342 630 2347
rect 681 2342 790 2347
rect 1025 2342 1126 2347
rect 1153 2342 1222 2347
rect 1321 2342 1494 2347
rect 873 2332 1038 2337
rect 1321 2327 1326 2342
rect 1489 2337 1494 2342
rect 2113 2342 2174 2347
rect 2617 2342 2670 2347
rect 2689 2342 2766 2347
rect 2857 2342 2958 2347
rect 2113 2337 2118 2342
rect 1489 2332 2030 2337
rect 2049 2332 2118 2337
rect 2193 2332 2606 2337
rect 1041 2322 1326 2327
rect 2025 2327 2030 2332
rect 2193 2327 2198 2332
rect 2025 2322 2198 2327
rect 2601 2327 2606 2332
rect 2689 2327 2694 2342
rect 2737 2332 2854 2337
rect 3017 2327 3022 2337
rect 2601 2322 2694 2327
rect 2905 2322 3088 2327
rect 2465 2317 2558 2322
rect 929 2312 1046 2317
rect 1041 2307 1046 2312
rect 1129 2312 1158 2317
rect 1337 2312 1614 2317
rect 1713 2312 1814 2317
rect 1833 2312 1942 2317
rect 1961 2312 2342 2317
rect 2441 2312 2470 2317
rect 2553 2312 2582 2317
rect 2721 2312 2742 2317
rect 1129 2307 1134 2312
rect 377 2302 454 2307
rect 513 2302 822 2307
rect 1041 2302 1134 2307
rect 1153 2302 1158 2312
rect 1833 2307 1838 2312
rect 1449 2302 1486 2307
rect 1537 2302 1566 2307
rect 817 2297 822 2302
rect 1561 2297 1566 2302
rect 1625 2302 1702 2307
rect 1625 2297 1630 2302
rect 817 2292 918 2297
rect 913 2287 918 2292
rect 993 2292 1022 2297
rect 1561 2292 1630 2297
rect 1697 2297 1702 2302
rect 1761 2302 1838 2307
rect 1937 2307 1942 2312
rect 1937 2302 2182 2307
rect 1761 2297 1766 2302
rect 2177 2297 2182 2302
rect 2353 2302 2382 2307
rect 2465 2302 2574 2307
rect 2609 2302 2894 2307
rect 2353 2297 2358 2302
rect 1697 2292 1766 2297
rect 1809 2292 2158 2297
rect 2177 2292 2358 2297
rect 2889 2297 2894 2302
rect 2969 2302 3088 2307
rect 2969 2297 2974 2302
rect 2889 2292 2974 2297
rect 993 2287 998 2292
rect 697 2282 726 2287
rect 721 2277 726 2282
rect 793 2282 822 2287
rect 913 2282 998 2287
rect 1785 2282 1910 2287
rect 1921 2282 2062 2287
rect 2521 2282 2590 2287
rect 793 2277 798 2282
rect 2585 2277 2590 2282
rect 2705 2282 2734 2287
rect 2705 2277 2710 2282
rect 721 2272 798 2277
rect 1057 2272 2566 2277
rect 2585 2272 2710 2277
rect 2025 2262 2094 2267
rect 2521 2262 2542 2267
rect 1617 2257 2006 2262
rect 1593 2252 1622 2257
rect 2001 2252 2214 2257
rect 385 2242 462 2247
rect 993 2242 1582 2247
rect 1577 2237 1582 2242
rect 1649 2242 2054 2247
rect 2305 2242 2606 2247
rect 2961 2242 3088 2247
rect 1649 2237 1654 2242
rect 2961 2237 2966 2242
rect 313 2232 350 2237
rect 921 2232 1006 2237
rect 1577 2232 1654 2237
rect 1737 2232 1806 2237
rect 1993 2232 2102 2237
rect 2697 2232 2966 2237
rect 1825 2227 1998 2232
rect 177 2222 214 2227
rect 177 2217 182 2222
rect 865 2217 870 2227
rect 897 2222 974 2227
rect 1153 2222 1270 2227
rect 1673 2222 1830 2227
rect 2017 2222 2046 2227
rect 2113 2222 2366 2227
rect 2425 2222 2470 2227
rect 1153 2217 1158 2222
rect 0 2212 182 2217
rect 225 2212 494 2217
rect 521 2212 630 2217
rect 865 2212 886 2217
rect 881 2207 886 2212
rect 1017 2212 1158 2217
rect 1553 2212 1654 2217
rect 1681 2212 1950 2217
rect 2017 2212 2022 2222
rect 2041 2217 2118 2222
rect 2465 2217 2470 2222
rect 2465 2212 2718 2217
rect 1017 2207 1022 2212
rect 1553 2207 1558 2212
rect 881 2202 1022 2207
rect 1193 2202 1222 2207
rect 1217 2197 1222 2202
rect 1281 2202 1310 2207
rect 1401 2202 1454 2207
rect 1537 2202 1558 2207
rect 1649 2207 1654 2212
rect 1649 2202 1718 2207
rect 1881 2202 2270 2207
rect 2321 2202 2494 2207
rect 1281 2197 1286 2202
rect 337 2192 358 2197
rect 1217 2192 1286 2197
rect 1537 2192 1542 2202
rect 1713 2197 1886 2202
rect 1561 2192 1694 2197
rect 1905 2192 2054 2197
rect 2289 2192 2342 2197
rect 2513 2192 2566 2197
rect 217 2182 334 2187
rect 617 2182 774 2187
rect 1481 2182 1558 2187
rect 1761 2182 1806 2187
rect 1993 2182 2182 2187
rect 2313 2182 2454 2187
rect 2737 2182 2766 2187
rect 81 2172 190 2177
rect 1417 2172 1470 2177
rect 1889 2172 1958 2177
rect 2121 2172 2230 2177
rect 2241 2172 2422 2177
rect 369 2162 454 2167
rect 369 2157 374 2162
rect 345 2152 374 2157
rect 449 2157 454 2162
rect 1081 2162 1166 2167
rect 1649 2162 1702 2167
rect 1713 2162 2150 2167
rect 2185 2162 2222 2167
rect 2233 2162 2358 2167
rect 2481 2162 2718 2167
rect 1081 2157 1086 2162
rect 449 2152 478 2157
rect 1057 2152 1086 2157
rect 1161 2157 1166 2162
rect 2481 2157 2486 2162
rect 1161 2152 1190 2157
rect 1449 2152 1654 2157
rect 1857 2152 1950 2157
rect 2217 2152 2486 2157
rect 2713 2157 2718 2162
rect 2737 2157 2742 2182
rect 2713 2152 2782 2157
rect 2849 2152 2926 2157
rect 1649 2147 1654 2152
rect 81 2142 294 2147
rect 905 2142 1038 2147
rect 1649 2142 1734 2147
rect 1753 2142 2206 2147
rect 81 2137 86 2142
rect 905 2137 910 2142
rect 0 2132 86 2137
rect 281 2132 726 2137
rect 881 2132 910 2137
rect 1033 2137 1038 2142
rect 1729 2137 1734 2142
rect 2201 2137 2206 2142
rect 2273 2142 2302 2147
rect 2713 2142 2862 2147
rect 2273 2137 2278 2142
rect 1033 2132 1150 2137
rect 1433 2132 1478 2137
rect 1729 2132 1758 2137
rect 2113 2132 2142 2137
rect 2201 2132 2278 2137
rect 2409 2132 2702 2137
rect 1753 2127 1934 2132
rect 2113 2127 2118 2132
rect 1321 2122 1358 2127
rect 1593 2122 1630 2127
rect 1929 2122 2118 2127
rect 2697 2127 2702 2132
rect 2697 2122 3088 2127
rect 905 2117 990 2122
rect 0 2112 30 2117
rect 25 2107 30 2112
rect 97 2112 230 2117
rect 345 2112 622 2117
rect 881 2112 910 2117
rect 985 2112 1246 2117
rect 1329 2112 1422 2117
rect 1537 2112 1566 2117
rect 1641 2112 1910 2117
rect 2161 2112 2246 2117
rect 2265 2112 2390 2117
rect 97 2107 102 2112
rect 1561 2107 1646 2112
rect 2265 2107 2270 2112
rect 25 2102 102 2107
rect 617 2102 838 2107
rect 873 2102 974 2107
rect 1089 2102 1174 2107
rect 129 2092 166 2097
rect 977 2092 1150 2097
rect 1169 2087 1174 2102
rect 1361 2102 1526 2107
rect 1361 2087 1366 2102
rect 1521 2097 1526 2102
rect 1713 2102 1790 2107
rect 1921 2102 2270 2107
rect 2385 2107 2390 2112
rect 2385 2102 2846 2107
rect 1713 2097 1718 2102
rect 1785 2097 1926 2102
rect 1449 2092 1502 2097
rect 1521 2092 1718 2097
rect 1737 2092 1766 2097
rect 2105 2092 2174 2097
rect 2857 2092 2918 2097
rect 2913 2087 2918 2092
rect 417 2082 606 2087
rect 601 2077 606 2082
rect 937 2082 1030 2087
rect 1169 2082 1366 2087
rect 1385 2082 1414 2087
rect 937 2077 942 2082
rect 1409 2077 1414 2082
rect 1833 2082 2094 2087
rect 1833 2077 1838 2082
rect 601 2072 942 2077
rect 961 2072 1046 2077
rect 1409 2072 1838 2077
rect 2089 2077 2094 2082
rect 2185 2082 2910 2087
rect 2913 2082 3088 2087
rect 2185 2077 2190 2082
rect 2089 2072 2190 2077
rect 2617 2072 2646 2077
rect 2641 2067 2646 2072
rect 2825 2072 2886 2077
rect 2905 2072 2910 2082
rect 2825 2067 2830 2072
rect 2641 2062 2830 2067
rect 2881 2067 2886 2072
rect 2881 2062 2934 2067
rect 1857 2052 2326 2057
rect 2377 2052 2558 2057
rect 1425 2042 1494 2047
rect 1721 2042 1894 2047
rect 2625 2042 2814 2047
rect 1425 2037 1430 2042
rect 385 2032 462 2037
rect 793 2032 958 2037
rect 1113 2032 1430 2037
rect 1489 2037 1494 2042
rect 1489 2032 1678 2037
rect 1737 2032 1838 2037
rect 129 2022 166 2027
rect 281 2022 342 2027
rect 2049 2022 2166 2027
rect 2417 2022 2758 2027
rect 2833 2022 2934 2027
rect 2049 2017 2054 2022
rect 665 2012 758 2017
rect 1441 2012 1478 2017
rect 1545 2012 1614 2017
rect 1873 2012 1974 2017
rect 2025 2012 2054 2017
rect 2161 2017 2166 2022
rect 2833 2017 2838 2022
rect 2161 2012 2342 2017
rect 2729 2012 2838 2017
rect 2929 2017 2934 2022
rect 2929 2012 2958 2017
rect 1545 2007 1550 2012
rect 0 2002 302 2007
rect 841 2002 950 2007
rect 961 2002 998 2007
rect 1225 2002 1262 2007
rect 1521 2002 1550 2007
rect 1609 2007 1614 2012
rect 1609 2002 1638 2007
rect 2793 1997 2910 2002
rect 3083 1997 3088 2017
rect 737 1992 766 1997
rect 1033 1992 1078 1997
rect 1401 1992 1542 1997
rect 1577 1992 1750 1997
rect 1929 1992 2150 1997
rect 2289 1992 2366 1997
rect 2577 1992 2798 1997
rect 2905 1992 3088 1997
rect 81 1982 198 1987
rect 785 1982 982 1987
rect 1105 1982 1246 1987
rect 1265 1982 1670 1987
rect 1825 1982 1910 1987
rect 785 1977 790 1982
rect 713 1972 790 1977
rect 977 1977 982 1982
rect 1265 1977 1270 1982
rect 977 1972 1270 1977
rect 809 1967 902 1972
rect 1401 1967 1662 1972
rect 1825 1967 1830 1982
rect 1905 1977 1910 1982
rect 2169 1982 2270 1987
rect 2809 1982 2894 1987
rect 2169 1977 2174 1982
rect 1905 1972 2030 1977
rect 2129 1972 2174 1977
rect 2265 1977 2270 1982
rect 2265 1972 2342 1977
rect 2513 1972 2582 1977
rect 2513 1967 2518 1972
rect 0 1962 278 1967
rect 721 1962 814 1967
rect 897 1962 966 1967
rect 1377 1962 1406 1967
rect 1657 1962 1854 1967
rect 2081 1962 2446 1967
rect 2489 1962 2518 1967
rect 2577 1967 2582 1972
rect 2577 1962 2870 1967
rect 985 1957 1238 1962
rect 745 1952 870 1957
rect 905 1952 990 1957
rect 1233 1952 1646 1957
rect 1873 1952 2270 1957
rect 2353 1952 2438 1957
rect 2537 1952 2670 1957
rect 1737 1947 1814 1952
rect 2265 1947 2358 1952
rect 2433 1947 2518 1952
rect 2721 1947 2822 1952
rect 97 1942 206 1947
rect 753 1942 870 1947
rect 945 1942 1158 1947
rect 1401 1942 1430 1947
rect 1505 1942 1550 1947
rect 1657 1942 1742 1947
rect 1809 1942 1838 1947
rect 2097 1942 2198 1947
rect 2377 1942 2414 1947
rect 2513 1942 2542 1947
rect 2681 1942 2726 1947
rect 2817 1942 2974 1947
rect 2993 1942 3088 1947
rect 1217 1937 1406 1942
rect 1545 1937 1662 1942
rect 1953 1937 2062 1942
rect 2537 1937 2686 1942
rect 2993 1937 2998 1942
rect 721 1932 742 1937
rect 721 1927 726 1932
rect 705 1922 726 1927
rect 737 1927 742 1932
rect 833 1932 1022 1937
rect 833 1927 838 1932
rect 1017 1927 1022 1932
rect 1217 1927 1222 1937
rect 1497 1932 1526 1937
rect 1521 1927 1526 1932
rect 1753 1932 1958 1937
rect 2057 1932 2086 1937
rect 1753 1927 1758 1932
rect 737 1922 838 1927
rect 857 1922 886 1927
rect 881 1917 886 1922
rect 969 1922 998 1927
rect 1017 1922 1222 1927
rect 1257 1922 1494 1927
rect 1521 1922 1758 1927
rect 1777 1922 1806 1927
rect 1833 1922 1862 1927
rect 1969 1922 2046 1927
rect 969 1917 974 1922
rect 249 1912 358 1917
rect 881 1912 974 1917
rect 1489 1907 1494 1922
rect 1777 1907 1782 1922
rect 1857 1917 1974 1922
rect 2081 1917 2086 1932
rect 2209 1932 2366 1937
rect 2737 1932 2806 1937
rect 2873 1932 2998 1937
rect 2209 1917 2214 1932
rect 2361 1927 2470 1932
rect 2465 1922 2566 1927
rect 2585 1922 2718 1927
rect 2969 1922 3088 1927
rect 2585 1917 2590 1922
rect 2081 1912 2214 1917
rect 2425 1912 2590 1917
rect 2713 1917 2718 1922
rect 2713 1912 2742 1917
rect 1081 1902 1126 1907
rect 1345 1902 1470 1907
rect 1489 1902 1782 1907
rect 1841 1902 1942 1907
rect 2241 1902 2974 1907
rect 1857 1892 1894 1897
rect 2145 1892 2230 1897
rect 2145 1887 2150 1892
rect 1 1877 6 1887
rect 873 1882 1350 1887
rect 1825 1882 2150 1887
rect 2225 1887 2230 1892
rect 2241 1887 2246 1902
rect 2969 1897 2974 1902
rect 3057 1902 3088 1907
rect 3057 1897 3062 1902
rect 2393 1892 2422 1897
rect 2225 1882 2246 1887
rect 2417 1887 2422 1892
rect 2513 1892 2542 1897
rect 2657 1892 2686 1897
rect 2513 1887 2518 1892
rect 2417 1882 2518 1887
rect 2681 1877 2686 1892
rect 2921 1892 2950 1897
rect 2969 1892 3062 1897
rect 2921 1877 2926 1892
rect 0 1872 6 1877
rect 1281 1872 1358 1877
rect 1385 1872 1774 1877
rect 2161 1872 2222 1877
rect 2681 1872 2926 1877
rect 0 1857 5 1872
rect 1385 1867 1390 1872
rect 169 1862 238 1867
rect 1001 1862 1086 1867
rect 1361 1862 1390 1867
rect 1769 1867 1774 1872
rect 1769 1862 1910 1867
rect 1001 1857 1006 1862
rect 0 1852 582 1857
rect 713 1852 822 1857
rect 713 1847 718 1852
rect 121 1842 150 1847
rect 145 1837 150 1842
rect 225 1842 302 1847
rect 689 1842 718 1847
rect 817 1847 822 1852
rect 865 1852 958 1857
rect 977 1852 1006 1857
rect 1081 1857 1086 1862
rect 1905 1857 1910 1862
rect 1081 1852 1270 1857
rect 1409 1852 1718 1857
rect 1905 1852 1926 1857
rect 2241 1852 2478 1857
rect 2497 1852 2590 1857
rect 865 1847 870 1852
rect 817 1842 870 1847
rect 953 1847 958 1852
rect 1409 1847 1414 1852
rect 953 1842 1414 1847
rect 1713 1847 1718 1852
rect 1713 1842 1742 1847
rect 1801 1842 2014 1847
rect 2073 1842 2214 1847
rect 225 1837 230 1842
rect 1433 1837 1518 1842
rect 2241 1837 2246 1852
rect 2473 1842 2478 1852
rect 2609 1842 2694 1847
rect 2473 1837 2614 1842
rect 2689 1837 2694 1842
rect 145 1832 230 1837
rect 857 1832 990 1837
rect 1017 1832 1118 1837
rect 1209 1832 1278 1837
rect 1401 1832 1438 1837
rect 1513 1832 2246 1837
rect 2689 1832 2710 1837
rect 2769 1832 2918 1837
rect 2705 1827 2710 1832
rect 249 1822 294 1827
rect 553 1822 726 1827
rect 737 1822 846 1827
rect 929 1822 1502 1827
rect 1825 1822 1894 1827
rect 1993 1822 2270 1827
rect 2369 1822 2686 1827
rect 2705 1822 2734 1827
rect 2841 1822 2870 1827
rect 1713 1817 1782 1822
rect 217 1812 278 1817
rect 769 1812 878 1817
rect 1057 1812 1238 1817
rect 1289 1812 1534 1817
rect 1569 1812 1670 1817
rect 1689 1812 1718 1817
rect 1777 1812 2054 1817
rect 2153 1812 2190 1817
rect 2369 1812 2374 1822
rect 2729 1817 2846 1822
rect 2385 1812 2414 1817
rect 2617 1812 2702 1817
rect 1569 1807 1574 1812
rect 297 1802 542 1807
rect 537 1797 542 1802
rect 641 1802 1446 1807
rect 1545 1802 1574 1807
rect 1665 1807 1670 1812
rect 2049 1807 2158 1812
rect 2385 1807 2390 1812
rect 1665 1802 1766 1807
rect 1865 1802 2030 1807
rect 2177 1802 2390 1807
rect 2497 1802 2598 1807
rect 2721 1802 2774 1807
rect 2841 1802 2982 1807
rect 641 1797 646 1802
rect 1441 1797 1550 1802
rect 2497 1797 2502 1802
rect 2593 1797 2726 1802
rect 537 1792 646 1797
rect 825 1792 1422 1797
rect 1585 1792 1630 1797
rect 1657 1792 1790 1797
rect 1809 1792 2502 1797
rect 2753 1792 2862 1797
rect 2753 1787 2758 1792
rect 665 1782 702 1787
rect 697 1777 702 1782
rect 825 1782 1134 1787
rect 1265 1782 1486 1787
rect 1569 1782 1638 1787
rect 1849 1782 1886 1787
rect 1913 1782 1990 1787
rect 2001 1782 2086 1787
rect 2193 1782 2230 1787
rect 2305 1782 2366 1787
rect 2385 1782 2414 1787
rect 2513 1782 2646 1787
rect 2673 1782 2758 1787
rect 825 1777 830 1782
rect 1129 1777 1270 1782
rect 89 1772 486 1777
rect 697 1772 830 1777
rect 921 1772 1014 1777
rect 1289 1772 1374 1777
rect 1497 1772 1558 1777
rect 1649 1772 1742 1777
rect 89 1767 94 1772
rect 0 1762 94 1767
rect 481 1767 486 1772
rect 1033 1767 1110 1772
rect 1369 1767 1502 1772
rect 1553 1767 1654 1772
rect 1737 1767 1742 1772
rect 1833 1772 1862 1777
rect 1881 1772 1942 1777
rect 1833 1767 1838 1772
rect 481 1762 510 1767
rect 873 1762 1038 1767
rect 1105 1762 1278 1767
rect 1737 1762 1838 1767
rect 1937 1767 1942 1772
rect 2073 1772 2126 1777
rect 2073 1767 2078 1772
rect 1937 1762 2078 1767
rect 2121 1767 2126 1772
rect 2193 1767 2198 1782
rect 2385 1777 2390 1782
rect 2217 1772 2246 1777
rect 2121 1762 2198 1767
rect 2241 1767 2246 1772
rect 2369 1772 2406 1777
rect 2369 1767 2374 1772
rect 2241 1762 2374 1767
rect 2401 1767 2406 1772
rect 2513 1772 2582 1777
rect 2513 1767 2518 1772
rect 2401 1762 2518 1767
rect 2577 1767 2582 1772
rect 2697 1772 2790 1777
rect 2697 1767 2702 1772
rect 2577 1762 2702 1767
rect 2721 1762 2958 1767
rect 2985 1762 3088 1767
rect 1273 1757 1350 1762
rect 545 1752 678 1757
rect 849 1752 1094 1757
rect 1345 1747 1350 1757
rect 1465 1752 1718 1757
rect 2673 1747 2822 1752
rect 0 1742 470 1747
rect 825 1742 910 1747
rect 961 1742 1014 1747
rect 1081 1742 1134 1747
rect 1265 1742 1326 1747
rect 1345 1742 1478 1747
rect 2537 1742 2630 1747
rect 2649 1742 2678 1747
rect 2817 1742 3088 1747
rect 2537 1737 2542 1742
rect 1177 1732 1262 1737
rect 1497 1732 1646 1737
rect 2393 1732 2542 1737
rect 2625 1737 2630 1742
rect 2625 1732 2806 1737
rect 2801 1727 2806 1732
rect 137 1722 326 1727
rect 961 1722 1126 1727
rect 1185 1722 1214 1727
rect 137 1717 142 1722
rect 0 1712 142 1717
rect 321 1717 326 1722
rect 1209 1717 1214 1722
rect 1273 1722 1390 1727
rect 1585 1722 1694 1727
rect 1897 1722 1982 1727
rect 2105 1722 2174 1727
rect 2297 1722 2790 1727
rect 2801 1722 2854 1727
rect 1273 1717 1278 1722
rect 2785 1717 2790 1722
rect 2849 1717 2854 1722
rect 3057 1722 3088 1727
rect 3057 1717 3062 1722
rect 321 1712 478 1717
rect 649 1712 846 1717
rect 1209 1712 1278 1717
rect 1361 1712 1942 1717
rect 2481 1712 2542 1717
rect 2537 1707 2542 1712
rect 2609 1712 2638 1717
rect 2785 1712 2830 1717
rect 2849 1712 3062 1717
rect 2609 1707 2614 1712
rect 153 1702 310 1707
rect 1601 1702 1686 1707
rect 1857 1702 1966 1707
rect 2121 1702 2518 1707
rect 2537 1702 2614 1707
rect 2785 1702 2822 1707
rect 0 1692 142 1697
rect 137 1687 142 1692
rect 265 1692 622 1697
rect 833 1692 1022 1697
rect 1057 1692 1262 1697
rect 265 1687 270 1692
rect 1057 1687 1062 1692
rect 137 1682 270 1687
rect 1033 1682 1062 1687
rect 1257 1687 1262 1692
rect 1417 1692 1582 1697
rect 1417 1687 1422 1692
rect 1577 1687 1710 1692
rect 2513 1687 2518 1702
rect 2785 1697 2790 1702
rect 2649 1692 2790 1697
rect 2649 1687 2654 1692
rect 1257 1682 1422 1687
rect 1705 1682 2494 1687
rect 2513 1682 2654 1687
rect 2873 1682 2934 1687
rect 2929 1677 2934 1682
rect 0 1672 94 1677
rect 89 1667 94 1672
rect 289 1672 342 1677
rect 289 1667 294 1672
rect 89 1662 294 1667
rect 337 1667 342 1672
rect 417 1672 446 1677
rect 825 1672 1030 1677
rect 1433 1672 1694 1677
rect 2809 1672 2902 1677
rect 2929 1672 3088 1677
rect 417 1667 422 1672
rect 337 1662 422 1667
rect 1025 1667 1030 1672
rect 1025 1662 1246 1667
rect 1529 1662 1558 1667
rect 1553 1657 1558 1662
rect 1633 1662 1662 1667
rect 2977 1662 3014 1667
rect 1633 1657 1638 1662
rect 721 1652 806 1657
rect 1553 1652 1638 1657
rect 1745 1652 2846 1657
rect 721 1647 726 1652
rect 0 1642 70 1647
rect 497 1642 566 1647
rect 697 1642 726 1647
rect 801 1647 806 1652
rect 2841 1647 2846 1652
rect 2977 1647 2982 1662
rect 801 1642 974 1647
rect 1121 1642 1158 1647
rect 497 1637 502 1642
rect 369 1632 414 1637
rect 473 1632 502 1637
rect 561 1637 566 1642
rect 561 1632 678 1637
rect 1089 1632 1150 1637
rect 761 1627 942 1632
rect 2353 1627 2358 1647
rect 2841 1642 2982 1647
rect 2569 1632 2686 1637
rect 2705 1632 2798 1637
rect 2705 1627 2710 1632
rect 737 1622 766 1627
rect 937 1622 966 1627
rect 993 1622 1206 1627
rect 1297 1622 1358 1627
rect 1705 1622 1806 1627
rect 2041 1622 2118 1627
rect 2337 1622 2630 1627
rect 2665 1622 2710 1627
rect 2793 1627 2798 1632
rect 2793 1622 2822 1627
rect 993 1617 998 1622
rect 25 1612 118 1617
rect 385 1612 550 1617
rect 753 1612 998 1617
rect 1089 1612 1158 1617
rect 1321 1612 1382 1617
rect 1609 1612 1718 1617
rect 2033 1612 2062 1617
rect 2617 1612 2862 1617
rect 25 1607 30 1612
rect 0 1602 30 1607
rect 113 1597 118 1612
rect 129 1602 198 1607
rect 217 1602 366 1607
rect 217 1597 222 1602
rect 113 1592 222 1597
rect 361 1597 366 1602
rect 417 1602 462 1607
rect 545 1602 622 1607
rect 721 1602 990 1607
rect 1025 1602 1134 1607
rect 1401 1602 1526 1607
rect 1545 1602 1758 1607
rect 2097 1602 2182 1607
rect 2409 1602 2694 1607
rect 417 1597 422 1602
rect 1401 1597 1406 1602
rect 361 1592 422 1597
rect 729 1592 822 1597
rect 1153 1592 1190 1597
rect 1369 1592 1406 1597
rect 1521 1597 1526 1602
rect 1521 1592 1550 1597
rect 1769 1592 1830 1597
rect 2305 1592 2390 1597
rect 2681 1592 2814 1597
rect 241 1587 342 1592
rect 441 1587 526 1592
rect 849 1587 974 1592
rect 1545 1587 1654 1592
rect 1769 1587 1774 1592
rect 2305 1587 2310 1592
rect 0 1582 246 1587
rect 337 1582 446 1587
rect 521 1582 718 1587
rect 833 1582 854 1587
rect 969 1582 998 1587
rect 1257 1582 1350 1587
rect 1441 1582 1502 1587
rect 1649 1582 1774 1587
rect 2281 1582 2310 1587
rect 2385 1587 2390 1592
rect 2385 1582 2430 1587
rect 2625 1582 2694 1587
rect 713 1577 838 1582
rect 1257 1577 1262 1582
rect 225 1572 510 1577
rect 865 1572 1262 1577
rect 1345 1577 1350 1582
rect 1345 1572 1582 1577
rect 2289 1572 2374 1577
rect 2441 1572 3088 1577
rect 105 1567 206 1572
rect 2369 1567 2446 1572
rect 0 1562 70 1567
rect 81 1562 110 1567
rect 201 1562 598 1567
rect 617 1562 846 1567
rect 1337 1562 1454 1567
rect 1497 1562 1630 1567
rect 2657 1562 2742 1567
rect 65 1557 70 1562
rect 617 1557 622 1562
rect 65 1552 622 1557
rect 841 1557 846 1562
rect 1017 1557 1094 1562
rect 841 1552 886 1557
rect 929 1552 1022 1557
rect 1089 1552 1158 1557
rect 1273 1552 1462 1557
rect 1657 1552 1814 1557
rect 1657 1547 1662 1552
rect 0 1542 54 1547
rect 49 1537 54 1542
rect 113 1542 270 1547
rect 633 1542 710 1547
rect 721 1542 862 1547
rect 1033 1542 1078 1547
rect 1281 1542 1414 1547
rect 1441 1542 1510 1547
rect 1633 1542 1662 1547
rect 1809 1547 1814 1552
rect 1857 1552 2006 1557
rect 1809 1542 1838 1547
rect 113 1537 118 1542
rect 265 1537 638 1542
rect 49 1532 118 1537
rect 161 1532 246 1537
rect 705 1532 710 1542
rect 1857 1537 1862 1552
rect 2001 1537 2006 1552
rect 2289 1552 2478 1557
rect 2289 1547 2294 1552
rect 2105 1542 2294 1547
rect 2473 1547 2478 1552
rect 2897 1552 2966 1557
rect 2897 1547 2902 1552
rect 2473 1542 2502 1547
rect 2561 1542 2606 1547
rect 2673 1542 2798 1547
rect 2873 1542 2902 1547
rect 2961 1547 2966 1552
rect 2961 1542 3088 1547
rect 945 1532 1054 1537
rect 1697 1532 1790 1537
rect 1817 1532 1862 1537
rect 1881 1532 1966 1537
rect 2001 1532 2150 1537
rect 705 1527 838 1532
rect 1217 1527 1318 1532
rect 1697 1527 1702 1532
rect 137 1522 654 1527
rect 833 1522 1006 1527
rect 1057 1522 1222 1527
rect 1313 1522 1702 1527
rect 1785 1527 1790 1532
rect 1881 1527 1886 1532
rect 1785 1522 1886 1527
rect 1961 1527 1966 1532
rect 1961 1522 1990 1527
rect 1057 1517 1062 1522
rect 2145 1517 2150 1532
rect 2305 1532 2502 1537
rect 2801 1532 2862 1537
rect 2921 1532 2950 1537
rect 2305 1517 2310 1532
rect 2857 1527 2926 1532
rect 2497 1522 2534 1527
rect 2529 1517 2534 1522
rect 2617 1522 2678 1527
rect 3057 1522 3088 1527
rect 2617 1517 2622 1522
rect 3057 1517 3062 1522
rect 0 1512 54 1517
rect 65 1512 302 1517
rect 737 1512 1062 1517
rect 1233 1512 1302 1517
rect 1713 1512 1814 1517
rect 1897 1512 1958 1517
rect 2145 1512 2310 1517
rect 2329 1512 2510 1517
rect 2529 1512 2622 1517
rect 2729 1512 2878 1517
rect 49 1507 54 1512
rect 2873 1507 2878 1512
rect 2977 1512 3062 1517
rect 2977 1507 2982 1512
rect 49 1502 766 1507
rect 777 1502 1102 1507
rect 1609 1502 1782 1507
rect 2873 1502 2982 1507
rect 0 1492 30 1497
rect 937 1492 1110 1497
rect 1217 1492 1590 1497
rect 1721 1492 1822 1497
rect 2337 1492 2430 1497
rect 25 1487 942 1492
rect 1217 1487 1222 1492
rect 1049 1482 1222 1487
rect 1585 1487 1590 1492
rect 1585 1482 1614 1487
rect 0 1472 702 1477
rect 753 1472 918 1477
rect 937 1472 1502 1477
rect 753 1467 758 1472
rect 729 1462 758 1467
rect 913 1467 918 1472
rect 1529 1467 1670 1472
rect 913 1462 1270 1467
rect 169 1457 238 1462
rect 145 1452 174 1457
rect 233 1452 942 1457
rect 1145 1452 1174 1457
rect 145 1447 150 1452
rect 937 1447 1046 1452
rect 1145 1447 1150 1452
rect 0 1442 150 1447
rect 169 1442 222 1447
rect 1041 1442 1150 1447
rect 1265 1447 1270 1462
rect 1449 1462 1534 1467
rect 1665 1462 2422 1467
rect 1449 1447 1454 1462
rect 2417 1457 2422 1462
rect 1545 1452 1654 1457
rect 2417 1452 3088 1457
rect 1265 1442 1454 1447
rect 1769 1442 1806 1447
rect 2201 1442 2270 1447
rect 513 1437 614 1442
rect 2201 1437 2206 1442
rect 369 1432 518 1437
rect 609 1432 1022 1437
rect 2177 1432 2206 1437
rect 2265 1437 2270 1442
rect 2265 1432 2294 1437
rect 137 1422 182 1427
rect 201 1422 278 1427
rect 369 1417 374 1432
rect 529 1422 582 1427
rect 0 1412 126 1417
rect 289 1412 374 1417
rect 393 1412 478 1417
rect 121 1407 294 1412
rect 593 1402 598 1427
rect 713 1422 758 1427
rect 1073 1422 1246 1427
rect 1473 1422 1582 1427
rect 1721 1422 1814 1427
rect 2217 1422 2286 1427
rect 2537 1422 2598 1427
rect 2897 1422 2950 1427
rect 689 1412 894 1417
rect 1177 1412 1278 1417
rect 2049 1412 2238 1417
rect 2569 1412 2926 1417
rect 689 1397 694 1412
rect 777 1402 1158 1407
rect 2785 1402 2878 1407
rect 0 1392 694 1397
rect 705 1392 758 1397
rect 769 1392 830 1397
rect 825 1387 830 1392
rect 945 1392 998 1397
rect 945 1387 950 1392
rect 553 1382 598 1387
rect 825 1382 950 1387
rect 993 1387 998 1392
rect 1121 1392 1150 1397
rect 1265 1392 1334 1397
rect 1609 1392 1702 1397
rect 1857 1392 1950 1397
rect 1121 1387 1126 1392
rect 2841 1387 2926 1392
rect 993 1382 1126 1387
rect 2609 1382 2766 1387
rect 2817 1382 2846 1387
rect 2921 1382 3088 1387
rect 785 1372 806 1377
rect 2433 1372 2534 1377
rect 2609 1367 2614 1382
rect 2761 1377 2766 1382
rect 2761 1372 2910 1377
rect 0 1362 670 1367
rect 753 1362 1406 1367
rect 2017 1362 2614 1367
rect 2633 1362 2662 1367
rect 2921 1362 3088 1367
rect 1009 1352 1038 1357
rect 1569 1352 1742 1357
rect 1569 1347 1574 1352
rect 0 1342 118 1347
rect 145 1342 206 1347
rect 217 1342 286 1347
rect 753 1342 870 1347
rect 881 1342 958 1347
rect 1137 1342 1574 1347
rect 1737 1347 1742 1352
rect 1737 1342 1974 1347
rect 2017 1342 2022 1362
rect 2657 1357 2662 1362
rect 2785 1357 2926 1362
rect 2657 1352 2790 1357
rect 2089 1342 2198 1347
rect 2497 1342 2542 1347
rect 2809 1342 2910 1347
rect 753 1337 758 1342
rect 977 1337 1102 1342
rect 2905 1337 2910 1342
rect 305 1332 446 1337
rect 305 1327 310 1332
rect 0 1322 310 1327
rect 441 1327 446 1332
rect 489 1332 758 1337
rect 865 1332 982 1337
rect 1097 1332 1126 1337
rect 489 1327 494 1332
rect 1121 1327 1126 1332
rect 1441 1332 1470 1337
rect 1657 1332 1726 1337
rect 2489 1332 2534 1337
rect 2905 1332 3014 1337
rect 1441 1327 1446 1332
rect 2529 1327 2534 1332
rect 2993 1327 2998 1332
rect 441 1322 494 1327
rect 993 1322 1078 1327
rect 1121 1322 1446 1327
rect 1585 1317 1590 1327
rect 1617 1322 1718 1327
rect 2353 1322 2446 1327
rect 2529 1322 2622 1327
rect 2761 1322 2886 1327
rect 2993 1322 3088 1327
rect 937 1312 1102 1317
rect 1465 1312 1590 1317
rect 1961 1312 2206 1317
rect 2257 1312 2366 1317
rect 2513 1312 2542 1317
rect 0 1302 758 1307
rect 793 1302 1030 1307
rect 1025 1297 1030 1302
rect 1113 1302 1406 1307
rect 2113 1302 2190 1307
rect 2737 1302 2766 1307
rect 1113 1297 1118 1302
rect 2761 1297 2766 1302
rect 2849 1302 2878 1307
rect 2849 1297 2854 1302
rect 1025 1292 1118 1297
rect 1521 1292 2022 1297
rect 2761 1292 2854 1297
rect 0 1282 910 1287
rect 985 1262 1150 1267
rect 1657 1262 2110 1267
rect 985 1257 990 1262
rect 0 1252 726 1257
rect 961 1252 990 1257
rect 1145 1257 1150 1262
rect 1145 1252 1174 1257
rect 1921 1252 1950 1257
rect 1945 1247 1950 1252
rect 2089 1252 2174 1257
rect 2089 1247 2094 1252
rect 1009 1242 1126 1247
rect 913 1237 1014 1242
rect 1121 1237 1126 1242
rect 1217 1242 1318 1247
rect 1497 1242 1734 1247
rect 1945 1242 2094 1247
rect 1217 1237 1222 1242
rect 0 1232 206 1237
rect 689 1232 806 1237
rect 889 1232 918 1237
rect 1121 1232 1222 1237
rect 1313 1237 1318 1242
rect 1313 1232 1526 1237
rect 1585 1232 1694 1237
rect 2113 1232 2230 1237
rect 2241 1232 2318 1237
rect 2833 1232 2982 1237
rect 689 1227 694 1232
rect 665 1222 694 1227
rect 801 1227 806 1232
rect 2241 1227 2246 1232
rect 801 1222 958 1227
rect 1025 1222 1110 1227
rect 1145 1222 1270 1227
rect 1441 1222 1558 1227
rect 1673 1222 1702 1227
rect 2209 1222 2246 1227
rect 2321 1222 2382 1227
rect 2729 1222 2774 1227
rect 953 1217 1030 1222
rect 1553 1217 1678 1222
rect 97 1212 246 1217
rect 377 1212 526 1217
rect 617 1212 702 1217
rect 745 1212 790 1217
rect 1073 1212 1302 1217
rect 1785 1212 1862 1217
rect 2081 1207 2086 1217
rect 2865 1212 2894 1217
rect 881 1202 1294 1207
rect 1313 1202 1398 1207
rect 1505 1202 1806 1207
rect 2081 1202 2118 1207
rect 2713 1202 2798 1207
rect 153 1192 270 1197
rect 769 1192 902 1197
rect 1089 1192 1254 1197
rect 1337 1192 1494 1197
rect 1809 1192 1838 1197
rect 2009 1192 2246 1197
rect 2785 1192 2854 1197
rect 1489 1187 1590 1192
rect 1809 1187 1814 1192
rect 2865 1187 2870 1212
rect 2889 1207 2894 1212
rect 2993 1212 3088 1217
rect 2993 1207 2998 1212
rect 2889 1202 2998 1207
rect 241 1182 494 1187
rect 1129 1182 1182 1187
rect 1585 1182 1814 1187
rect 2257 1182 2326 1187
rect 2761 1182 2870 1187
rect 1953 1177 2070 1182
rect 921 1172 1070 1177
rect 1225 1172 1382 1177
rect 1425 1172 1566 1177
rect 1929 1172 1958 1177
rect 2065 1172 2126 1177
rect 921 1167 926 1172
rect 241 1162 334 1167
rect 705 1162 926 1167
rect 1065 1167 1070 1172
rect 1425 1167 1430 1172
rect 1065 1162 1174 1167
rect 1401 1162 1430 1167
rect 1561 1167 1566 1172
rect 2121 1167 2126 1172
rect 2257 1172 2286 1177
rect 2569 1172 2622 1177
rect 2257 1167 2262 1172
rect 1561 1162 2054 1167
rect 2121 1162 2262 1167
rect 2817 1162 2950 1167
rect 1257 1157 1350 1162
rect 385 1152 446 1157
rect 513 1152 686 1157
rect 1233 1152 1262 1157
rect 1345 1152 1550 1157
rect 2601 1152 2702 1157
rect 513 1137 518 1152
rect 489 1132 518 1137
rect 681 1137 686 1152
rect 769 1142 838 1147
rect 913 1142 1334 1147
rect 1913 1142 2102 1147
rect 2337 1137 2342 1147
rect 2745 1142 2886 1147
rect 681 1132 742 1137
rect 1281 1132 1414 1137
rect 1497 1132 1726 1137
rect 2161 1132 2342 1137
rect 2441 1132 2526 1137
rect 1113 1127 1222 1132
rect 2441 1127 2446 1132
rect 217 1122 558 1127
rect 641 1122 750 1127
rect 1025 1122 1118 1127
rect 1217 1122 1270 1127
rect 1425 1122 1486 1127
rect 1577 1122 1606 1127
rect 2049 1122 2110 1127
rect 2417 1122 2446 1127
rect 2521 1127 2526 1132
rect 2521 1122 2550 1127
rect 2737 1122 2878 1127
rect 2897 1122 3088 1127
rect 1265 1117 1430 1122
rect 1481 1117 1582 1122
rect 2049 1117 2054 1122
rect 2897 1117 2902 1122
rect 145 1112 230 1117
rect 497 1112 582 1117
rect 593 1112 622 1117
rect 761 1112 886 1117
rect 953 1112 1022 1117
rect 1153 1112 1206 1117
rect 1985 1112 2054 1117
rect 2081 1112 2182 1117
rect 2345 1112 2398 1117
rect 2425 1112 2534 1117
rect 2809 1112 2902 1117
rect 617 1107 766 1112
rect 1321 1102 1350 1107
rect 1345 1097 1350 1102
rect 1409 1102 1438 1107
rect 1481 1102 1534 1107
rect 2145 1102 2198 1107
rect 1409 1097 1414 1102
rect 113 1092 142 1097
rect 137 1087 142 1092
rect 241 1092 614 1097
rect 241 1087 246 1092
rect 137 1082 246 1087
rect 609 1087 614 1092
rect 713 1092 910 1097
rect 1105 1092 1246 1097
rect 1345 1092 1414 1097
rect 2337 1092 2446 1097
rect 713 1087 718 1092
rect 609 1082 718 1087
rect 1041 1082 1102 1087
rect 2113 1082 2174 1087
rect 2081 1072 2190 1077
rect 481 1062 590 1067
rect 481 1057 486 1062
rect 457 1052 486 1057
rect 585 1057 590 1062
rect 737 1062 830 1067
rect 737 1057 742 1062
rect 585 1052 742 1057
rect 825 1057 830 1062
rect 873 1062 1294 1067
rect 1417 1062 1486 1067
rect 1721 1062 1910 1067
rect 2713 1062 2750 1067
rect 873 1057 878 1062
rect 825 1052 878 1057
rect 1289 1057 1294 1062
rect 1289 1052 1318 1057
rect 769 1042 878 1047
rect 993 1042 1166 1047
rect 1625 1042 1678 1047
rect 2713 1042 2790 1047
rect 265 1032 294 1037
rect 313 1032 438 1037
rect 481 1032 574 1037
rect 753 1032 798 1037
rect 809 1032 982 1037
rect 1177 1032 1334 1037
rect 1425 1032 1558 1037
rect 2521 1032 2566 1037
rect 2753 1032 2886 1037
rect 313 1027 318 1032
rect 161 1022 318 1027
rect 433 1027 438 1032
rect 977 1027 1070 1032
rect 1177 1027 1182 1032
rect 1425 1027 1430 1032
rect 433 1022 518 1027
rect 513 1017 518 1022
rect 585 1022 646 1027
rect 1065 1022 1182 1027
rect 1305 1022 1430 1027
rect 1553 1027 1558 1032
rect 1553 1022 1582 1027
rect 1721 1022 1854 1027
rect 1921 1022 2078 1027
rect 2265 1022 2326 1027
rect 2449 1022 2542 1027
rect 2681 1022 2734 1027
rect 585 1017 590 1022
rect 513 1012 590 1017
rect 761 1012 1046 1017
rect 1489 1007 1494 1017
rect 1785 1012 1862 1017
rect 1921 1007 1926 1022
rect 169 1002 494 1007
rect 1065 1002 1246 1007
rect 929 997 1070 1002
rect 1241 997 1246 1002
rect 1441 1002 1494 1007
rect 1521 1002 1622 1007
rect 1889 1002 1926 1007
rect 2073 1007 2078 1022
rect 2793 1012 3088 1017
rect 2073 1002 2206 1007
rect 1441 997 1446 1002
rect 561 992 814 997
rect 905 992 934 997
rect 1241 992 1446 997
rect 1465 992 1678 997
rect 1937 992 2062 997
rect 2505 992 2606 997
rect 2721 992 2774 997
rect 561 987 566 992
rect 193 982 374 987
rect 369 977 374 982
rect 505 982 566 987
rect 689 982 1230 987
rect 2449 982 2526 987
rect 2793 982 3062 987
rect 505 977 510 982
rect 1625 977 1694 982
rect 2641 977 2718 982
rect 2793 977 2798 982
rect 369 972 510 977
rect 609 972 910 977
rect 1081 972 1126 977
rect 1553 972 1630 977
rect 1689 972 1718 977
rect 1945 972 2046 977
rect 2081 972 2150 977
rect 2617 972 2646 977
rect 2713 972 2798 977
rect 3057 977 3062 982
rect 3057 972 3088 977
rect 2081 967 2086 972
rect 201 962 350 967
rect 577 962 694 967
rect 721 957 726 967
rect 953 962 1054 967
rect 1241 962 1342 967
rect 1361 962 1526 967
rect 1641 962 1670 967
rect 953 957 958 962
rect 105 952 182 957
rect 721 952 958 957
rect 1049 957 1054 962
rect 1361 957 1366 962
rect 1049 952 1366 957
rect 1521 957 1526 962
rect 1665 957 1670 962
rect 1729 962 1862 967
rect 1953 962 2086 967
rect 2145 967 2150 972
rect 2145 962 2230 967
rect 2497 962 2702 967
rect 1729 957 1734 962
rect 1521 952 1598 957
rect 1665 952 1734 957
rect 2697 957 2702 962
rect 2809 962 2934 967
rect 2809 957 2814 962
rect 2697 952 2814 957
rect 2937 952 3088 957
rect 105 947 110 952
rect 81 942 110 947
rect 177 947 182 952
rect 177 942 278 947
rect 273 937 278 942
rect 345 942 470 947
rect 497 942 710 947
rect 345 937 350 942
rect 705 937 710 942
rect 785 942 814 947
rect 969 942 1038 947
rect 1169 942 1278 947
rect 785 937 790 942
rect 1273 937 1278 942
rect 1377 942 1430 947
rect 2041 942 2134 947
rect 2441 942 2486 947
rect 1377 937 1382 942
rect 2481 937 2486 942
rect 2553 942 2606 947
rect 2553 937 2558 942
rect 121 932 174 937
rect 273 932 350 937
rect 369 932 406 937
rect 113 922 206 927
rect 641 917 646 937
rect 705 932 790 937
rect 841 932 1022 937
rect 1185 932 1214 937
rect 1273 932 1382 937
rect 1417 932 1510 937
rect 2481 932 2558 937
rect 2601 937 2606 942
rect 2841 942 2926 947
rect 2841 937 2846 942
rect 2601 932 2846 937
rect 2921 937 2926 942
rect 2921 932 2998 937
rect 1057 922 1150 927
rect 865 917 1062 922
rect 1145 917 1150 922
rect 1185 917 1190 932
rect 2993 927 2998 932
rect 1201 922 1254 927
rect 2993 922 3088 927
rect 393 912 502 917
rect 641 912 870 917
rect 1145 912 1230 917
rect 1257 912 1326 917
rect 1577 912 1710 917
rect 2113 912 2406 917
rect 2865 912 2982 917
rect 881 902 1294 907
rect 1433 902 1638 907
rect 2025 902 2126 907
rect 2457 902 2638 907
rect 3057 902 3088 907
rect 1313 897 1414 902
rect 3057 897 3062 902
rect 833 892 862 897
rect 1017 892 1318 897
rect 1409 892 1478 897
rect 2729 892 3062 897
rect 857 887 1022 892
rect 1569 887 1678 892
rect 1041 882 1574 887
rect 1673 882 1702 887
rect 2385 882 2446 887
rect 2441 877 2446 882
rect 2561 882 2590 887
rect 2561 877 2566 882
rect 225 872 1030 877
rect 1025 867 1030 872
rect 1121 872 1182 877
rect 1225 872 1254 877
rect 1585 872 1662 877
rect 2441 872 2566 877
rect 1121 867 1126 872
rect 1249 867 1414 872
rect 1025 862 1126 867
rect 1409 857 1414 867
rect 1585 857 1590 872
rect 1609 862 1638 867
rect 793 852 870 857
rect 865 847 870 852
rect 1145 852 1390 857
rect 1409 852 1590 857
rect 1633 857 1638 862
rect 1713 862 1966 867
rect 2817 862 2886 867
rect 1713 857 1718 862
rect 2817 857 2822 862
rect 1633 852 1718 857
rect 2793 852 2822 857
rect 2881 857 2886 862
rect 2881 852 2910 857
rect 1145 847 1150 852
rect 489 842 582 847
rect 865 842 1150 847
rect 489 837 494 842
rect 385 832 494 837
rect 577 837 582 842
rect 577 832 622 837
rect 817 832 846 837
rect 1281 832 1358 837
rect 2073 832 2134 837
rect 2689 832 2830 837
rect 2865 832 2998 837
rect 129 822 222 827
rect 1169 822 1654 827
rect 2633 822 2726 827
rect 1169 817 1174 822
rect 2721 817 2726 822
rect 465 812 566 817
rect 761 812 846 817
rect 1033 812 1174 817
rect 1185 812 1406 817
rect 2113 812 2494 817
rect 2721 812 3088 817
rect 193 807 302 812
rect 1425 807 1534 812
rect 169 802 198 807
rect 297 802 518 807
rect 1089 802 1430 807
rect 1529 802 1718 807
rect 193 792 286 797
rect 497 792 678 797
rect 737 792 798 797
rect 1009 792 1518 797
rect 2537 792 2742 797
rect 2737 787 2742 792
rect 2865 792 2894 797
rect 2865 787 2870 792
rect 1121 782 1150 787
rect 1321 782 1494 787
rect 2737 782 2870 787
rect 2929 782 3088 787
rect 1145 777 1326 782
rect 313 772 446 777
rect 569 772 630 777
rect 825 772 982 777
rect 1345 772 1478 777
rect 825 767 830 772
rect 801 762 830 767
rect 977 767 982 772
rect 977 762 1334 767
rect 1329 757 1334 762
rect 1577 762 1766 767
rect 1577 757 1582 762
rect 825 752 886 757
rect 1329 752 1422 757
rect 1441 752 1582 757
rect 1761 757 1766 762
rect 1761 752 1790 757
rect 2817 752 2886 757
rect 1441 747 1446 752
rect 337 742 742 747
rect 889 742 966 747
rect 1081 742 1158 747
rect 1177 742 1318 747
rect 225 732 358 737
rect 409 732 438 737
rect 433 727 438 732
rect 553 732 582 737
rect 553 727 558 732
rect 433 722 558 727
rect 1153 717 1158 742
rect 1313 737 1318 742
rect 1377 742 1446 747
rect 2593 742 2742 747
rect 1377 737 1382 742
rect 2593 737 2598 742
rect 1313 732 1382 737
rect 1401 732 1830 737
rect 2209 732 2598 737
rect 1401 717 1406 732
rect 1913 722 1950 727
rect 2993 722 3088 727
rect 1153 712 1406 717
rect 1641 712 1710 717
rect 1817 712 1966 717
rect 441 702 822 707
rect 2297 692 2454 697
rect 2505 682 2558 687
rect 945 672 1030 677
rect 945 667 950 672
rect 921 662 950 667
rect 1025 667 1030 672
rect 1073 672 1230 677
rect 1073 667 1078 672
rect 1025 662 1078 667
rect 1225 667 1230 672
rect 1361 672 1478 677
rect 1361 667 1366 672
rect 1225 662 1366 667
rect 1473 667 1478 672
rect 1473 662 1566 667
rect 2769 662 3006 667
rect 625 652 694 657
rect 625 647 630 652
rect 601 642 630 647
rect 689 647 694 652
rect 2585 652 2662 657
rect 2585 647 2590 652
rect 689 642 1214 647
rect 1209 637 1214 642
rect 1297 642 1462 647
rect 2097 642 2182 647
rect 2561 642 2590 647
rect 2657 647 2662 652
rect 2769 647 2774 662
rect 3001 657 3006 662
rect 3001 652 3088 657
rect 2657 642 2774 647
rect 2785 642 2870 647
rect 1297 637 1302 642
rect 2097 637 2102 642
rect 265 632 350 637
rect 577 632 678 637
rect 905 632 982 637
rect 1209 632 1302 637
rect 1593 632 1686 637
rect 2073 632 2102 637
rect 2177 637 2182 642
rect 2177 632 2206 637
rect 2433 632 2686 637
rect 2681 627 2686 632
rect 2785 632 2990 637
rect 2785 627 2790 632
rect 2985 627 2990 632
rect 3057 632 3088 637
rect 3057 627 3062 632
rect 201 622 678 627
rect 969 622 1086 627
rect 1113 622 1190 627
rect 1417 622 1470 627
rect 2241 622 2406 627
rect 2681 622 2790 627
rect 2849 622 2934 627
rect 2985 622 3062 627
rect 321 612 358 617
rect 529 612 622 617
rect 673 607 678 622
rect 2241 617 2246 622
rect 697 612 886 617
rect 1321 612 1390 617
rect 1561 612 1622 617
rect 1649 612 1950 617
rect 2057 612 2246 617
rect 2577 612 2662 617
rect 697 607 702 612
rect 137 602 222 607
rect 673 602 702 607
rect 881 607 886 612
rect 881 602 1174 607
rect 2225 602 2230 612
rect 2681 602 2782 607
rect 1169 597 1174 602
rect 2681 597 2686 602
rect 321 592 350 597
rect 513 592 598 597
rect 609 592 750 597
rect 1169 592 1198 597
rect 1841 592 1902 597
rect 2569 592 2686 597
rect 2777 597 2782 602
rect 2777 592 2806 597
rect 593 587 598 592
rect 201 582 278 587
rect 465 582 550 587
rect 593 582 1014 587
rect 1009 577 1014 582
rect 1137 582 1166 587
rect 1697 582 1822 587
rect 1137 577 1142 582
rect 1697 577 1702 582
rect 89 572 190 577
rect 185 567 190 572
rect 273 572 422 577
rect 1009 572 1142 577
rect 1473 572 1702 577
rect 1817 577 1822 582
rect 1921 582 1974 587
rect 1921 577 1926 582
rect 2697 577 2878 582
rect 1817 572 1926 577
rect 2305 572 2374 577
rect 273 567 278 572
rect 2305 567 2310 572
rect 185 562 278 567
rect 297 562 326 567
rect 409 562 462 567
rect 657 562 734 567
rect 1417 562 1446 567
rect 1529 562 1558 567
rect 1649 562 1878 567
rect 1977 562 2310 567
rect 2369 567 2374 572
rect 2481 572 2702 577
rect 2873 572 3006 577
rect 2481 567 2486 572
rect 2369 562 2486 567
rect 2713 562 2758 567
rect 2777 562 2862 567
rect 321 557 414 562
rect 1441 557 1534 562
rect 481 552 630 557
rect 785 552 926 557
rect 1297 552 1398 557
rect 2321 552 2462 557
rect 2481 552 2622 557
rect 481 547 486 552
rect 225 542 326 547
rect 449 542 486 547
rect 625 547 630 552
rect 1297 547 1302 552
rect 625 542 654 547
rect 721 542 830 547
rect 721 537 726 542
rect 825 537 830 542
rect 905 542 1030 547
rect 1201 542 1302 547
rect 1393 547 1398 552
rect 1393 542 1462 547
rect 1697 542 1798 547
rect 905 537 910 542
rect 1201 537 1206 542
rect 1697 537 1702 542
rect 641 532 726 537
rect 737 532 806 537
rect 825 532 910 537
rect 1017 532 1206 537
rect 1313 532 1702 537
rect 1793 537 1798 542
rect 1881 542 1910 547
rect 1881 537 1886 542
rect 1793 532 1886 537
rect 2681 532 2750 537
rect 2681 527 2686 532
rect 345 522 630 527
rect 1697 522 1774 527
rect 2433 522 2686 527
rect 2745 527 2750 532
rect 2745 522 2774 527
rect 777 512 870 517
rect 1001 512 1094 517
rect 1201 512 1326 517
rect 2025 512 2198 517
rect 2481 512 2486 522
rect 2697 512 2734 517
rect 2817 512 2950 517
rect 505 502 574 507
rect 1929 502 2022 507
rect 2073 502 2110 507
rect 505 497 510 502
rect 249 492 510 497
rect 569 497 574 502
rect 1065 497 1142 502
rect 569 492 598 497
rect 833 492 1070 497
rect 1137 492 1270 497
rect 833 487 838 492
rect 1265 487 1270 492
rect 1337 492 1478 497
rect 1337 487 1342 492
rect 209 482 238 487
rect 233 477 238 482
rect 337 482 550 487
rect 337 477 342 482
rect 233 472 342 477
rect 545 477 550 482
rect 609 482 838 487
rect 857 482 886 487
rect 609 477 614 482
rect 545 472 614 477
rect 881 477 886 482
rect 993 482 1126 487
rect 993 477 998 482
rect 881 472 998 477
rect 1121 477 1126 482
rect 1217 482 1246 487
rect 1265 482 1342 487
rect 2769 482 3088 487
rect 1217 477 1222 482
rect 1121 472 1222 477
rect 1921 472 2134 477
rect 465 452 710 457
rect 513 432 622 437
rect 2153 432 2318 437
rect 1161 422 1238 427
rect 1161 417 1166 422
rect 1137 412 1166 417
rect 1233 417 1238 422
rect 1537 422 1710 427
rect 2529 422 2582 427
rect 2633 422 2726 427
rect 2753 422 2830 427
rect 1233 412 1262 417
rect 1537 407 1542 422
rect 177 402 542 407
rect 1185 402 1294 407
rect 1513 402 1542 407
rect 1705 407 1710 422
rect 1777 412 1918 417
rect 2145 412 2222 417
rect 2145 407 2150 412
rect 1705 402 1734 407
rect 2121 402 2150 407
rect 2217 407 2222 412
rect 2217 402 2406 407
rect 801 392 934 397
rect 1033 392 1150 397
rect 1385 392 1486 397
rect 1505 392 1694 397
rect 457 382 558 387
rect 761 382 814 387
rect 1041 382 1070 387
rect 1065 377 1070 382
rect 1153 382 1414 387
rect 1153 377 1158 382
rect 1065 372 1158 377
rect 1409 377 1414 382
rect 1505 377 1510 392
rect 1689 387 1694 392
rect 1825 392 1854 397
rect 2105 392 2206 397
rect 1825 387 1830 392
rect 1689 382 1830 387
rect 2465 382 2574 387
rect 2465 377 2470 382
rect 1409 372 1510 377
rect 2393 372 2470 377
rect 2569 377 2574 382
rect 2569 372 2838 377
rect 2313 362 2406 367
rect 177 352 358 357
rect 705 352 790 357
rect 1177 352 1390 357
rect 1569 352 1662 357
rect 2153 352 2238 357
rect 2257 352 2566 357
rect 705 347 710 352
rect 89 342 246 347
rect 473 342 662 347
rect 681 342 710 347
rect 785 347 790 352
rect 2153 347 2158 352
rect 785 342 814 347
rect 921 342 966 347
rect 1505 342 1558 347
rect 473 327 478 342
rect 0 322 270 327
rect 449 322 478 327
rect 657 327 662 342
rect 1553 337 1558 342
rect 1641 342 1670 347
rect 2049 342 2158 347
rect 2233 347 2238 352
rect 2233 342 2254 347
rect 1641 337 1646 342
rect 2249 337 2254 342
rect 2385 342 2414 347
rect 2385 337 2390 342
rect 985 332 1110 337
rect 1553 332 1646 337
rect 2065 332 2102 337
rect 985 327 990 332
rect 657 322 694 327
rect 721 322 990 327
rect 1105 327 1110 332
rect 2097 327 2102 332
rect 2169 332 2222 337
rect 2249 332 2390 337
rect 2753 332 2966 337
rect 2169 327 2174 332
rect 1105 322 1134 327
rect 1849 322 1942 327
rect 1977 322 2078 327
rect 2097 322 2174 327
rect 233 312 302 317
rect 433 312 662 317
rect 1601 312 1718 317
rect 2209 312 2262 317
rect 2329 312 2510 317
rect 2553 312 2614 317
rect 2817 312 2846 317
rect 2841 307 2846 312
rect 2945 312 2974 317
rect 2945 307 2950 312
rect 593 302 1342 307
rect 1433 302 1542 307
rect 1777 302 1870 307
rect 2065 302 2134 307
rect 2289 302 2358 307
rect 2841 302 2950 307
rect 801 272 1166 277
rect 2081 262 2166 267
rect 2225 262 2462 267
rect 1121 252 1526 257
rect 2225 247 2230 262
rect 545 242 622 247
rect 753 242 862 247
rect 881 242 926 247
rect 1681 242 1782 247
rect 753 237 758 242
rect 497 232 758 237
rect 857 237 862 242
rect 1681 237 1686 242
rect 857 232 878 237
rect 873 227 878 232
rect 937 232 1198 237
rect 1545 232 1638 237
rect 1657 232 1686 237
rect 1777 237 1782 242
rect 1825 242 1910 247
rect 1929 242 2022 247
rect 2201 242 2230 247
rect 2457 247 2462 262
rect 2457 242 2622 247
rect 2689 242 2774 247
rect 1825 237 1830 242
rect 1777 232 1830 237
rect 1905 237 1910 242
rect 2689 237 2694 242
rect 1905 232 2446 237
rect 2633 232 2694 237
rect 2769 237 2774 242
rect 2769 232 2798 237
rect 937 227 942 232
rect 1545 227 1550 232
rect 873 222 942 227
rect 1441 222 1550 227
rect 1633 227 1638 232
rect 2441 227 2518 232
rect 2633 227 2638 232
rect 1633 222 1878 227
rect 2513 222 2638 227
rect 2897 222 2974 227
rect 1873 217 1878 222
rect 769 212 846 217
rect 1297 212 1430 217
rect 1425 207 1430 212
rect 1529 212 1622 217
rect 1529 207 1534 212
rect 97 202 174 207
rect 561 202 678 207
rect 905 202 1270 207
rect 1425 202 1534 207
rect 1617 207 1622 212
rect 1753 212 1782 217
rect 1873 212 2286 217
rect 2321 212 2374 217
rect 1753 207 1758 212
rect 2369 207 2374 212
rect 2465 212 2494 217
rect 2705 212 2814 217
rect 2465 207 2470 212
rect 1617 202 1646 207
rect 1729 202 1758 207
rect 2249 202 2350 207
rect 2369 202 2470 207
rect 561 197 566 202
rect 377 192 462 197
rect 537 192 566 197
rect 673 197 678 202
rect 1641 197 1734 202
rect 673 192 966 197
rect 1561 192 1590 197
rect 1585 187 1590 192
rect 1785 192 1862 197
rect 1785 187 1790 192
rect 385 182 518 187
rect 1009 182 1142 187
rect 1585 182 1790 187
rect 1857 187 1862 192
rect 1937 192 2022 197
rect 1937 187 1942 192
rect 1857 182 1942 187
rect 2113 182 2166 187
rect 1009 177 1014 182
rect 433 172 462 177
rect 457 167 462 172
rect 529 172 1014 177
rect 1449 172 1534 177
rect 529 167 534 172
rect 1449 167 1454 172
rect 457 162 534 167
rect 1425 162 1454 167
rect 1529 167 1534 172
rect 2721 172 2854 177
rect 2721 167 2726 172
rect 1529 162 1558 167
rect 2697 162 2726 167
rect 2849 167 2854 172
rect 2849 162 2878 167
rect 337 152 414 157
rect 625 152 718 157
rect 753 152 910 157
rect 1585 152 1694 157
rect 2073 152 2182 157
rect 2609 152 2902 157
rect 337 147 342 152
rect 89 142 342 147
rect 409 147 414 152
rect 1585 147 1590 152
rect 409 142 606 147
rect 905 142 942 147
rect 1057 142 1166 147
rect 1417 142 1502 147
rect 1561 142 1590 147
rect 1689 147 1694 152
rect 1689 142 2062 147
rect 2193 142 2542 147
rect 601 137 774 142
rect 905 137 910 142
rect 2057 137 2198 142
rect 769 132 910 137
rect 1185 132 1254 137
rect 1321 132 1510 137
rect 1057 127 1134 132
rect 1185 127 1190 132
rect 353 122 422 127
rect 681 122 750 127
rect 929 122 1062 127
rect 1129 122 1190 127
rect 1249 127 1254 132
rect 1697 127 1702 137
rect 1249 122 1342 127
rect 1337 117 1342 122
rect 1449 122 1686 127
rect 1697 122 1718 127
rect 2137 122 2190 127
rect 1449 117 1454 122
rect 273 112 374 117
rect 1073 112 1118 117
rect 1113 107 1118 112
rect 1193 112 1246 117
rect 1337 112 1454 117
rect 1473 112 1566 117
rect 1689 112 1742 117
rect 1961 112 2110 117
rect 2553 112 2630 117
rect 2689 112 2766 117
rect 1193 107 1198 112
rect 377 102 670 107
rect 665 97 670 102
rect 761 102 886 107
rect 1113 102 1198 107
rect 1241 107 1246 112
rect 1241 102 1318 107
rect 761 97 766 102
rect 1313 97 1318 102
rect 1537 102 1566 107
rect 2145 102 2278 107
rect 1537 97 1542 102
rect 665 92 766 97
rect 993 92 1094 97
rect 1313 92 1542 97
rect 2625 87 2630 112
rect 2745 102 2878 107
rect 2793 87 2902 92
rect 2625 82 2798 87
rect 2897 82 2990 87
rect 2617 72 2646 77
rect 2641 67 2646 72
rect 2761 72 2862 77
rect 2761 67 2766 72
rect 873 62 1334 67
rect 1569 62 1598 67
rect 2641 62 2766 67
rect 2857 67 2862 72
rect 2929 72 2958 77
rect 2929 67 2934 72
rect 2857 62 2934 67
rect 2545 42 2758 47
use AND2X2  AND2X2_0
timestamp 1713400504
transform 1 0 744 0 1 2570
box -8 -3 40 105
use AND2X2  AND2X2_1
timestamp 1713400504
transform 1 0 640 0 -1 2570
box -8 -3 40 105
use AND2X2  AND2X2_2
timestamp 1713400504
transform 1 0 504 0 -1 2570
box -8 -3 40 105
use AND2X2  AND2X2_3
timestamp 1713400504
transform 1 0 272 0 1 1970
box -8 -3 40 105
use AND2X2  AND2X2_4
timestamp 1713400504
transform 1 0 1352 0 -1 1770
box -8 -3 40 105
use AND2X2  AND2X2_5
timestamp 1713400504
transform 1 0 1304 0 1 1370
box -8 -3 40 105
use AND2X2  AND2X2_6
timestamp 1713400504
transform 1 0 1936 0 1 770
box -8 -3 40 105
use AND2X2  AND2X2_7
timestamp 1713400504
transform 1 0 856 0 1 2570
box -8 -3 40 105
use AND2X2  AND2X2_8
timestamp 1713400504
transform 1 0 1312 0 1 170
box -8 -3 40 105
use AND2X2  AND2X2_9
timestamp 1713400504
transform 1 0 2296 0 -1 2370
box -8 -3 40 105
use AND2X2  AND2X2_10
timestamp 1713400504
transform 1 0 2320 0 1 770
box -8 -3 40 105
use AND2X2  AND2X2_11
timestamp 1713400504
transform 1 0 1664 0 1 970
box -8 -3 40 105
use AND2X2  AND2X2_12
timestamp 1713400504
transform 1 0 2080 0 -1 570
box -8 -3 40 105
use AND2X2  AND2X2_13
timestamp 1713400504
transform 1 0 2944 0 1 170
box -8 -3 40 105
use AND2X2  AND2X2_14
timestamp 1713400504
transform 1 0 2776 0 1 570
box -8 -3 40 105
use AOI21X1  AOI21X1_0
timestamp 1713400504
transform 1 0 1096 0 -1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_1
timestamp 1713400504
transform 1 0 248 0 1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_2
timestamp 1713400504
transform 1 0 224 0 -1 370
box -7 -3 39 105
use AOI21X1  AOI21X1_3
timestamp 1713400504
transform 1 0 2432 0 -1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_4
timestamp 1713400504
transform 1 0 2344 0 1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_5
timestamp 1713400504
transform 1 0 2592 0 -1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_6
timestamp 1713400504
transform 1 0 2520 0 1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_7
timestamp 1713400504
transform 1 0 2704 0 -1 2170
box -7 -3 39 105
use AOI21X1  AOI21X1_8
timestamp 1713400504
transform 1 0 1672 0 -1 2170
box -7 -3 39 105
use AOI21X1  AOI21X1_9
timestamp 1713400504
transform 1 0 2496 0 -1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_10
timestamp 1713400504
transform 1 0 1448 0 1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_11
timestamp 1713400504
transform 1 0 1648 0 1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_12
timestamp 1713400504
transform 1 0 1736 0 1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_13
timestamp 1713400504
transform 1 0 1752 0 -1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_14
timestamp 1713400504
transform 1 0 1160 0 -1 2170
box -7 -3 39 105
use AOI21X1  AOI21X1_15
timestamp 1713400504
transform 1 0 1216 0 -1 2370
box -7 -3 39 105
use AOI21X1  AOI21X1_16
timestamp 1713400504
transform 1 0 1360 0 1 570
box -7 -3 39 105
use AOI21X1  AOI21X1_17
timestamp 1713400504
transform 1 0 1440 0 1 370
box -7 -3 39 105
use AOI21X1  AOI21X1_18
timestamp 1713400504
transform 1 0 1152 0 -1 1570
box -7 -3 39 105
use AOI21X1  AOI21X1_19
timestamp 1713400504
transform 1 0 1224 0 1 1570
box -7 -3 39 105
use AOI21X1  AOI21X1_20
timestamp 1713400504
transform 1 0 1032 0 1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_21
timestamp 1713400504
transform 1 0 1120 0 1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_22
timestamp 1713400504
transform 1 0 2136 0 1 170
box -7 -3 39 105
use AOI21X1  AOI21X1_23
timestamp 1713400504
transform 1 0 2920 0 -1 570
box -7 -3 39 105
use AOI21X1  AOI21X1_24
timestamp 1713400504
transform 1 0 2952 0 1 570
box -7 -3 39 105
use AOI21X1  AOI21X1_25
timestamp 1713400504
transform 1 0 2904 0 1 370
box -7 -3 39 105
use AOI21X1  AOI21X1_26
timestamp 1713400504
transform 1 0 2704 0 -1 570
box -7 -3 39 105
use AOI21X1  AOI21X1_27
timestamp 1713400504
transform 1 0 2568 0 1 570
box -7 -3 39 105
use AOI21X1  AOI21X1_28
timestamp 1713400504
transform 1 0 2640 0 1 570
box -7 -3 39 105
use AOI21X1  AOI21X1_29
timestamp 1713400504
transform 1 0 2696 0 1 170
box -7 -3 39 105
use AOI22X1  AOI22X1_0
timestamp 1713400504
transform 1 0 2328 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_1
timestamp 1713400504
transform 1 0 2400 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_2
timestamp 1713400504
transform 1 0 2864 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_3
timestamp 1713400504
transform 1 0 2864 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_4
timestamp 1713400504
transform 1 0 2688 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_5
timestamp 1713400504
transform 1 0 2752 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_6
timestamp 1713400504
transform 1 0 2728 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_7
timestamp 1713400504
transform 1 0 2832 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_8
timestamp 1713400504
transform 1 0 2736 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_9
timestamp 1713400504
transform 1 0 2768 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_10
timestamp 1713400504
transform 1 0 1720 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_11
timestamp 1713400504
transform 1 0 1736 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_12
timestamp 1713400504
transform 1 0 2720 0 -1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_13
timestamp 1713400504
transform 1 0 2376 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_14
timestamp 1713400504
transform 1 0 1352 0 1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_15
timestamp 1713400504
transform 1 0 1408 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_16
timestamp 1713400504
transform 1 0 2480 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_17
timestamp 1713400504
transform 1 0 1920 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_18
timestamp 1713400504
transform 1 0 2528 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_19
timestamp 1713400504
transform 1 0 2608 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_20
timestamp 1713400504
transform 1 0 1832 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_21
timestamp 1713400504
transform 1 0 1744 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_22
timestamp 1713400504
transform 1 0 1088 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_23
timestamp 1713400504
transform 1 0 1672 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_24
timestamp 1713400504
transform 1 0 1448 0 1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_25
timestamp 1713400504
transform 1 0 1432 0 -1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_26
timestamp 1713400504
transform 1 0 1504 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_27
timestamp 1713400504
transform 1 0 1616 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_28
timestamp 1713400504
transform 1 0 2192 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_29
timestamp 1713400504
transform 1 0 2144 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_30
timestamp 1713400504
transform 1 0 1896 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_31
timestamp 1713400504
transform 1 0 1600 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_32
timestamp 1713400504
transform 1 0 1704 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_33
timestamp 1713400504
transform 1 0 1920 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_34
timestamp 1713400504
transform 1 0 1448 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_35
timestamp 1713400504
transform 1 0 1688 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_36
timestamp 1713400504
transform 1 0 1664 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_37
timestamp 1713400504
transform 1 0 1560 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_38
timestamp 1713400504
transform 1 0 1400 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_39
timestamp 1713400504
transform 1 0 1488 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_40
timestamp 1713400504
transform 1 0 1304 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_41
timestamp 1713400504
transform 1 0 1464 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_42
timestamp 1713400504
transform 1 0 1600 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_43
timestamp 1713400504
transform 1 0 1568 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_44
timestamp 1713400504
transform 1 0 1456 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_45
timestamp 1713400504
transform 1 0 1576 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_46
timestamp 1713400504
transform 1 0 1464 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_47
timestamp 1713400504
transform 1 0 1448 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_48
timestamp 1713400504
transform 1 0 1272 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_49
timestamp 1713400504
transform 1 0 1520 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_50
timestamp 1713400504
transform 1 0 1256 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_51
timestamp 1713400504
transform 1 0 1208 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_52
timestamp 1713400504
transform 1 0 2688 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_53
timestamp 1713400504
transform 1 0 2744 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_54
timestamp 1713400504
transform 1 0 2776 0 -1 370
box -8 -3 46 105
use BUFX2  BUFX2_0
timestamp 1713400504
transform 1 0 2688 0 1 1370
box -5 -3 28 105
use BUFX2  BUFX2_1
timestamp 1713400504
transform 1 0 2160 0 -1 1570
box -5 -3 28 105
use BUFX2  BUFX2_2
timestamp 1713400504
transform 1 0 728 0 1 1370
box -5 -3 28 105
use BUFX2  BUFX2_3
timestamp 1713400504
transform 1 0 2984 0 -1 770
box -5 -3 28 105
use BUFX2  BUFX2_4
timestamp 1713400504
transform 1 0 2512 0 -1 1370
box -5 -3 28 105
use BUFX2  BUFX2_5
timestamp 1713400504
transform 1 0 336 0 -1 370
box -5 -3 28 105
use BUFX2  BUFX2_6
timestamp 1713400504
transform 1 0 2192 0 1 2170
box -5 -3 28 105
use BUFX2  BUFX2_7
timestamp 1713400504
transform 1 0 2200 0 1 1770
box -5 -3 28 105
use BUFX2  BUFX2_8
timestamp 1713400504
transform 1 0 2160 0 1 2170
box -5 -3 28 105
use BUFX2  BUFX2_9
timestamp 1713400504
transform 1 0 704 0 1 1370
box -5 -3 28 105
use BUFX2  BUFX2_10
timestamp 1713400504
transform 1 0 608 0 1 1370
box -5 -3 28 105
use BUFX2  BUFX2_11
timestamp 1713400504
transform 1 0 584 0 1 1370
box -5 -3 28 105
use BUFX2  BUFX2_12
timestamp 1713400504
transform 1 0 2656 0 -1 1370
box -5 -3 28 105
use BUFX2  BUFX2_13
timestamp 1713400504
transform 1 0 2664 0 1 1370
box -5 -3 28 105
use BUFX2  BUFX2_14
timestamp 1713400504
transform 1 0 2168 0 1 1770
box -5 -3 28 105
use BUFX2  BUFX2_15
timestamp 1713400504
transform 1 0 2096 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_16
timestamp 1713400504
transform 1 0 2232 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_17
timestamp 1713400504
transform 1 0 2096 0 1 1570
box -5 -3 28 105
use BUFX2  BUFX2_18
timestamp 1713400504
transform 1 0 2440 0 -1 1970
box -5 -3 28 105
use BUFX2  BUFX2_19
timestamp 1713400504
transform 1 0 2128 0 1 1970
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_0
timestamp 1713400504
transform 1 0 1464 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_1
timestamp 1713400504
transform 1 0 80 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_2
timestamp 1713400504
transform 1 0 72 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_3
timestamp 1713400504
transform 1 0 584 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_4
timestamp 1713400504
transform 1 0 376 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_5
timestamp 1713400504
transform 1 0 80 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_6
timestamp 1713400504
transform 1 0 224 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_7
timestamp 1713400504
transform 1 0 408 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_8
timestamp 1713400504
transform 1 0 72 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_9
timestamp 1713400504
transform 1 0 80 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_10
timestamp 1713400504
transform 1 0 72 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_11
timestamp 1713400504
transform 1 0 240 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_12
timestamp 1713400504
transform 1 0 456 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_13
timestamp 1713400504
transform 1 0 400 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_14
timestamp 1713400504
transform 1 0 600 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_15
timestamp 1713400504
transform 1 0 928 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_16
timestamp 1713400504
transform 1 0 952 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_17
timestamp 1713400504
transform 1 0 616 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_18
timestamp 1713400504
transform 1 0 792 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_19
timestamp 1713400504
transform 1 0 568 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_20
timestamp 1713400504
transform 1 0 704 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_21
timestamp 1713400504
transform 1 0 464 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_22
timestamp 1713400504
transform 1 0 880 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_23
timestamp 1713400504
transform 1 0 496 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_24
timestamp 1713400504
transform 1 0 384 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_25
timestamp 1713400504
transform 1 0 128 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_26
timestamp 1713400504
transform 1 0 80 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_27
timestamp 1713400504
transform 1 0 424 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_28
timestamp 1713400504
transform 1 0 1024 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_29
timestamp 1713400504
transform 1 0 784 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_30
timestamp 1713400504
transform 1 0 1032 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_31
timestamp 1713400504
transform 1 0 1128 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_32
timestamp 1713400504
transform 1 0 1056 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_33
timestamp 1713400504
transform 1 0 832 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_34
timestamp 1713400504
transform 1 0 1704 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_35
timestamp 1713400504
transform 1 0 1864 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_36
timestamp 1713400504
transform 1 0 1840 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_37
timestamp 1713400504
transform 1 0 1568 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_38
timestamp 1713400504
transform 1 0 1640 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_39
timestamp 1713400504
transform 1 0 1696 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_40
timestamp 1713400504
transform 1 0 1976 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_41
timestamp 1713400504
transform 1 0 2072 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_42
timestamp 1713400504
transform 1 0 1704 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_43
timestamp 1713400504
transform 1 0 1800 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_44
timestamp 1713400504
transform 1 0 1696 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_45
timestamp 1713400504
transform 1 0 1504 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_46
timestamp 1713400504
transform 1 0 1456 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_47
timestamp 1713400504
transform 1 0 1552 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_48
timestamp 1713400504
transform 1 0 1432 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_49
timestamp 1713400504
transform 1 0 1536 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_50
timestamp 1713400504
transform 1 0 1984 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_51
timestamp 1713400504
transform 1 0 1984 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_52
timestamp 1713400504
transform 1 0 2216 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_53
timestamp 1713400504
transform 1 0 2312 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_54
timestamp 1713400504
transform 1 0 2400 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_55
timestamp 1713400504
transform 1 0 2200 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_56
timestamp 1713400504
transform 1 0 2712 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_57
timestamp 1713400504
transform 1 0 2720 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_58
timestamp 1713400504
transform 1 0 2752 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_59
timestamp 1713400504
transform 1 0 2448 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_60
timestamp 1713400504
transform 1 0 2400 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_61
timestamp 1713400504
transform 1 0 2544 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_62
timestamp 1713400504
transform 1 0 2768 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_63
timestamp 1713400504
transform 1 0 2768 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_64
timestamp 1713400504
transform 1 0 2200 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_65
timestamp 1713400504
transform 1 0 2152 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_66
timestamp 1713400504
transform 1 0 2208 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_67
timestamp 1713400504
transform 1 0 1600 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_68
timestamp 1713400504
transform 1 0 1360 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_69
timestamp 1713400504
transform 1 0 1608 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_70
timestamp 1713400504
transform 1 0 1288 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_71
timestamp 1713400504
transform 1 0 1160 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_72
timestamp 1713400504
transform 1 0 1056 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_73
timestamp 1713400504
transform 1 0 968 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_74
timestamp 1713400504
transform 1 0 1064 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_75
timestamp 1713400504
transform 1 0 1648 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_76
timestamp 1713400504
transform 1 0 1840 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_77
timestamp 1713400504
transform 1 0 2040 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_78
timestamp 1713400504
transform 1 0 2496 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_79
timestamp 1713400504
transform 1 0 2592 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_80
timestamp 1713400504
transform 1 0 2808 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_81
timestamp 1713400504
transform 1 0 2912 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_82
timestamp 1713400504
transform 1 0 2920 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_83
timestamp 1713400504
transform 1 0 2920 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_84
timestamp 1713400504
transform 1 0 2616 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_85
timestamp 1713400504
transform 1 0 2760 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_86
timestamp 1713400504
transform 1 0 2912 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_87
timestamp 1713400504
transform 1 0 2912 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_88
timestamp 1713400504
transform 1 0 2912 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_89
timestamp 1713400504
transform 1 0 2864 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_90
timestamp 1713400504
transform 1 0 2576 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_91
timestamp 1713400504
transform 1 0 2560 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_92
timestamp 1713400504
transform 1 0 2912 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_93
timestamp 1713400504
transform 1 0 2920 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_94
timestamp 1713400504
transform 1 0 2672 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_95
timestamp 1713400504
transform 1 0 2920 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_96
timestamp 1713400504
transform 1 0 2624 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_97
timestamp 1713400504
transform 1 0 2544 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_98
timestamp 1713400504
transform 1 0 2856 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_99
timestamp 1713400504
transform 1 0 2920 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_100
timestamp 1713400504
transform 1 0 2488 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_101
timestamp 1713400504
transform 1 0 2528 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_102
timestamp 1713400504
transform 1 0 2344 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_103
timestamp 1713400504
transform 1 0 2448 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_104
timestamp 1713400504
transform 1 0 2528 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_105
timestamp 1713400504
transform 1 0 2760 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_106
timestamp 1713400504
transform 1 0 2560 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_107
timestamp 1713400504
transform 1 0 2472 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_108
timestamp 1713400504
transform 1 0 2464 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_109
timestamp 1713400504
transform 1 0 2424 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_110
timestamp 1713400504
transform 1 0 2432 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_111
timestamp 1713400504
transform 1 0 2520 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_112
timestamp 1713400504
transform 1 0 1928 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_113
timestamp 1713400504
transform 1 0 1928 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_114
timestamp 1713400504
transform 1 0 2312 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_115
timestamp 1713400504
transform 1 0 1976 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_116
timestamp 1713400504
transform 1 0 2312 0 -1 170
box -8 -3 104 105
use FAX1  FAX1_0
timestamp 1713400504
transform 1 0 312 0 1 2370
box -5 -3 126 105
use FAX1  FAX1_1
timestamp 1713400504
transform 1 0 224 0 1 2170
box -5 -3 126 105
use FAX1  FAX1_2
timestamp 1713400504
transform 1 0 704 0 -1 2570
box -5 -3 126 105
use FAX1  FAX1_3
timestamp 1713400504
transform 1 0 680 0 1 2370
box -5 -3 126 105
use FAX1  FAX1_4
timestamp 1713400504
transform 1 0 528 0 1 2370
box -5 -3 126 105
use FAX1  FAX1_5
timestamp 1713400504
transform 1 0 512 0 -1 2370
box -5 -3 126 105
use FAX1  FAX1_6
timestamp 1713400504
transform 1 0 368 0 -1 2370
box -5 -3 126 105
use FAX1  FAX1_7
timestamp 1713400504
transform 1 0 704 0 -1 2170
box -5 -3 126 105
use FAX1  FAX1_8
timestamp 1713400504
transform 1 0 520 0 1 2170
box -5 -3 126 105
use FILL  FILL_0
timestamp 1713400504
transform 1 0 3008 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1
timestamp 1713400504
transform 1 0 3000 0 -1 2970
box -8 -3 16 105
use FILL  FILL_2
timestamp 1713400504
transform 1 0 2992 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3
timestamp 1713400504
transform 1 0 2984 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4
timestamp 1713400504
transform 1 0 2976 0 -1 2970
box -8 -3 16 105
use FILL  FILL_5
timestamp 1713400504
transform 1 0 2968 0 -1 2970
box -8 -3 16 105
use FILL  FILL_6
timestamp 1713400504
transform 1 0 2960 0 -1 2970
box -8 -3 16 105
use FILL  FILL_7
timestamp 1713400504
transform 1 0 2952 0 -1 2970
box -8 -3 16 105
use FILL  FILL_8
timestamp 1713400504
transform 1 0 2944 0 -1 2970
box -8 -3 16 105
use FILL  FILL_9
timestamp 1713400504
transform 1 0 2936 0 -1 2970
box -8 -3 16 105
use FILL  FILL_10
timestamp 1713400504
transform 1 0 2928 0 -1 2970
box -8 -3 16 105
use FILL  FILL_11
timestamp 1713400504
transform 1 0 2920 0 -1 2970
box -8 -3 16 105
use FILL  FILL_12
timestamp 1713400504
transform 1 0 2912 0 -1 2970
box -8 -3 16 105
use FILL  FILL_13
timestamp 1713400504
transform 1 0 2904 0 -1 2970
box -8 -3 16 105
use FILL  FILL_14
timestamp 1713400504
transform 1 0 2896 0 -1 2970
box -8 -3 16 105
use FILL  FILL_15
timestamp 1713400504
transform 1 0 2888 0 -1 2970
box -8 -3 16 105
use FILL  FILL_16
timestamp 1713400504
transform 1 0 2880 0 -1 2970
box -8 -3 16 105
use FILL  FILL_17
timestamp 1713400504
transform 1 0 2872 0 -1 2970
box -8 -3 16 105
use FILL  FILL_18
timestamp 1713400504
transform 1 0 2864 0 -1 2970
box -8 -3 16 105
use FILL  FILL_19
timestamp 1713400504
transform 1 0 2856 0 -1 2970
box -8 -3 16 105
use FILL  FILL_20
timestamp 1713400504
transform 1 0 2848 0 -1 2970
box -8 -3 16 105
use FILL  FILL_21
timestamp 1713400504
transform 1 0 2840 0 -1 2970
box -8 -3 16 105
use FILL  FILL_22
timestamp 1713400504
transform 1 0 2832 0 -1 2970
box -8 -3 16 105
use FILL  FILL_23
timestamp 1713400504
transform 1 0 2824 0 -1 2970
box -8 -3 16 105
use FILL  FILL_24
timestamp 1713400504
transform 1 0 2816 0 -1 2970
box -8 -3 16 105
use FILL  FILL_25
timestamp 1713400504
transform 1 0 2808 0 -1 2970
box -8 -3 16 105
use FILL  FILL_26
timestamp 1713400504
transform 1 0 2800 0 -1 2970
box -8 -3 16 105
use FILL  FILL_27
timestamp 1713400504
transform 1 0 2792 0 -1 2970
box -8 -3 16 105
use FILL  FILL_28
timestamp 1713400504
transform 1 0 2784 0 -1 2970
box -8 -3 16 105
use FILL  FILL_29
timestamp 1713400504
transform 1 0 2736 0 -1 2970
box -8 -3 16 105
use FILL  FILL_30
timestamp 1713400504
transform 1 0 2728 0 -1 2970
box -8 -3 16 105
use FILL  FILL_31
timestamp 1713400504
transform 1 0 2720 0 -1 2970
box -8 -3 16 105
use FILL  FILL_32
timestamp 1713400504
transform 1 0 2696 0 -1 2970
box -8 -3 16 105
use FILL  FILL_33
timestamp 1713400504
transform 1 0 2688 0 -1 2970
box -8 -3 16 105
use FILL  FILL_34
timestamp 1713400504
transform 1 0 2488 0 -1 2970
box -8 -3 16 105
use FILL  FILL_35
timestamp 1713400504
transform 1 0 2480 0 -1 2970
box -8 -3 16 105
use FILL  FILL_36
timestamp 1713400504
transform 1 0 2472 0 -1 2970
box -8 -3 16 105
use FILL  FILL_37
timestamp 1713400504
transform 1 0 2424 0 -1 2970
box -8 -3 16 105
use FILL  FILL_38
timestamp 1713400504
transform 1 0 2416 0 -1 2970
box -8 -3 16 105
use FILL  FILL_39
timestamp 1713400504
transform 1 0 2408 0 -1 2970
box -8 -3 16 105
use FILL  FILL_40
timestamp 1713400504
transform 1 0 2208 0 -1 2970
box -8 -3 16 105
use FILL  FILL_41
timestamp 1713400504
transform 1 0 2200 0 -1 2970
box -8 -3 16 105
use FILL  FILL_42
timestamp 1713400504
transform 1 0 2192 0 -1 2970
box -8 -3 16 105
use FILL  FILL_43
timestamp 1713400504
transform 1 0 2144 0 -1 2970
box -8 -3 16 105
use FILL  FILL_44
timestamp 1713400504
transform 1 0 2136 0 -1 2970
box -8 -3 16 105
use FILL  FILL_45
timestamp 1713400504
transform 1 0 2032 0 -1 2970
box -8 -3 16 105
use FILL  FILL_46
timestamp 1713400504
transform 1 0 2024 0 -1 2970
box -8 -3 16 105
use FILL  FILL_47
timestamp 1713400504
transform 1 0 1976 0 -1 2970
box -8 -3 16 105
use FILL  FILL_48
timestamp 1713400504
transform 1 0 1968 0 -1 2970
box -8 -3 16 105
use FILL  FILL_49
timestamp 1713400504
transform 1 0 1960 0 -1 2970
box -8 -3 16 105
use FILL  FILL_50
timestamp 1713400504
transform 1 0 1936 0 -1 2970
box -8 -3 16 105
use FILL  FILL_51
timestamp 1713400504
transform 1 0 1832 0 -1 2970
box -8 -3 16 105
use FILL  FILL_52
timestamp 1713400504
transform 1 0 1824 0 -1 2970
box -8 -3 16 105
use FILL  FILL_53
timestamp 1713400504
transform 1 0 1776 0 -1 2970
box -8 -3 16 105
use FILL  FILL_54
timestamp 1713400504
transform 1 0 1768 0 -1 2970
box -8 -3 16 105
use FILL  FILL_55
timestamp 1713400504
transform 1 0 1744 0 -1 2970
box -8 -3 16 105
use FILL  FILL_56
timestamp 1713400504
transform 1 0 1544 0 -1 2970
box -8 -3 16 105
use FILL  FILL_57
timestamp 1713400504
transform 1 0 1424 0 -1 2970
box -8 -3 16 105
use FILL  FILL_58
timestamp 1713400504
transform 1 0 1400 0 -1 2970
box -8 -3 16 105
use FILL  FILL_59
timestamp 1713400504
transform 1 0 1392 0 -1 2970
box -8 -3 16 105
use FILL  FILL_60
timestamp 1713400504
transform 1 0 1384 0 -1 2970
box -8 -3 16 105
use FILL  FILL_61
timestamp 1713400504
transform 1 0 1376 0 -1 2970
box -8 -3 16 105
use FILL  FILL_62
timestamp 1713400504
transform 1 0 1368 0 -1 2970
box -8 -3 16 105
use FILL  FILL_63
timestamp 1713400504
transform 1 0 1320 0 -1 2970
box -8 -3 16 105
use FILL  FILL_64
timestamp 1713400504
transform 1 0 1312 0 -1 2970
box -8 -3 16 105
use FILL  FILL_65
timestamp 1713400504
transform 1 0 1304 0 -1 2970
box -8 -3 16 105
use FILL  FILL_66
timestamp 1713400504
transform 1 0 1280 0 -1 2970
box -8 -3 16 105
use FILL  FILL_67
timestamp 1713400504
transform 1 0 1272 0 -1 2970
box -8 -3 16 105
use FILL  FILL_68
timestamp 1713400504
transform 1 0 1264 0 -1 2970
box -8 -3 16 105
use FILL  FILL_69
timestamp 1713400504
transform 1 0 1256 0 -1 2970
box -8 -3 16 105
use FILL  FILL_70
timestamp 1713400504
transform 1 0 1208 0 -1 2970
box -8 -3 16 105
use FILL  FILL_71
timestamp 1713400504
transform 1 0 1200 0 -1 2970
box -8 -3 16 105
use FILL  FILL_72
timestamp 1713400504
transform 1 0 1192 0 -1 2970
box -8 -3 16 105
use FILL  FILL_73
timestamp 1713400504
transform 1 0 1184 0 -1 2970
box -8 -3 16 105
use FILL  FILL_74
timestamp 1713400504
transform 1 0 1160 0 -1 2970
box -8 -3 16 105
use FILL  FILL_75
timestamp 1713400504
transform 1 0 960 0 -1 2970
box -8 -3 16 105
use FILL  FILL_76
timestamp 1713400504
transform 1 0 920 0 -1 2970
box -8 -3 16 105
use FILL  FILL_77
timestamp 1713400504
transform 1 0 832 0 -1 2970
box -8 -3 16 105
use FILL  FILL_78
timestamp 1713400504
transform 1 0 824 0 -1 2970
box -8 -3 16 105
use FILL  FILL_79
timestamp 1713400504
transform 1 0 768 0 -1 2970
box -8 -3 16 105
use FILL  FILL_80
timestamp 1713400504
transform 1 0 760 0 -1 2970
box -8 -3 16 105
use FILL  FILL_81
timestamp 1713400504
transform 1 0 672 0 -1 2970
box -8 -3 16 105
use FILL  FILL_82
timestamp 1713400504
transform 1 0 664 0 -1 2970
box -8 -3 16 105
use FILL  FILL_83
timestamp 1713400504
transform 1 0 608 0 -1 2970
box -8 -3 16 105
use FILL  FILL_84
timestamp 1713400504
transform 1 0 600 0 -1 2970
box -8 -3 16 105
use FILL  FILL_85
timestamp 1713400504
transform 1 0 592 0 -1 2970
box -8 -3 16 105
use FILL  FILL_86
timestamp 1713400504
transform 1 0 560 0 -1 2970
box -8 -3 16 105
use FILL  FILL_87
timestamp 1713400504
transform 1 0 552 0 -1 2970
box -8 -3 16 105
use FILL  FILL_88
timestamp 1713400504
transform 1 0 544 0 -1 2970
box -8 -3 16 105
use FILL  FILL_89
timestamp 1713400504
transform 1 0 536 0 -1 2970
box -8 -3 16 105
use FILL  FILL_90
timestamp 1713400504
transform 1 0 528 0 -1 2970
box -8 -3 16 105
use FILL  FILL_91
timestamp 1713400504
transform 1 0 520 0 -1 2970
box -8 -3 16 105
use FILL  FILL_92
timestamp 1713400504
transform 1 0 480 0 -1 2970
box -8 -3 16 105
use FILL  FILL_93
timestamp 1713400504
transform 1 0 472 0 -1 2970
box -8 -3 16 105
use FILL  FILL_94
timestamp 1713400504
transform 1 0 464 0 -1 2970
box -8 -3 16 105
use FILL  FILL_95
timestamp 1713400504
transform 1 0 456 0 -1 2970
box -8 -3 16 105
use FILL  FILL_96
timestamp 1713400504
transform 1 0 416 0 -1 2970
box -8 -3 16 105
use FILL  FILL_97
timestamp 1713400504
transform 1 0 408 0 -1 2970
box -8 -3 16 105
use FILL  FILL_98
timestamp 1713400504
transform 1 0 400 0 -1 2970
box -8 -3 16 105
use FILL  FILL_99
timestamp 1713400504
transform 1 0 312 0 -1 2970
box -8 -3 16 105
use FILL  FILL_100
timestamp 1713400504
transform 1 0 304 0 -1 2970
box -8 -3 16 105
use FILL  FILL_101
timestamp 1713400504
transform 1 0 296 0 -1 2970
box -8 -3 16 105
use FILL  FILL_102
timestamp 1713400504
transform 1 0 240 0 -1 2970
box -8 -3 16 105
use FILL  FILL_103
timestamp 1713400504
transform 1 0 232 0 -1 2970
box -8 -3 16 105
use FILL  FILL_104
timestamp 1713400504
transform 1 0 224 0 -1 2970
box -8 -3 16 105
use FILL  FILL_105
timestamp 1713400504
transform 1 0 216 0 -1 2970
box -8 -3 16 105
use FILL  FILL_106
timestamp 1713400504
transform 1 0 208 0 -1 2970
box -8 -3 16 105
use FILL  FILL_107
timestamp 1713400504
transform 1 0 184 0 -1 2970
box -8 -3 16 105
use FILL  FILL_108
timestamp 1713400504
transform 1 0 176 0 -1 2970
box -8 -3 16 105
use FILL  FILL_109
timestamp 1713400504
transform 1 0 136 0 -1 2970
box -8 -3 16 105
use FILL  FILL_110
timestamp 1713400504
transform 1 0 128 0 -1 2970
box -8 -3 16 105
use FILL  FILL_111
timestamp 1713400504
transform 1 0 120 0 -1 2970
box -8 -3 16 105
use FILL  FILL_112
timestamp 1713400504
transform 1 0 112 0 -1 2970
box -8 -3 16 105
use FILL  FILL_113
timestamp 1713400504
transform 1 0 104 0 -1 2970
box -8 -3 16 105
use FILL  FILL_114
timestamp 1713400504
transform 1 0 96 0 -1 2970
box -8 -3 16 105
use FILL  FILL_115
timestamp 1713400504
transform 1 0 88 0 -1 2970
box -8 -3 16 105
use FILL  FILL_116
timestamp 1713400504
transform 1 0 80 0 -1 2970
box -8 -3 16 105
use FILL  FILL_117
timestamp 1713400504
transform 1 0 72 0 -1 2970
box -8 -3 16 105
use FILL  FILL_118
timestamp 1713400504
transform 1 0 3008 0 1 2770
box -8 -3 16 105
use FILL  FILL_119
timestamp 1713400504
transform 1 0 2904 0 1 2770
box -8 -3 16 105
use FILL  FILL_120
timestamp 1713400504
transform 1 0 2800 0 1 2770
box -8 -3 16 105
use FILL  FILL_121
timestamp 1713400504
transform 1 0 2776 0 1 2770
box -8 -3 16 105
use FILL  FILL_122
timestamp 1713400504
transform 1 0 2768 0 1 2770
box -8 -3 16 105
use FILL  FILL_123
timestamp 1713400504
transform 1 0 2760 0 1 2770
box -8 -3 16 105
use FILL  FILL_124
timestamp 1713400504
transform 1 0 2752 0 1 2770
box -8 -3 16 105
use FILL  FILL_125
timestamp 1713400504
transform 1 0 2744 0 1 2770
box -8 -3 16 105
use FILL  FILL_126
timestamp 1713400504
transform 1 0 2696 0 1 2770
box -8 -3 16 105
use FILL  FILL_127
timestamp 1713400504
transform 1 0 2688 0 1 2770
box -8 -3 16 105
use FILL  FILL_128
timestamp 1713400504
transform 1 0 2680 0 1 2770
box -8 -3 16 105
use FILL  FILL_129
timestamp 1713400504
transform 1 0 2672 0 1 2770
box -8 -3 16 105
use FILL  FILL_130
timestamp 1713400504
transform 1 0 2664 0 1 2770
box -8 -3 16 105
use FILL  FILL_131
timestamp 1713400504
transform 1 0 2624 0 1 2770
box -8 -3 16 105
use FILL  FILL_132
timestamp 1713400504
transform 1 0 2616 0 1 2770
box -8 -3 16 105
use FILL  FILL_133
timestamp 1713400504
transform 1 0 2608 0 1 2770
box -8 -3 16 105
use FILL  FILL_134
timestamp 1713400504
transform 1 0 2600 0 1 2770
box -8 -3 16 105
use FILL  FILL_135
timestamp 1713400504
transform 1 0 2560 0 1 2770
box -8 -3 16 105
use FILL  FILL_136
timestamp 1713400504
transform 1 0 2552 0 1 2770
box -8 -3 16 105
use FILL  FILL_137
timestamp 1713400504
transform 1 0 2544 0 1 2770
box -8 -3 16 105
use FILL  FILL_138
timestamp 1713400504
transform 1 0 2520 0 1 2770
box -8 -3 16 105
use FILL  FILL_139
timestamp 1713400504
transform 1 0 2512 0 1 2770
box -8 -3 16 105
use FILL  FILL_140
timestamp 1713400504
transform 1 0 2488 0 1 2770
box -8 -3 16 105
use FILL  FILL_141
timestamp 1713400504
transform 1 0 2480 0 1 2770
box -8 -3 16 105
use FILL  FILL_142
timestamp 1713400504
transform 1 0 2472 0 1 2770
box -8 -3 16 105
use FILL  FILL_143
timestamp 1713400504
transform 1 0 2464 0 1 2770
box -8 -3 16 105
use FILL  FILL_144
timestamp 1713400504
transform 1 0 2456 0 1 2770
box -8 -3 16 105
use FILL  FILL_145
timestamp 1713400504
transform 1 0 2416 0 1 2770
box -8 -3 16 105
use FILL  FILL_146
timestamp 1713400504
transform 1 0 2408 0 1 2770
box -8 -3 16 105
use FILL  FILL_147
timestamp 1713400504
transform 1 0 2400 0 1 2770
box -8 -3 16 105
use FILL  FILL_148
timestamp 1713400504
transform 1 0 2376 0 1 2770
box -8 -3 16 105
use FILL  FILL_149
timestamp 1713400504
transform 1 0 2368 0 1 2770
box -8 -3 16 105
use FILL  FILL_150
timestamp 1713400504
transform 1 0 2360 0 1 2770
box -8 -3 16 105
use FILL  FILL_151
timestamp 1713400504
transform 1 0 2320 0 1 2770
box -8 -3 16 105
use FILL  FILL_152
timestamp 1713400504
transform 1 0 2312 0 1 2770
box -8 -3 16 105
use FILL  FILL_153
timestamp 1713400504
transform 1 0 2304 0 1 2770
box -8 -3 16 105
use FILL  FILL_154
timestamp 1713400504
transform 1 0 2280 0 1 2770
box -8 -3 16 105
use FILL  FILL_155
timestamp 1713400504
transform 1 0 2272 0 1 2770
box -8 -3 16 105
use FILL  FILL_156
timestamp 1713400504
transform 1 0 2264 0 1 2770
box -8 -3 16 105
use FILL  FILL_157
timestamp 1713400504
transform 1 0 2256 0 1 2770
box -8 -3 16 105
use FILL  FILL_158
timestamp 1713400504
transform 1 0 2216 0 1 2770
box -8 -3 16 105
use FILL  FILL_159
timestamp 1713400504
transform 1 0 2208 0 1 2770
box -8 -3 16 105
use FILL  FILL_160
timestamp 1713400504
transform 1 0 2184 0 1 2770
box -8 -3 16 105
use FILL  FILL_161
timestamp 1713400504
transform 1 0 2176 0 1 2770
box -8 -3 16 105
use FILL  FILL_162
timestamp 1713400504
transform 1 0 2168 0 1 2770
box -8 -3 16 105
use FILL  FILL_163
timestamp 1713400504
transform 1 0 2160 0 1 2770
box -8 -3 16 105
use FILL  FILL_164
timestamp 1713400504
transform 1 0 2120 0 1 2770
box -8 -3 16 105
use FILL  FILL_165
timestamp 1713400504
transform 1 0 2112 0 1 2770
box -8 -3 16 105
use FILL  FILL_166
timestamp 1713400504
transform 1 0 2088 0 1 2770
box -8 -3 16 105
use FILL  FILL_167
timestamp 1713400504
transform 1 0 2080 0 1 2770
box -8 -3 16 105
use FILL  FILL_168
timestamp 1713400504
transform 1 0 1976 0 1 2770
box -8 -3 16 105
use FILL  FILL_169
timestamp 1713400504
transform 1 0 1968 0 1 2770
box -8 -3 16 105
use FILL  FILL_170
timestamp 1713400504
transform 1 0 1960 0 1 2770
box -8 -3 16 105
use FILL  FILL_171
timestamp 1713400504
transform 1 0 1920 0 1 2770
box -8 -3 16 105
use FILL  FILL_172
timestamp 1713400504
transform 1 0 1912 0 1 2770
box -8 -3 16 105
use FILL  FILL_173
timestamp 1713400504
transform 1 0 1904 0 1 2770
box -8 -3 16 105
use FILL  FILL_174
timestamp 1713400504
transform 1 0 1896 0 1 2770
box -8 -3 16 105
use FILL  FILL_175
timestamp 1713400504
transform 1 0 1888 0 1 2770
box -8 -3 16 105
use FILL  FILL_176
timestamp 1713400504
transform 1 0 1856 0 1 2770
box -8 -3 16 105
use FILL  FILL_177
timestamp 1713400504
transform 1 0 1848 0 1 2770
box -8 -3 16 105
use FILL  FILL_178
timestamp 1713400504
transform 1 0 1840 0 1 2770
box -8 -3 16 105
use FILL  FILL_179
timestamp 1713400504
transform 1 0 1808 0 1 2770
box -8 -3 16 105
use FILL  FILL_180
timestamp 1713400504
transform 1 0 1800 0 1 2770
box -8 -3 16 105
use FILL  FILL_181
timestamp 1713400504
transform 1 0 1792 0 1 2770
box -8 -3 16 105
use FILL  FILL_182
timestamp 1713400504
transform 1 0 1784 0 1 2770
box -8 -3 16 105
use FILL  FILL_183
timestamp 1713400504
transform 1 0 1752 0 1 2770
box -8 -3 16 105
use FILL  FILL_184
timestamp 1713400504
transform 1 0 1744 0 1 2770
box -8 -3 16 105
use FILL  FILL_185
timestamp 1713400504
transform 1 0 1736 0 1 2770
box -8 -3 16 105
use FILL  FILL_186
timestamp 1713400504
transform 1 0 1728 0 1 2770
box -8 -3 16 105
use FILL  FILL_187
timestamp 1713400504
transform 1 0 1720 0 1 2770
box -8 -3 16 105
use FILL  FILL_188
timestamp 1713400504
transform 1 0 1712 0 1 2770
box -8 -3 16 105
use FILL  FILL_189
timestamp 1713400504
transform 1 0 1664 0 1 2770
box -8 -3 16 105
use FILL  FILL_190
timestamp 1713400504
transform 1 0 1656 0 1 2770
box -8 -3 16 105
use FILL  FILL_191
timestamp 1713400504
transform 1 0 1648 0 1 2770
box -8 -3 16 105
use FILL  FILL_192
timestamp 1713400504
transform 1 0 1640 0 1 2770
box -8 -3 16 105
use FILL  FILL_193
timestamp 1713400504
transform 1 0 1632 0 1 2770
box -8 -3 16 105
use FILL  FILL_194
timestamp 1713400504
transform 1 0 1528 0 1 2770
box -8 -3 16 105
use FILL  FILL_195
timestamp 1713400504
transform 1 0 1520 0 1 2770
box -8 -3 16 105
use FILL  FILL_196
timestamp 1713400504
transform 1 0 1512 0 1 2770
box -8 -3 16 105
use FILL  FILL_197
timestamp 1713400504
transform 1 0 1504 0 1 2770
box -8 -3 16 105
use FILL  FILL_198
timestamp 1713400504
transform 1 0 1480 0 1 2770
box -8 -3 16 105
use FILL  FILL_199
timestamp 1713400504
transform 1 0 1472 0 1 2770
box -8 -3 16 105
use FILL  FILL_200
timestamp 1713400504
transform 1 0 1464 0 1 2770
box -8 -3 16 105
use FILL  FILL_201
timestamp 1713400504
transform 1 0 1456 0 1 2770
box -8 -3 16 105
use FILL  FILL_202
timestamp 1713400504
transform 1 0 1448 0 1 2770
box -8 -3 16 105
use FILL  FILL_203
timestamp 1713400504
transform 1 0 1400 0 1 2770
box -8 -3 16 105
use FILL  FILL_204
timestamp 1713400504
transform 1 0 1392 0 1 2770
box -8 -3 16 105
use FILL  FILL_205
timestamp 1713400504
transform 1 0 1384 0 1 2770
box -8 -3 16 105
use FILL  FILL_206
timestamp 1713400504
transform 1 0 1376 0 1 2770
box -8 -3 16 105
use FILL  FILL_207
timestamp 1713400504
transform 1 0 1368 0 1 2770
box -8 -3 16 105
use FILL  FILL_208
timestamp 1713400504
transform 1 0 1360 0 1 2770
box -8 -3 16 105
use FILL  FILL_209
timestamp 1713400504
transform 1 0 1328 0 1 2770
box -8 -3 16 105
use FILL  FILL_210
timestamp 1713400504
transform 1 0 1320 0 1 2770
box -8 -3 16 105
use FILL  FILL_211
timestamp 1713400504
transform 1 0 1312 0 1 2770
box -8 -3 16 105
use FILL  FILL_212
timestamp 1713400504
transform 1 0 1304 0 1 2770
box -8 -3 16 105
use FILL  FILL_213
timestamp 1713400504
transform 1 0 1296 0 1 2770
box -8 -3 16 105
use FILL  FILL_214
timestamp 1713400504
transform 1 0 1256 0 1 2770
box -8 -3 16 105
use FILL  FILL_215
timestamp 1713400504
transform 1 0 1248 0 1 2770
box -8 -3 16 105
use FILL  FILL_216
timestamp 1713400504
transform 1 0 1240 0 1 2770
box -8 -3 16 105
use FILL  FILL_217
timestamp 1713400504
transform 1 0 1232 0 1 2770
box -8 -3 16 105
use FILL  FILL_218
timestamp 1713400504
transform 1 0 1224 0 1 2770
box -8 -3 16 105
use FILL  FILL_219
timestamp 1713400504
transform 1 0 1216 0 1 2770
box -8 -3 16 105
use FILL  FILL_220
timestamp 1713400504
transform 1 0 1208 0 1 2770
box -8 -3 16 105
use FILL  FILL_221
timestamp 1713400504
transform 1 0 1168 0 1 2770
box -8 -3 16 105
use FILL  FILL_222
timestamp 1713400504
transform 1 0 1160 0 1 2770
box -8 -3 16 105
use FILL  FILL_223
timestamp 1713400504
transform 1 0 1152 0 1 2770
box -8 -3 16 105
use FILL  FILL_224
timestamp 1713400504
transform 1 0 1144 0 1 2770
box -8 -3 16 105
use FILL  FILL_225
timestamp 1713400504
transform 1 0 1136 0 1 2770
box -8 -3 16 105
use FILL  FILL_226
timestamp 1713400504
transform 1 0 1128 0 1 2770
box -8 -3 16 105
use FILL  FILL_227
timestamp 1713400504
transform 1 0 1104 0 1 2770
box -8 -3 16 105
use FILL  FILL_228
timestamp 1713400504
transform 1 0 1096 0 1 2770
box -8 -3 16 105
use FILL  FILL_229
timestamp 1713400504
transform 1 0 1088 0 1 2770
box -8 -3 16 105
use FILL  FILL_230
timestamp 1713400504
transform 1 0 1080 0 1 2770
box -8 -3 16 105
use FILL  FILL_231
timestamp 1713400504
transform 1 0 1072 0 1 2770
box -8 -3 16 105
use FILL  FILL_232
timestamp 1713400504
transform 1 0 1064 0 1 2770
box -8 -3 16 105
use FILL  FILL_233
timestamp 1713400504
transform 1 0 1056 0 1 2770
box -8 -3 16 105
use FILL  FILL_234
timestamp 1713400504
transform 1 0 1048 0 1 2770
box -8 -3 16 105
use FILL  FILL_235
timestamp 1713400504
transform 1 0 1040 0 1 2770
box -8 -3 16 105
use FILL  FILL_236
timestamp 1713400504
transform 1 0 1032 0 1 2770
box -8 -3 16 105
use FILL  FILL_237
timestamp 1713400504
transform 1 0 1024 0 1 2770
box -8 -3 16 105
use FILL  FILL_238
timestamp 1713400504
transform 1 0 1016 0 1 2770
box -8 -3 16 105
use FILL  FILL_239
timestamp 1713400504
transform 1 0 992 0 1 2770
box -8 -3 16 105
use FILL  FILL_240
timestamp 1713400504
transform 1 0 984 0 1 2770
box -8 -3 16 105
use FILL  FILL_241
timestamp 1713400504
transform 1 0 976 0 1 2770
box -8 -3 16 105
use FILL  FILL_242
timestamp 1713400504
transform 1 0 968 0 1 2770
box -8 -3 16 105
use FILL  FILL_243
timestamp 1713400504
transform 1 0 960 0 1 2770
box -8 -3 16 105
use FILL  FILL_244
timestamp 1713400504
transform 1 0 952 0 1 2770
box -8 -3 16 105
use FILL  FILL_245
timestamp 1713400504
transform 1 0 896 0 1 2770
box -8 -3 16 105
use FILL  FILL_246
timestamp 1713400504
transform 1 0 888 0 1 2770
box -8 -3 16 105
use FILL  FILL_247
timestamp 1713400504
transform 1 0 880 0 1 2770
box -8 -3 16 105
use FILL  FILL_248
timestamp 1713400504
transform 1 0 856 0 1 2770
box -8 -3 16 105
use FILL  FILL_249
timestamp 1713400504
transform 1 0 848 0 1 2770
box -8 -3 16 105
use FILL  FILL_250
timestamp 1713400504
transform 1 0 840 0 1 2770
box -8 -3 16 105
use FILL  FILL_251
timestamp 1713400504
transform 1 0 832 0 1 2770
box -8 -3 16 105
use FILL  FILL_252
timestamp 1713400504
transform 1 0 776 0 1 2770
box -8 -3 16 105
use FILL  FILL_253
timestamp 1713400504
transform 1 0 768 0 1 2770
box -8 -3 16 105
use FILL  FILL_254
timestamp 1713400504
transform 1 0 760 0 1 2770
box -8 -3 16 105
use FILL  FILL_255
timestamp 1713400504
transform 1 0 752 0 1 2770
box -8 -3 16 105
use FILL  FILL_256
timestamp 1713400504
transform 1 0 728 0 1 2770
box -8 -3 16 105
use FILL  FILL_257
timestamp 1713400504
transform 1 0 720 0 1 2770
box -8 -3 16 105
use FILL  FILL_258
timestamp 1713400504
transform 1 0 712 0 1 2770
box -8 -3 16 105
use FILL  FILL_259
timestamp 1713400504
transform 1 0 656 0 1 2770
box -8 -3 16 105
use FILL  FILL_260
timestamp 1713400504
transform 1 0 648 0 1 2770
box -8 -3 16 105
use FILL  FILL_261
timestamp 1713400504
transform 1 0 640 0 1 2770
box -8 -3 16 105
use FILL  FILL_262
timestamp 1713400504
transform 1 0 632 0 1 2770
box -8 -3 16 105
use FILL  FILL_263
timestamp 1713400504
transform 1 0 552 0 1 2770
box -8 -3 16 105
use FILL  FILL_264
timestamp 1713400504
transform 1 0 544 0 1 2770
box -8 -3 16 105
use FILL  FILL_265
timestamp 1713400504
transform 1 0 536 0 1 2770
box -8 -3 16 105
use FILL  FILL_266
timestamp 1713400504
transform 1 0 528 0 1 2770
box -8 -3 16 105
use FILL  FILL_267
timestamp 1713400504
transform 1 0 472 0 1 2770
box -8 -3 16 105
use FILL  FILL_268
timestamp 1713400504
transform 1 0 464 0 1 2770
box -8 -3 16 105
use FILL  FILL_269
timestamp 1713400504
transform 1 0 456 0 1 2770
box -8 -3 16 105
use FILL  FILL_270
timestamp 1713400504
transform 1 0 432 0 1 2770
box -8 -3 16 105
use FILL  FILL_271
timestamp 1713400504
transform 1 0 424 0 1 2770
box -8 -3 16 105
use FILL  FILL_272
timestamp 1713400504
transform 1 0 336 0 1 2770
box -8 -3 16 105
use FILL  FILL_273
timestamp 1713400504
transform 1 0 328 0 1 2770
box -8 -3 16 105
use FILL  FILL_274
timestamp 1713400504
transform 1 0 272 0 1 2770
box -8 -3 16 105
use FILL  FILL_275
timestamp 1713400504
transform 1 0 264 0 1 2770
box -8 -3 16 105
use FILL  FILL_276
timestamp 1713400504
transform 1 0 256 0 1 2770
box -8 -3 16 105
use FILL  FILL_277
timestamp 1713400504
transform 1 0 232 0 1 2770
box -8 -3 16 105
use FILL  FILL_278
timestamp 1713400504
transform 1 0 224 0 1 2770
box -8 -3 16 105
use FILL  FILL_279
timestamp 1713400504
transform 1 0 136 0 1 2770
box -8 -3 16 105
use FILL  FILL_280
timestamp 1713400504
transform 1 0 128 0 1 2770
box -8 -3 16 105
use FILL  FILL_281
timestamp 1713400504
transform 1 0 72 0 1 2770
box -8 -3 16 105
use FILL  FILL_282
timestamp 1713400504
transform 1 0 3008 0 -1 2770
box -8 -3 16 105
use FILL  FILL_283
timestamp 1713400504
transform 1 0 3000 0 -1 2770
box -8 -3 16 105
use FILL  FILL_284
timestamp 1713400504
transform 1 0 2992 0 -1 2770
box -8 -3 16 105
use FILL  FILL_285
timestamp 1713400504
transform 1 0 2968 0 -1 2770
box -8 -3 16 105
use FILL  FILL_286
timestamp 1713400504
transform 1 0 2960 0 -1 2770
box -8 -3 16 105
use FILL  FILL_287
timestamp 1713400504
transform 1 0 2952 0 -1 2770
box -8 -3 16 105
use FILL  FILL_288
timestamp 1713400504
transform 1 0 2944 0 -1 2770
box -8 -3 16 105
use FILL  FILL_289
timestamp 1713400504
transform 1 0 2936 0 -1 2770
box -8 -3 16 105
use FILL  FILL_290
timestamp 1713400504
transform 1 0 2928 0 -1 2770
box -8 -3 16 105
use FILL  FILL_291
timestamp 1713400504
transform 1 0 2920 0 -1 2770
box -8 -3 16 105
use FILL  FILL_292
timestamp 1713400504
transform 1 0 2872 0 -1 2770
box -8 -3 16 105
use FILL  FILL_293
timestamp 1713400504
transform 1 0 2864 0 -1 2770
box -8 -3 16 105
use FILL  FILL_294
timestamp 1713400504
transform 1 0 2856 0 -1 2770
box -8 -3 16 105
use FILL  FILL_295
timestamp 1713400504
transform 1 0 2848 0 -1 2770
box -8 -3 16 105
use FILL  FILL_296
timestamp 1713400504
transform 1 0 2824 0 -1 2770
box -8 -3 16 105
use FILL  FILL_297
timestamp 1713400504
transform 1 0 2816 0 -1 2770
box -8 -3 16 105
use FILL  FILL_298
timestamp 1713400504
transform 1 0 2808 0 -1 2770
box -8 -3 16 105
use FILL  FILL_299
timestamp 1713400504
transform 1 0 2704 0 -1 2770
box -8 -3 16 105
use FILL  FILL_300
timestamp 1713400504
transform 1 0 2696 0 -1 2770
box -8 -3 16 105
use FILL  FILL_301
timestamp 1713400504
transform 1 0 2688 0 -1 2770
box -8 -3 16 105
use FILL  FILL_302
timestamp 1713400504
transform 1 0 2680 0 -1 2770
box -8 -3 16 105
use FILL  FILL_303
timestamp 1713400504
transform 1 0 2640 0 -1 2770
box -8 -3 16 105
use FILL  FILL_304
timestamp 1713400504
transform 1 0 2608 0 -1 2770
box -8 -3 16 105
use FILL  FILL_305
timestamp 1713400504
transform 1 0 2600 0 -1 2770
box -8 -3 16 105
use FILL  FILL_306
timestamp 1713400504
transform 1 0 2592 0 -1 2770
box -8 -3 16 105
use FILL  FILL_307
timestamp 1713400504
transform 1 0 2584 0 -1 2770
box -8 -3 16 105
use FILL  FILL_308
timestamp 1713400504
transform 1 0 2576 0 -1 2770
box -8 -3 16 105
use FILL  FILL_309
timestamp 1713400504
transform 1 0 2568 0 -1 2770
box -8 -3 16 105
use FILL  FILL_310
timestamp 1713400504
transform 1 0 2520 0 -1 2770
box -8 -3 16 105
use FILL  FILL_311
timestamp 1713400504
transform 1 0 2512 0 -1 2770
box -8 -3 16 105
use FILL  FILL_312
timestamp 1713400504
transform 1 0 2504 0 -1 2770
box -8 -3 16 105
use FILL  FILL_313
timestamp 1713400504
transform 1 0 2496 0 -1 2770
box -8 -3 16 105
use FILL  FILL_314
timestamp 1713400504
transform 1 0 2488 0 -1 2770
box -8 -3 16 105
use FILL  FILL_315
timestamp 1713400504
transform 1 0 2448 0 -1 2770
box -8 -3 16 105
use FILL  FILL_316
timestamp 1713400504
transform 1 0 2440 0 -1 2770
box -8 -3 16 105
use FILL  FILL_317
timestamp 1713400504
transform 1 0 2432 0 -1 2770
box -8 -3 16 105
use FILL  FILL_318
timestamp 1713400504
transform 1 0 2424 0 -1 2770
box -8 -3 16 105
use FILL  FILL_319
timestamp 1713400504
transform 1 0 2416 0 -1 2770
box -8 -3 16 105
use FILL  FILL_320
timestamp 1713400504
transform 1 0 2368 0 -1 2770
box -8 -3 16 105
use FILL  FILL_321
timestamp 1713400504
transform 1 0 2360 0 -1 2770
box -8 -3 16 105
use FILL  FILL_322
timestamp 1713400504
transform 1 0 2352 0 -1 2770
box -8 -3 16 105
use FILL  FILL_323
timestamp 1713400504
transform 1 0 2344 0 -1 2770
box -8 -3 16 105
use FILL  FILL_324
timestamp 1713400504
transform 1 0 2336 0 -1 2770
box -8 -3 16 105
use FILL  FILL_325
timestamp 1713400504
transform 1 0 2296 0 -1 2770
box -8 -3 16 105
use FILL  FILL_326
timestamp 1713400504
transform 1 0 2192 0 -1 2770
box -8 -3 16 105
use FILL  FILL_327
timestamp 1713400504
transform 1 0 2184 0 -1 2770
box -8 -3 16 105
use FILL  FILL_328
timestamp 1713400504
transform 1 0 2176 0 -1 2770
box -8 -3 16 105
use FILL  FILL_329
timestamp 1713400504
transform 1 0 2144 0 -1 2770
box -8 -3 16 105
use FILL  FILL_330
timestamp 1713400504
transform 1 0 2136 0 -1 2770
box -8 -3 16 105
use FILL  FILL_331
timestamp 1713400504
transform 1 0 2096 0 -1 2770
box -8 -3 16 105
use FILL  FILL_332
timestamp 1713400504
transform 1 0 2088 0 -1 2770
box -8 -3 16 105
use FILL  FILL_333
timestamp 1713400504
transform 1 0 2080 0 -1 2770
box -8 -3 16 105
use FILL  FILL_334
timestamp 1713400504
transform 1 0 1976 0 -1 2770
box -8 -3 16 105
use FILL  FILL_335
timestamp 1713400504
transform 1 0 1968 0 -1 2770
box -8 -3 16 105
use FILL  FILL_336
timestamp 1713400504
transform 1 0 1960 0 -1 2770
box -8 -3 16 105
use FILL  FILL_337
timestamp 1713400504
transform 1 0 1912 0 -1 2770
box -8 -3 16 105
use FILL  FILL_338
timestamp 1713400504
transform 1 0 1904 0 -1 2770
box -8 -3 16 105
use FILL  FILL_339
timestamp 1713400504
transform 1 0 1896 0 -1 2770
box -8 -3 16 105
use FILL  FILL_340
timestamp 1713400504
transform 1 0 1888 0 -1 2770
box -8 -3 16 105
use FILL  FILL_341
timestamp 1713400504
transform 1 0 1880 0 -1 2770
box -8 -3 16 105
use FILL  FILL_342
timestamp 1713400504
transform 1 0 1872 0 -1 2770
box -8 -3 16 105
use FILL  FILL_343
timestamp 1713400504
transform 1 0 1824 0 -1 2770
box -8 -3 16 105
use FILL  FILL_344
timestamp 1713400504
transform 1 0 1816 0 -1 2770
box -8 -3 16 105
use FILL  FILL_345
timestamp 1713400504
transform 1 0 1808 0 -1 2770
box -8 -3 16 105
use FILL  FILL_346
timestamp 1713400504
transform 1 0 1800 0 -1 2770
box -8 -3 16 105
use FILL  FILL_347
timestamp 1713400504
transform 1 0 1792 0 -1 2770
box -8 -3 16 105
use FILL  FILL_348
timestamp 1713400504
transform 1 0 1784 0 -1 2770
box -8 -3 16 105
use FILL  FILL_349
timestamp 1713400504
transform 1 0 1736 0 -1 2770
box -8 -3 16 105
use FILL  FILL_350
timestamp 1713400504
transform 1 0 1728 0 -1 2770
box -8 -3 16 105
use FILL  FILL_351
timestamp 1713400504
transform 1 0 1720 0 -1 2770
box -8 -3 16 105
use FILL  FILL_352
timestamp 1713400504
transform 1 0 1712 0 -1 2770
box -8 -3 16 105
use FILL  FILL_353
timestamp 1713400504
transform 1 0 1704 0 -1 2770
box -8 -3 16 105
use FILL  FILL_354
timestamp 1713400504
transform 1 0 1680 0 -1 2770
box -8 -3 16 105
use FILL  FILL_355
timestamp 1713400504
transform 1 0 1672 0 -1 2770
box -8 -3 16 105
use FILL  FILL_356
timestamp 1713400504
transform 1 0 1632 0 -1 2770
box -8 -3 16 105
use FILL  FILL_357
timestamp 1713400504
transform 1 0 1624 0 -1 2770
box -8 -3 16 105
use FILL  FILL_358
timestamp 1713400504
transform 1 0 1616 0 -1 2770
box -8 -3 16 105
use FILL  FILL_359
timestamp 1713400504
transform 1 0 1608 0 -1 2770
box -8 -3 16 105
use FILL  FILL_360
timestamp 1713400504
transform 1 0 1568 0 -1 2770
box -8 -3 16 105
use FILL  FILL_361
timestamp 1713400504
transform 1 0 1560 0 -1 2770
box -8 -3 16 105
use FILL  FILL_362
timestamp 1713400504
transform 1 0 1552 0 -1 2770
box -8 -3 16 105
use FILL  FILL_363
timestamp 1713400504
transform 1 0 1544 0 -1 2770
box -8 -3 16 105
use FILL  FILL_364
timestamp 1713400504
transform 1 0 1504 0 -1 2770
box -8 -3 16 105
use FILL  FILL_365
timestamp 1713400504
transform 1 0 1496 0 -1 2770
box -8 -3 16 105
use FILL  FILL_366
timestamp 1713400504
transform 1 0 1488 0 -1 2770
box -8 -3 16 105
use FILL  FILL_367
timestamp 1713400504
transform 1 0 1448 0 -1 2770
box -8 -3 16 105
use FILL  FILL_368
timestamp 1713400504
transform 1 0 1440 0 -1 2770
box -8 -3 16 105
use FILL  FILL_369
timestamp 1713400504
transform 1 0 1432 0 -1 2770
box -8 -3 16 105
use FILL  FILL_370
timestamp 1713400504
transform 1 0 1424 0 -1 2770
box -8 -3 16 105
use FILL  FILL_371
timestamp 1713400504
transform 1 0 1400 0 -1 2770
box -8 -3 16 105
use FILL  FILL_372
timestamp 1713400504
transform 1 0 1392 0 -1 2770
box -8 -3 16 105
use FILL  FILL_373
timestamp 1713400504
transform 1 0 1352 0 -1 2770
box -8 -3 16 105
use FILL  FILL_374
timestamp 1713400504
transform 1 0 1344 0 -1 2770
box -8 -3 16 105
use FILL  FILL_375
timestamp 1713400504
transform 1 0 1336 0 -1 2770
box -8 -3 16 105
use FILL  FILL_376
timestamp 1713400504
transform 1 0 1328 0 -1 2770
box -8 -3 16 105
use FILL  FILL_377
timestamp 1713400504
transform 1 0 1296 0 -1 2770
box -8 -3 16 105
use FILL  FILL_378
timestamp 1713400504
transform 1 0 1288 0 -1 2770
box -8 -3 16 105
use FILL  FILL_379
timestamp 1713400504
transform 1 0 1280 0 -1 2770
box -8 -3 16 105
use FILL  FILL_380
timestamp 1713400504
transform 1 0 1272 0 -1 2770
box -8 -3 16 105
use FILL  FILL_381
timestamp 1713400504
transform 1 0 1232 0 -1 2770
box -8 -3 16 105
use FILL  FILL_382
timestamp 1713400504
transform 1 0 1224 0 -1 2770
box -8 -3 16 105
use FILL  FILL_383
timestamp 1713400504
transform 1 0 1216 0 -1 2770
box -8 -3 16 105
use FILL  FILL_384
timestamp 1713400504
transform 1 0 1208 0 -1 2770
box -8 -3 16 105
use FILL  FILL_385
timestamp 1713400504
transform 1 0 1168 0 -1 2770
box -8 -3 16 105
use FILL  FILL_386
timestamp 1713400504
transform 1 0 1160 0 -1 2770
box -8 -3 16 105
use FILL  FILL_387
timestamp 1713400504
transform 1 0 1152 0 -1 2770
box -8 -3 16 105
use FILL  FILL_388
timestamp 1713400504
transform 1 0 1144 0 -1 2770
box -8 -3 16 105
use FILL  FILL_389
timestamp 1713400504
transform 1 0 1136 0 -1 2770
box -8 -3 16 105
use FILL  FILL_390
timestamp 1713400504
transform 1 0 1128 0 -1 2770
box -8 -3 16 105
use FILL  FILL_391
timestamp 1713400504
transform 1 0 1080 0 -1 2770
box -8 -3 16 105
use FILL  FILL_392
timestamp 1713400504
transform 1 0 1072 0 -1 2770
box -8 -3 16 105
use FILL  FILL_393
timestamp 1713400504
transform 1 0 1064 0 -1 2770
box -8 -3 16 105
use FILL  FILL_394
timestamp 1713400504
transform 1 0 1056 0 -1 2770
box -8 -3 16 105
use FILL  FILL_395
timestamp 1713400504
transform 1 0 1048 0 -1 2770
box -8 -3 16 105
use FILL  FILL_396
timestamp 1713400504
transform 1 0 992 0 -1 2770
box -8 -3 16 105
use FILL  FILL_397
timestamp 1713400504
transform 1 0 984 0 -1 2770
box -8 -3 16 105
use FILL  FILL_398
timestamp 1713400504
transform 1 0 976 0 -1 2770
box -8 -3 16 105
use FILL  FILL_399
timestamp 1713400504
transform 1 0 944 0 -1 2770
box -8 -3 16 105
use FILL  FILL_400
timestamp 1713400504
transform 1 0 880 0 -1 2770
box -8 -3 16 105
use FILL  FILL_401
timestamp 1713400504
transform 1 0 848 0 -1 2770
box -8 -3 16 105
use FILL  FILL_402
timestamp 1713400504
transform 1 0 840 0 -1 2770
box -8 -3 16 105
use FILL  FILL_403
timestamp 1713400504
transform 1 0 832 0 -1 2770
box -8 -3 16 105
use FILL  FILL_404
timestamp 1713400504
transform 1 0 752 0 -1 2770
box -8 -3 16 105
use FILL  FILL_405
timestamp 1713400504
transform 1 0 744 0 -1 2770
box -8 -3 16 105
use FILL  FILL_406
timestamp 1713400504
transform 1 0 736 0 -1 2770
box -8 -3 16 105
use FILL  FILL_407
timestamp 1713400504
transform 1 0 648 0 -1 2770
box -8 -3 16 105
use FILL  FILL_408
timestamp 1713400504
transform 1 0 640 0 -1 2770
box -8 -3 16 105
use FILL  FILL_409
timestamp 1713400504
transform 1 0 632 0 -1 2770
box -8 -3 16 105
use FILL  FILL_410
timestamp 1713400504
transform 1 0 608 0 -1 2770
box -8 -3 16 105
use FILL  FILL_411
timestamp 1713400504
transform 1 0 576 0 -1 2770
box -8 -3 16 105
use FILL  FILL_412
timestamp 1713400504
transform 1 0 568 0 -1 2770
box -8 -3 16 105
use FILL  FILL_413
timestamp 1713400504
transform 1 0 456 0 -1 2770
box -8 -3 16 105
use FILL  FILL_414
timestamp 1713400504
transform 1 0 448 0 -1 2770
box -8 -3 16 105
use FILL  FILL_415
timestamp 1713400504
transform 1 0 440 0 -1 2770
box -8 -3 16 105
use FILL  FILL_416
timestamp 1713400504
transform 1 0 432 0 -1 2770
box -8 -3 16 105
use FILL  FILL_417
timestamp 1713400504
transform 1 0 344 0 -1 2770
box -8 -3 16 105
use FILL  FILL_418
timestamp 1713400504
transform 1 0 336 0 -1 2770
box -8 -3 16 105
use FILL  FILL_419
timestamp 1713400504
transform 1 0 312 0 -1 2770
box -8 -3 16 105
use FILL  FILL_420
timestamp 1713400504
transform 1 0 256 0 -1 2770
box -8 -3 16 105
use FILL  FILL_421
timestamp 1713400504
transform 1 0 248 0 -1 2770
box -8 -3 16 105
use FILL  FILL_422
timestamp 1713400504
transform 1 0 240 0 -1 2770
box -8 -3 16 105
use FILL  FILL_423
timestamp 1713400504
transform 1 0 136 0 -1 2770
box -8 -3 16 105
use FILL  FILL_424
timestamp 1713400504
transform 1 0 128 0 -1 2770
box -8 -3 16 105
use FILL  FILL_425
timestamp 1713400504
transform 1 0 72 0 -1 2770
box -8 -3 16 105
use FILL  FILL_426
timestamp 1713400504
transform 1 0 2912 0 1 2570
box -8 -3 16 105
use FILL  FILL_427
timestamp 1713400504
transform 1 0 2904 0 1 2570
box -8 -3 16 105
use FILL  FILL_428
timestamp 1713400504
transform 1 0 2880 0 1 2570
box -8 -3 16 105
use FILL  FILL_429
timestamp 1713400504
transform 1 0 2872 0 1 2570
box -8 -3 16 105
use FILL  FILL_430
timestamp 1713400504
transform 1 0 2864 0 1 2570
box -8 -3 16 105
use FILL  FILL_431
timestamp 1713400504
transform 1 0 2816 0 1 2570
box -8 -3 16 105
use FILL  FILL_432
timestamp 1713400504
transform 1 0 2808 0 1 2570
box -8 -3 16 105
use FILL  FILL_433
timestamp 1713400504
transform 1 0 2800 0 1 2570
box -8 -3 16 105
use FILL  FILL_434
timestamp 1713400504
transform 1 0 2792 0 1 2570
box -8 -3 16 105
use FILL  FILL_435
timestamp 1713400504
transform 1 0 2784 0 1 2570
box -8 -3 16 105
use FILL  FILL_436
timestamp 1713400504
transform 1 0 2744 0 1 2570
box -8 -3 16 105
use FILL  FILL_437
timestamp 1713400504
transform 1 0 2736 0 1 2570
box -8 -3 16 105
use FILL  FILL_438
timestamp 1713400504
transform 1 0 2728 0 1 2570
box -8 -3 16 105
use FILL  FILL_439
timestamp 1713400504
transform 1 0 2688 0 1 2570
box -8 -3 16 105
use FILL  FILL_440
timestamp 1713400504
transform 1 0 2680 0 1 2570
box -8 -3 16 105
use FILL  FILL_441
timestamp 1713400504
transform 1 0 2672 0 1 2570
box -8 -3 16 105
use FILL  FILL_442
timestamp 1713400504
transform 1 0 2664 0 1 2570
box -8 -3 16 105
use FILL  FILL_443
timestamp 1713400504
transform 1 0 2656 0 1 2570
box -8 -3 16 105
use FILL  FILL_444
timestamp 1713400504
transform 1 0 2648 0 1 2570
box -8 -3 16 105
use FILL  FILL_445
timestamp 1713400504
transform 1 0 2600 0 1 2570
box -8 -3 16 105
use FILL  FILL_446
timestamp 1713400504
transform 1 0 2592 0 1 2570
box -8 -3 16 105
use FILL  FILL_447
timestamp 1713400504
transform 1 0 2584 0 1 2570
box -8 -3 16 105
use FILL  FILL_448
timestamp 1713400504
transform 1 0 2576 0 1 2570
box -8 -3 16 105
use FILL  FILL_449
timestamp 1713400504
transform 1 0 2568 0 1 2570
box -8 -3 16 105
use FILL  FILL_450
timestamp 1713400504
transform 1 0 2520 0 1 2570
box -8 -3 16 105
use FILL  FILL_451
timestamp 1713400504
transform 1 0 2512 0 1 2570
box -8 -3 16 105
use FILL  FILL_452
timestamp 1713400504
transform 1 0 2504 0 1 2570
box -8 -3 16 105
use FILL  FILL_453
timestamp 1713400504
transform 1 0 2496 0 1 2570
box -8 -3 16 105
use FILL  FILL_454
timestamp 1713400504
transform 1 0 2392 0 1 2570
box -8 -3 16 105
use FILL  FILL_455
timestamp 1713400504
transform 1 0 2384 0 1 2570
box -8 -3 16 105
use FILL  FILL_456
timestamp 1713400504
transform 1 0 2344 0 1 2570
box -8 -3 16 105
use FILL  FILL_457
timestamp 1713400504
transform 1 0 2336 0 1 2570
box -8 -3 16 105
use FILL  FILL_458
timestamp 1713400504
transform 1 0 2328 0 1 2570
box -8 -3 16 105
use FILL  FILL_459
timestamp 1713400504
transform 1 0 2320 0 1 2570
box -8 -3 16 105
use FILL  FILL_460
timestamp 1713400504
transform 1 0 2288 0 1 2570
box -8 -3 16 105
use FILL  FILL_461
timestamp 1713400504
transform 1 0 2280 0 1 2570
box -8 -3 16 105
use FILL  FILL_462
timestamp 1713400504
transform 1 0 2272 0 1 2570
box -8 -3 16 105
use FILL  FILL_463
timestamp 1713400504
transform 1 0 2240 0 1 2570
box -8 -3 16 105
use FILL  FILL_464
timestamp 1713400504
transform 1 0 2232 0 1 2570
box -8 -3 16 105
use FILL  FILL_465
timestamp 1713400504
transform 1 0 2224 0 1 2570
box -8 -3 16 105
use FILL  FILL_466
timestamp 1713400504
transform 1 0 2216 0 1 2570
box -8 -3 16 105
use FILL  FILL_467
timestamp 1713400504
transform 1 0 2184 0 1 2570
box -8 -3 16 105
use FILL  FILL_468
timestamp 1713400504
transform 1 0 2176 0 1 2570
box -8 -3 16 105
use FILL  FILL_469
timestamp 1713400504
transform 1 0 2152 0 1 2570
box -8 -3 16 105
use FILL  FILL_470
timestamp 1713400504
transform 1 0 2144 0 1 2570
box -8 -3 16 105
use FILL  FILL_471
timestamp 1713400504
transform 1 0 2136 0 1 2570
box -8 -3 16 105
use FILL  FILL_472
timestamp 1713400504
transform 1 0 2128 0 1 2570
box -8 -3 16 105
use FILL  FILL_473
timestamp 1713400504
transform 1 0 2096 0 1 2570
box -8 -3 16 105
use FILL  FILL_474
timestamp 1713400504
transform 1 0 2088 0 1 2570
box -8 -3 16 105
use FILL  FILL_475
timestamp 1713400504
transform 1 0 2080 0 1 2570
box -8 -3 16 105
use FILL  FILL_476
timestamp 1713400504
transform 1 0 2040 0 1 2570
box -8 -3 16 105
use FILL  FILL_477
timestamp 1713400504
transform 1 0 2032 0 1 2570
box -8 -3 16 105
use FILL  FILL_478
timestamp 1713400504
transform 1 0 2024 0 1 2570
box -8 -3 16 105
use FILL  FILL_479
timestamp 1713400504
transform 1 0 2016 0 1 2570
box -8 -3 16 105
use FILL  FILL_480
timestamp 1713400504
transform 1 0 2008 0 1 2570
box -8 -3 16 105
use FILL  FILL_481
timestamp 1713400504
transform 1 0 2000 0 1 2570
box -8 -3 16 105
use FILL  FILL_482
timestamp 1713400504
transform 1 0 1960 0 1 2570
box -8 -3 16 105
use FILL  FILL_483
timestamp 1713400504
transform 1 0 1952 0 1 2570
box -8 -3 16 105
use FILL  FILL_484
timestamp 1713400504
transform 1 0 1944 0 1 2570
box -8 -3 16 105
use FILL  FILL_485
timestamp 1713400504
transform 1 0 1912 0 1 2570
box -8 -3 16 105
use FILL  FILL_486
timestamp 1713400504
transform 1 0 1904 0 1 2570
box -8 -3 16 105
use FILL  FILL_487
timestamp 1713400504
transform 1 0 1896 0 1 2570
box -8 -3 16 105
use FILL  FILL_488
timestamp 1713400504
transform 1 0 1864 0 1 2570
box -8 -3 16 105
use FILL  FILL_489
timestamp 1713400504
transform 1 0 1856 0 1 2570
box -8 -3 16 105
use FILL  FILL_490
timestamp 1713400504
transform 1 0 1832 0 1 2570
box -8 -3 16 105
use FILL  FILL_491
timestamp 1713400504
transform 1 0 1824 0 1 2570
box -8 -3 16 105
use FILL  FILL_492
timestamp 1713400504
transform 1 0 1816 0 1 2570
box -8 -3 16 105
use FILL  FILL_493
timestamp 1713400504
transform 1 0 1808 0 1 2570
box -8 -3 16 105
use FILL  FILL_494
timestamp 1713400504
transform 1 0 1776 0 1 2570
box -8 -3 16 105
use FILL  FILL_495
timestamp 1713400504
transform 1 0 1768 0 1 2570
box -8 -3 16 105
use FILL  FILL_496
timestamp 1713400504
transform 1 0 1760 0 1 2570
box -8 -3 16 105
use FILL  FILL_497
timestamp 1713400504
transform 1 0 1720 0 1 2570
box -8 -3 16 105
use FILL  FILL_498
timestamp 1713400504
transform 1 0 1712 0 1 2570
box -8 -3 16 105
use FILL  FILL_499
timestamp 1713400504
transform 1 0 1704 0 1 2570
box -8 -3 16 105
use FILL  FILL_500
timestamp 1713400504
transform 1 0 1600 0 1 2570
box -8 -3 16 105
use FILL  FILL_501
timestamp 1713400504
transform 1 0 1560 0 1 2570
box -8 -3 16 105
use FILL  FILL_502
timestamp 1713400504
transform 1 0 1552 0 1 2570
box -8 -3 16 105
use FILL  FILL_503
timestamp 1713400504
transform 1 0 1448 0 1 2570
box -8 -3 16 105
use FILL  FILL_504
timestamp 1713400504
transform 1 0 1440 0 1 2570
box -8 -3 16 105
use FILL  FILL_505
timestamp 1713400504
transform 1 0 1432 0 1 2570
box -8 -3 16 105
use FILL  FILL_506
timestamp 1713400504
transform 1 0 1392 0 1 2570
box -8 -3 16 105
use FILL  FILL_507
timestamp 1713400504
transform 1 0 1384 0 1 2570
box -8 -3 16 105
use FILL  FILL_508
timestamp 1713400504
transform 1 0 1280 0 1 2570
box -8 -3 16 105
use FILL  FILL_509
timestamp 1713400504
transform 1 0 1272 0 1 2570
box -8 -3 16 105
use FILL  FILL_510
timestamp 1713400504
transform 1 0 1264 0 1 2570
box -8 -3 16 105
use FILL  FILL_511
timestamp 1713400504
transform 1 0 1256 0 1 2570
box -8 -3 16 105
use FILL  FILL_512
timestamp 1713400504
transform 1 0 1208 0 1 2570
box -8 -3 16 105
use FILL  FILL_513
timestamp 1713400504
transform 1 0 1200 0 1 2570
box -8 -3 16 105
use FILL  FILL_514
timestamp 1713400504
transform 1 0 1192 0 1 2570
box -8 -3 16 105
use FILL  FILL_515
timestamp 1713400504
transform 1 0 1184 0 1 2570
box -8 -3 16 105
use FILL  FILL_516
timestamp 1713400504
transform 1 0 1160 0 1 2570
box -8 -3 16 105
use FILL  FILL_517
timestamp 1713400504
transform 1 0 1152 0 1 2570
box -8 -3 16 105
use FILL  FILL_518
timestamp 1713400504
transform 1 0 1048 0 1 2570
box -8 -3 16 105
use FILL  FILL_519
timestamp 1713400504
transform 1 0 968 0 1 2570
box -8 -3 16 105
use FILL  FILL_520
timestamp 1713400504
transform 1 0 960 0 1 2570
box -8 -3 16 105
use FILL  FILL_521
timestamp 1713400504
transform 1 0 952 0 1 2570
box -8 -3 16 105
use FILL  FILL_522
timestamp 1713400504
transform 1 0 944 0 1 2570
box -8 -3 16 105
use FILL  FILL_523
timestamp 1713400504
transform 1 0 912 0 1 2570
box -8 -3 16 105
use FILL  FILL_524
timestamp 1713400504
transform 1 0 904 0 1 2570
box -8 -3 16 105
use FILL  FILL_525
timestamp 1713400504
transform 1 0 896 0 1 2570
box -8 -3 16 105
use FILL  FILL_526
timestamp 1713400504
transform 1 0 888 0 1 2570
box -8 -3 16 105
use FILL  FILL_527
timestamp 1713400504
transform 1 0 848 0 1 2570
box -8 -3 16 105
use FILL  FILL_528
timestamp 1713400504
transform 1 0 784 0 1 2570
box -8 -3 16 105
use FILL  FILL_529
timestamp 1713400504
transform 1 0 776 0 1 2570
box -8 -3 16 105
use FILL  FILL_530
timestamp 1713400504
transform 1 0 736 0 1 2570
box -8 -3 16 105
use FILL  FILL_531
timestamp 1713400504
transform 1 0 672 0 1 2570
box -8 -3 16 105
use FILL  FILL_532
timestamp 1713400504
transform 1 0 664 0 1 2570
box -8 -3 16 105
use FILL  FILL_533
timestamp 1713400504
transform 1 0 608 0 1 2570
box -8 -3 16 105
use FILL  FILL_534
timestamp 1713400504
transform 1 0 600 0 1 2570
box -8 -3 16 105
use FILL  FILL_535
timestamp 1713400504
transform 1 0 576 0 1 2570
box -8 -3 16 105
use FILL  FILL_536
timestamp 1713400504
transform 1 0 568 0 1 2570
box -8 -3 16 105
use FILL  FILL_537
timestamp 1713400504
transform 1 0 560 0 1 2570
box -8 -3 16 105
use FILL  FILL_538
timestamp 1713400504
transform 1 0 552 0 1 2570
box -8 -3 16 105
use FILL  FILL_539
timestamp 1713400504
transform 1 0 528 0 1 2570
box -8 -3 16 105
use FILL  FILL_540
timestamp 1713400504
transform 1 0 520 0 1 2570
box -8 -3 16 105
use FILL  FILL_541
timestamp 1713400504
transform 1 0 464 0 1 2570
box -8 -3 16 105
use FILL  FILL_542
timestamp 1713400504
transform 1 0 456 0 1 2570
box -8 -3 16 105
use FILL  FILL_543
timestamp 1713400504
transform 1 0 448 0 1 2570
box -8 -3 16 105
use FILL  FILL_544
timestamp 1713400504
transform 1 0 440 0 1 2570
box -8 -3 16 105
use FILL  FILL_545
timestamp 1713400504
transform 1 0 432 0 1 2570
box -8 -3 16 105
use FILL  FILL_546
timestamp 1713400504
transform 1 0 408 0 1 2570
box -8 -3 16 105
use FILL  FILL_547
timestamp 1713400504
transform 1 0 376 0 1 2570
box -8 -3 16 105
use FILL  FILL_548
timestamp 1713400504
transform 1 0 368 0 1 2570
box -8 -3 16 105
use FILL  FILL_549
timestamp 1713400504
transform 1 0 360 0 1 2570
box -8 -3 16 105
use FILL  FILL_550
timestamp 1713400504
transform 1 0 296 0 1 2570
box -8 -3 16 105
use FILL  FILL_551
timestamp 1713400504
transform 1 0 288 0 1 2570
box -8 -3 16 105
use FILL  FILL_552
timestamp 1713400504
transform 1 0 232 0 1 2570
box -8 -3 16 105
use FILL  FILL_553
timestamp 1713400504
transform 1 0 224 0 1 2570
box -8 -3 16 105
use FILL  FILL_554
timestamp 1713400504
transform 1 0 216 0 1 2570
box -8 -3 16 105
use FILL  FILL_555
timestamp 1713400504
transform 1 0 208 0 1 2570
box -8 -3 16 105
use FILL  FILL_556
timestamp 1713400504
transform 1 0 176 0 1 2570
box -8 -3 16 105
use FILL  FILL_557
timestamp 1713400504
transform 1 0 168 0 1 2570
box -8 -3 16 105
use FILL  FILL_558
timestamp 1713400504
transform 1 0 104 0 1 2570
box -8 -3 16 105
use FILL  FILL_559
timestamp 1713400504
transform 1 0 96 0 1 2570
box -8 -3 16 105
use FILL  FILL_560
timestamp 1713400504
transform 1 0 72 0 1 2570
box -8 -3 16 105
use FILL  FILL_561
timestamp 1713400504
transform 1 0 3008 0 -1 2570
box -8 -3 16 105
use FILL  FILL_562
timestamp 1713400504
transform 1 0 3000 0 -1 2570
box -8 -3 16 105
use FILL  FILL_563
timestamp 1713400504
transform 1 0 2992 0 -1 2570
box -8 -3 16 105
use FILL  FILL_564
timestamp 1713400504
transform 1 0 2984 0 -1 2570
box -8 -3 16 105
use FILL  FILL_565
timestamp 1713400504
transform 1 0 2936 0 -1 2570
box -8 -3 16 105
use FILL  FILL_566
timestamp 1713400504
transform 1 0 2928 0 -1 2570
box -8 -3 16 105
use FILL  FILL_567
timestamp 1713400504
transform 1 0 2920 0 -1 2570
box -8 -3 16 105
use FILL  FILL_568
timestamp 1713400504
transform 1 0 2912 0 -1 2570
box -8 -3 16 105
use FILL  FILL_569
timestamp 1713400504
transform 1 0 2904 0 -1 2570
box -8 -3 16 105
use FILL  FILL_570
timestamp 1713400504
transform 1 0 2896 0 -1 2570
box -8 -3 16 105
use FILL  FILL_571
timestamp 1713400504
transform 1 0 2888 0 -1 2570
box -8 -3 16 105
use FILL  FILL_572
timestamp 1713400504
transform 1 0 2840 0 -1 2570
box -8 -3 16 105
use FILL  FILL_573
timestamp 1713400504
transform 1 0 2832 0 -1 2570
box -8 -3 16 105
use FILL  FILL_574
timestamp 1713400504
transform 1 0 2824 0 -1 2570
box -8 -3 16 105
use FILL  FILL_575
timestamp 1713400504
transform 1 0 2816 0 -1 2570
box -8 -3 16 105
use FILL  FILL_576
timestamp 1713400504
transform 1 0 2712 0 -1 2570
box -8 -3 16 105
use FILL  FILL_577
timestamp 1713400504
transform 1 0 2704 0 -1 2570
box -8 -3 16 105
use FILL  FILL_578
timestamp 1713400504
transform 1 0 2696 0 -1 2570
box -8 -3 16 105
use FILL  FILL_579
timestamp 1713400504
transform 1 0 2688 0 -1 2570
box -8 -3 16 105
use FILL  FILL_580
timestamp 1713400504
transform 1 0 2648 0 -1 2570
box -8 -3 16 105
use FILL  FILL_581
timestamp 1713400504
transform 1 0 2640 0 -1 2570
box -8 -3 16 105
use FILL  FILL_582
timestamp 1713400504
transform 1 0 2632 0 -1 2570
box -8 -3 16 105
use FILL  FILL_583
timestamp 1713400504
transform 1 0 2624 0 -1 2570
box -8 -3 16 105
use FILL  FILL_584
timestamp 1713400504
transform 1 0 2592 0 -1 2570
box -8 -3 16 105
use FILL  FILL_585
timestamp 1713400504
transform 1 0 2584 0 -1 2570
box -8 -3 16 105
use FILL  FILL_586
timestamp 1713400504
transform 1 0 2576 0 -1 2570
box -8 -3 16 105
use FILL  FILL_587
timestamp 1713400504
transform 1 0 2568 0 -1 2570
box -8 -3 16 105
use FILL  FILL_588
timestamp 1713400504
transform 1 0 2560 0 -1 2570
box -8 -3 16 105
use FILL  FILL_589
timestamp 1713400504
transform 1 0 2528 0 -1 2570
box -8 -3 16 105
use FILL  FILL_590
timestamp 1713400504
transform 1 0 2520 0 -1 2570
box -8 -3 16 105
use FILL  FILL_591
timestamp 1713400504
transform 1 0 2488 0 -1 2570
box -8 -3 16 105
use FILL  FILL_592
timestamp 1713400504
transform 1 0 2480 0 -1 2570
box -8 -3 16 105
use FILL  FILL_593
timestamp 1713400504
transform 1 0 2472 0 -1 2570
box -8 -3 16 105
use FILL  FILL_594
timestamp 1713400504
transform 1 0 2464 0 -1 2570
box -8 -3 16 105
use FILL  FILL_595
timestamp 1713400504
transform 1 0 2456 0 -1 2570
box -8 -3 16 105
use FILL  FILL_596
timestamp 1713400504
transform 1 0 2416 0 -1 2570
box -8 -3 16 105
use FILL  FILL_597
timestamp 1713400504
transform 1 0 2408 0 -1 2570
box -8 -3 16 105
use FILL  FILL_598
timestamp 1713400504
transform 1 0 2400 0 -1 2570
box -8 -3 16 105
use FILL  FILL_599
timestamp 1713400504
transform 1 0 2392 0 -1 2570
box -8 -3 16 105
use FILL  FILL_600
timestamp 1713400504
transform 1 0 2360 0 -1 2570
box -8 -3 16 105
use FILL  FILL_601
timestamp 1713400504
transform 1 0 2352 0 -1 2570
box -8 -3 16 105
use FILL  FILL_602
timestamp 1713400504
transform 1 0 2344 0 -1 2570
box -8 -3 16 105
use FILL  FILL_603
timestamp 1713400504
transform 1 0 2312 0 -1 2570
box -8 -3 16 105
use FILL  FILL_604
timestamp 1713400504
transform 1 0 2304 0 -1 2570
box -8 -3 16 105
use FILL  FILL_605
timestamp 1713400504
transform 1 0 2296 0 -1 2570
box -8 -3 16 105
use FILL  FILL_606
timestamp 1713400504
transform 1 0 2288 0 -1 2570
box -8 -3 16 105
use FILL  FILL_607
timestamp 1713400504
transform 1 0 2256 0 -1 2570
box -8 -3 16 105
use FILL  FILL_608
timestamp 1713400504
transform 1 0 2248 0 -1 2570
box -8 -3 16 105
use FILL  FILL_609
timestamp 1713400504
transform 1 0 2240 0 -1 2570
box -8 -3 16 105
use FILL  FILL_610
timestamp 1713400504
transform 1 0 2208 0 -1 2570
box -8 -3 16 105
use FILL  FILL_611
timestamp 1713400504
transform 1 0 2200 0 -1 2570
box -8 -3 16 105
use FILL  FILL_612
timestamp 1713400504
transform 1 0 2192 0 -1 2570
box -8 -3 16 105
use FILL  FILL_613
timestamp 1713400504
transform 1 0 2184 0 -1 2570
box -8 -3 16 105
use FILL  FILL_614
timestamp 1713400504
transform 1 0 2152 0 -1 2570
box -8 -3 16 105
use FILL  FILL_615
timestamp 1713400504
transform 1 0 2144 0 -1 2570
box -8 -3 16 105
use FILL  FILL_616
timestamp 1713400504
transform 1 0 2136 0 -1 2570
box -8 -3 16 105
use FILL  FILL_617
timestamp 1713400504
transform 1 0 2128 0 -1 2570
box -8 -3 16 105
use FILL  FILL_618
timestamp 1713400504
transform 1 0 2096 0 -1 2570
box -8 -3 16 105
use FILL  FILL_619
timestamp 1713400504
transform 1 0 2088 0 -1 2570
box -8 -3 16 105
use FILL  FILL_620
timestamp 1713400504
transform 1 0 2080 0 -1 2570
box -8 -3 16 105
use FILL  FILL_621
timestamp 1713400504
transform 1 0 2048 0 -1 2570
box -8 -3 16 105
use FILL  FILL_622
timestamp 1713400504
transform 1 0 2040 0 -1 2570
box -8 -3 16 105
use FILL  FILL_623
timestamp 1713400504
transform 1 0 2032 0 -1 2570
box -8 -3 16 105
use FILL  FILL_624
timestamp 1713400504
transform 1 0 2024 0 -1 2570
box -8 -3 16 105
use FILL  FILL_625
timestamp 1713400504
transform 1 0 1992 0 -1 2570
box -8 -3 16 105
use FILL  FILL_626
timestamp 1713400504
transform 1 0 1984 0 -1 2570
box -8 -3 16 105
use FILL  FILL_627
timestamp 1713400504
transform 1 0 1976 0 -1 2570
box -8 -3 16 105
use FILL  FILL_628
timestamp 1713400504
transform 1 0 1968 0 -1 2570
box -8 -3 16 105
use FILL  FILL_629
timestamp 1713400504
transform 1 0 1936 0 -1 2570
box -8 -3 16 105
use FILL  FILL_630
timestamp 1713400504
transform 1 0 1928 0 -1 2570
box -8 -3 16 105
use FILL  FILL_631
timestamp 1713400504
transform 1 0 1896 0 -1 2570
box -8 -3 16 105
use FILL  FILL_632
timestamp 1713400504
transform 1 0 1888 0 -1 2570
box -8 -3 16 105
use FILL  FILL_633
timestamp 1713400504
transform 1 0 1880 0 -1 2570
box -8 -3 16 105
use FILL  FILL_634
timestamp 1713400504
transform 1 0 1872 0 -1 2570
box -8 -3 16 105
use FILL  FILL_635
timestamp 1713400504
transform 1 0 1864 0 -1 2570
box -8 -3 16 105
use FILL  FILL_636
timestamp 1713400504
transform 1 0 1808 0 -1 2570
box -8 -3 16 105
use FILL  FILL_637
timestamp 1713400504
transform 1 0 1800 0 -1 2570
box -8 -3 16 105
use FILL  FILL_638
timestamp 1713400504
transform 1 0 1792 0 -1 2570
box -8 -3 16 105
use FILL  FILL_639
timestamp 1713400504
transform 1 0 1784 0 -1 2570
box -8 -3 16 105
use FILL  FILL_640
timestamp 1713400504
transform 1 0 1776 0 -1 2570
box -8 -3 16 105
use FILL  FILL_641
timestamp 1713400504
transform 1 0 1768 0 -1 2570
box -8 -3 16 105
use FILL  FILL_642
timestamp 1713400504
transform 1 0 1720 0 -1 2570
box -8 -3 16 105
use FILL  FILL_643
timestamp 1713400504
transform 1 0 1712 0 -1 2570
box -8 -3 16 105
use FILL  FILL_644
timestamp 1713400504
transform 1 0 1704 0 -1 2570
box -8 -3 16 105
use FILL  FILL_645
timestamp 1713400504
transform 1 0 1696 0 -1 2570
box -8 -3 16 105
use FILL  FILL_646
timestamp 1713400504
transform 1 0 1688 0 -1 2570
box -8 -3 16 105
use FILL  FILL_647
timestamp 1713400504
transform 1 0 1680 0 -1 2570
box -8 -3 16 105
use FILL  FILL_648
timestamp 1713400504
transform 1 0 1656 0 -1 2570
box -8 -3 16 105
use FILL  FILL_649
timestamp 1713400504
transform 1 0 1616 0 -1 2570
box -8 -3 16 105
use FILL  FILL_650
timestamp 1713400504
transform 1 0 1608 0 -1 2570
box -8 -3 16 105
use FILL  FILL_651
timestamp 1713400504
transform 1 0 1600 0 -1 2570
box -8 -3 16 105
use FILL  FILL_652
timestamp 1713400504
transform 1 0 1496 0 -1 2570
box -8 -3 16 105
use FILL  FILL_653
timestamp 1713400504
transform 1 0 1472 0 -1 2570
box -8 -3 16 105
use FILL  FILL_654
timestamp 1713400504
transform 1 0 1464 0 -1 2570
box -8 -3 16 105
use FILL  FILL_655
timestamp 1713400504
transform 1 0 1456 0 -1 2570
box -8 -3 16 105
use FILL  FILL_656
timestamp 1713400504
transform 1 0 1448 0 -1 2570
box -8 -3 16 105
use FILL  FILL_657
timestamp 1713400504
transform 1 0 1400 0 -1 2570
box -8 -3 16 105
use FILL  FILL_658
timestamp 1713400504
transform 1 0 1392 0 -1 2570
box -8 -3 16 105
use FILL  FILL_659
timestamp 1713400504
transform 1 0 1384 0 -1 2570
box -8 -3 16 105
use FILL  FILL_660
timestamp 1713400504
transform 1 0 1376 0 -1 2570
box -8 -3 16 105
use FILL  FILL_661
timestamp 1713400504
transform 1 0 1368 0 -1 2570
box -8 -3 16 105
use FILL  FILL_662
timestamp 1713400504
transform 1 0 1344 0 -1 2570
box -8 -3 16 105
use FILL  FILL_663
timestamp 1713400504
transform 1 0 1336 0 -1 2570
box -8 -3 16 105
use FILL  FILL_664
timestamp 1713400504
transform 1 0 1328 0 -1 2570
box -8 -3 16 105
use FILL  FILL_665
timestamp 1713400504
transform 1 0 1320 0 -1 2570
box -8 -3 16 105
use FILL  FILL_666
timestamp 1713400504
transform 1 0 1272 0 -1 2570
box -8 -3 16 105
use FILL  FILL_667
timestamp 1713400504
transform 1 0 1264 0 -1 2570
box -8 -3 16 105
use FILL  FILL_668
timestamp 1713400504
transform 1 0 1256 0 -1 2570
box -8 -3 16 105
use FILL  FILL_669
timestamp 1713400504
transform 1 0 1152 0 -1 2570
box -8 -3 16 105
use FILL  FILL_670
timestamp 1713400504
transform 1 0 1144 0 -1 2570
box -8 -3 16 105
use FILL  FILL_671
timestamp 1713400504
transform 1 0 1136 0 -1 2570
box -8 -3 16 105
use FILL  FILL_672
timestamp 1713400504
transform 1 0 1128 0 -1 2570
box -8 -3 16 105
use FILL  FILL_673
timestamp 1713400504
transform 1 0 1080 0 -1 2570
box -8 -3 16 105
use FILL  FILL_674
timestamp 1713400504
transform 1 0 1072 0 -1 2570
box -8 -3 16 105
use FILL  FILL_675
timestamp 1713400504
transform 1 0 1064 0 -1 2570
box -8 -3 16 105
use FILL  FILL_676
timestamp 1713400504
transform 1 0 1056 0 -1 2570
box -8 -3 16 105
use FILL  FILL_677
timestamp 1713400504
transform 1 0 1048 0 -1 2570
box -8 -3 16 105
use FILL  FILL_678
timestamp 1713400504
transform 1 0 1040 0 -1 2570
box -8 -3 16 105
use FILL  FILL_679
timestamp 1713400504
transform 1 0 1032 0 -1 2570
box -8 -3 16 105
use FILL  FILL_680
timestamp 1713400504
transform 1 0 984 0 -1 2570
box -8 -3 16 105
use FILL  FILL_681
timestamp 1713400504
transform 1 0 976 0 -1 2570
box -8 -3 16 105
use FILL  FILL_682
timestamp 1713400504
transform 1 0 968 0 -1 2570
box -8 -3 16 105
use FILL  FILL_683
timestamp 1713400504
transform 1 0 960 0 -1 2570
box -8 -3 16 105
use FILL  FILL_684
timestamp 1713400504
transform 1 0 952 0 -1 2570
box -8 -3 16 105
use FILL  FILL_685
timestamp 1713400504
transform 1 0 944 0 -1 2570
box -8 -3 16 105
use FILL  FILL_686
timestamp 1713400504
transform 1 0 936 0 -1 2570
box -8 -3 16 105
use FILL  FILL_687
timestamp 1713400504
transform 1 0 904 0 -1 2570
box -8 -3 16 105
use FILL  FILL_688
timestamp 1713400504
transform 1 0 840 0 -1 2570
box -8 -3 16 105
use FILL  FILL_689
timestamp 1713400504
transform 1 0 832 0 -1 2570
box -8 -3 16 105
use FILL  FILL_690
timestamp 1713400504
transform 1 0 824 0 -1 2570
box -8 -3 16 105
use FILL  FILL_691
timestamp 1713400504
transform 1 0 696 0 -1 2570
box -8 -3 16 105
use FILL  FILL_692
timestamp 1713400504
transform 1 0 688 0 -1 2570
box -8 -3 16 105
use FILL  FILL_693
timestamp 1713400504
transform 1 0 680 0 -1 2570
box -8 -3 16 105
use FILL  FILL_694
timestamp 1713400504
transform 1 0 672 0 -1 2570
box -8 -3 16 105
use FILL  FILL_695
timestamp 1713400504
transform 1 0 632 0 -1 2570
box -8 -3 16 105
use FILL  FILL_696
timestamp 1713400504
transform 1 0 624 0 -1 2570
box -8 -3 16 105
use FILL  FILL_697
timestamp 1713400504
transform 1 0 560 0 -1 2570
box -8 -3 16 105
use FILL  FILL_698
timestamp 1713400504
transform 1 0 552 0 -1 2570
box -8 -3 16 105
use FILL  FILL_699
timestamp 1713400504
transform 1 0 544 0 -1 2570
box -8 -3 16 105
use FILL  FILL_700
timestamp 1713400504
transform 1 0 536 0 -1 2570
box -8 -3 16 105
use FILL  FILL_701
timestamp 1713400504
transform 1 0 496 0 -1 2570
box -8 -3 16 105
use FILL  FILL_702
timestamp 1713400504
transform 1 0 488 0 -1 2570
box -8 -3 16 105
use FILL  FILL_703
timestamp 1713400504
transform 1 0 424 0 -1 2570
box -8 -3 16 105
use FILL  FILL_704
timestamp 1713400504
transform 1 0 416 0 -1 2570
box -8 -3 16 105
use FILL  FILL_705
timestamp 1713400504
transform 1 0 408 0 -1 2570
box -8 -3 16 105
use FILL  FILL_706
timestamp 1713400504
transform 1 0 400 0 -1 2570
box -8 -3 16 105
use FILL  FILL_707
timestamp 1713400504
transform 1 0 392 0 -1 2570
box -8 -3 16 105
use FILL  FILL_708
timestamp 1713400504
transform 1 0 368 0 -1 2570
box -8 -3 16 105
use FILL  FILL_709
timestamp 1713400504
transform 1 0 360 0 -1 2570
box -8 -3 16 105
use FILL  FILL_710
timestamp 1713400504
transform 1 0 352 0 -1 2570
box -8 -3 16 105
use FILL  FILL_711
timestamp 1713400504
transform 1 0 296 0 -1 2570
box -8 -3 16 105
use FILL  FILL_712
timestamp 1713400504
transform 1 0 288 0 -1 2570
box -8 -3 16 105
use FILL  FILL_713
timestamp 1713400504
transform 1 0 280 0 -1 2570
box -8 -3 16 105
use FILL  FILL_714
timestamp 1713400504
transform 1 0 272 0 -1 2570
box -8 -3 16 105
use FILL  FILL_715
timestamp 1713400504
transform 1 0 264 0 -1 2570
box -8 -3 16 105
use FILL  FILL_716
timestamp 1713400504
transform 1 0 256 0 -1 2570
box -8 -3 16 105
use FILL  FILL_717
timestamp 1713400504
transform 1 0 232 0 -1 2570
box -8 -3 16 105
use FILL  FILL_718
timestamp 1713400504
transform 1 0 224 0 -1 2570
box -8 -3 16 105
use FILL  FILL_719
timestamp 1713400504
transform 1 0 216 0 -1 2570
box -8 -3 16 105
use FILL  FILL_720
timestamp 1713400504
transform 1 0 184 0 -1 2570
box -8 -3 16 105
use FILL  FILL_721
timestamp 1713400504
transform 1 0 176 0 -1 2570
box -8 -3 16 105
use FILL  FILL_722
timestamp 1713400504
transform 1 0 168 0 -1 2570
box -8 -3 16 105
use FILL  FILL_723
timestamp 1713400504
transform 1 0 160 0 -1 2570
box -8 -3 16 105
use FILL  FILL_724
timestamp 1713400504
transform 1 0 152 0 -1 2570
box -8 -3 16 105
use FILL  FILL_725
timestamp 1713400504
transform 1 0 144 0 -1 2570
box -8 -3 16 105
use FILL  FILL_726
timestamp 1713400504
transform 1 0 88 0 -1 2570
box -8 -3 16 105
use FILL  FILL_727
timestamp 1713400504
transform 1 0 80 0 -1 2570
box -8 -3 16 105
use FILL  FILL_728
timestamp 1713400504
transform 1 0 72 0 -1 2570
box -8 -3 16 105
use FILL  FILL_729
timestamp 1713400504
transform 1 0 3008 0 1 2370
box -8 -3 16 105
use FILL  FILL_730
timestamp 1713400504
transform 1 0 3000 0 1 2370
box -8 -3 16 105
use FILL  FILL_731
timestamp 1713400504
transform 1 0 2992 0 1 2370
box -8 -3 16 105
use FILL  FILL_732
timestamp 1713400504
transform 1 0 2952 0 1 2370
box -8 -3 16 105
use FILL  FILL_733
timestamp 1713400504
transform 1 0 2944 0 1 2370
box -8 -3 16 105
use FILL  FILL_734
timestamp 1713400504
transform 1 0 2936 0 1 2370
box -8 -3 16 105
use FILL  FILL_735
timestamp 1713400504
transform 1 0 2928 0 1 2370
box -8 -3 16 105
use FILL  FILL_736
timestamp 1713400504
transform 1 0 2920 0 1 2370
box -8 -3 16 105
use FILL  FILL_737
timestamp 1713400504
transform 1 0 2912 0 1 2370
box -8 -3 16 105
use FILL  FILL_738
timestamp 1713400504
transform 1 0 2872 0 1 2370
box -8 -3 16 105
use FILL  FILL_739
timestamp 1713400504
transform 1 0 2864 0 1 2370
box -8 -3 16 105
use FILL  FILL_740
timestamp 1713400504
transform 1 0 2856 0 1 2370
box -8 -3 16 105
use FILL  FILL_741
timestamp 1713400504
transform 1 0 2816 0 1 2370
box -8 -3 16 105
use FILL  FILL_742
timestamp 1713400504
transform 1 0 2808 0 1 2370
box -8 -3 16 105
use FILL  FILL_743
timestamp 1713400504
transform 1 0 2800 0 1 2370
box -8 -3 16 105
use FILL  FILL_744
timestamp 1713400504
transform 1 0 2792 0 1 2370
box -8 -3 16 105
use FILL  FILL_745
timestamp 1713400504
transform 1 0 2784 0 1 2370
box -8 -3 16 105
use FILL  FILL_746
timestamp 1713400504
transform 1 0 2752 0 1 2370
box -8 -3 16 105
use FILL  FILL_747
timestamp 1713400504
transform 1 0 2728 0 1 2370
box -8 -3 16 105
use FILL  FILL_748
timestamp 1713400504
transform 1 0 2720 0 1 2370
box -8 -3 16 105
use FILL  FILL_749
timestamp 1713400504
transform 1 0 2712 0 1 2370
box -8 -3 16 105
use FILL  FILL_750
timestamp 1713400504
transform 1 0 2704 0 1 2370
box -8 -3 16 105
use FILL  FILL_751
timestamp 1713400504
transform 1 0 2696 0 1 2370
box -8 -3 16 105
use FILL  FILL_752
timestamp 1713400504
transform 1 0 2688 0 1 2370
box -8 -3 16 105
use FILL  FILL_753
timestamp 1713400504
transform 1 0 2648 0 1 2370
box -8 -3 16 105
use FILL  FILL_754
timestamp 1713400504
transform 1 0 2640 0 1 2370
box -8 -3 16 105
use FILL  FILL_755
timestamp 1713400504
transform 1 0 2632 0 1 2370
box -8 -3 16 105
use FILL  FILL_756
timestamp 1713400504
transform 1 0 2624 0 1 2370
box -8 -3 16 105
use FILL  FILL_757
timestamp 1713400504
transform 1 0 2584 0 1 2370
box -8 -3 16 105
use FILL  FILL_758
timestamp 1713400504
transform 1 0 2576 0 1 2370
box -8 -3 16 105
use FILL  FILL_759
timestamp 1713400504
transform 1 0 2568 0 1 2370
box -8 -3 16 105
use FILL  FILL_760
timestamp 1713400504
transform 1 0 2560 0 1 2370
box -8 -3 16 105
use FILL  FILL_761
timestamp 1713400504
transform 1 0 2552 0 1 2370
box -8 -3 16 105
use FILL  FILL_762
timestamp 1713400504
transform 1 0 2512 0 1 2370
box -8 -3 16 105
use FILL  FILL_763
timestamp 1713400504
transform 1 0 2504 0 1 2370
box -8 -3 16 105
use FILL  FILL_764
timestamp 1713400504
transform 1 0 2496 0 1 2370
box -8 -3 16 105
use FILL  FILL_765
timestamp 1713400504
transform 1 0 2472 0 1 2370
box -8 -3 16 105
use FILL  FILL_766
timestamp 1713400504
transform 1 0 2464 0 1 2370
box -8 -3 16 105
use FILL  FILL_767
timestamp 1713400504
transform 1 0 2456 0 1 2370
box -8 -3 16 105
use FILL  FILL_768
timestamp 1713400504
transform 1 0 2448 0 1 2370
box -8 -3 16 105
use FILL  FILL_769
timestamp 1713400504
transform 1 0 2416 0 1 2370
box -8 -3 16 105
use FILL  FILL_770
timestamp 1713400504
transform 1 0 2408 0 1 2370
box -8 -3 16 105
use FILL  FILL_771
timestamp 1713400504
transform 1 0 2400 0 1 2370
box -8 -3 16 105
use FILL  FILL_772
timestamp 1713400504
transform 1 0 2392 0 1 2370
box -8 -3 16 105
use FILL  FILL_773
timestamp 1713400504
transform 1 0 2384 0 1 2370
box -8 -3 16 105
use FILL  FILL_774
timestamp 1713400504
transform 1 0 2352 0 1 2370
box -8 -3 16 105
use FILL  FILL_775
timestamp 1713400504
transform 1 0 2344 0 1 2370
box -8 -3 16 105
use FILL  FILL_776
timestamp 1713400504
transform 1 0 2336 0 1 2370
box -8 -3 16 105
use FILL  FILL_777
timestamp 1713400504
transform 1 0 2328 0 1 2370
box -8 -3 16 105
use FILL  FILL_778
timestamp 1713400504
transform 1 0 2320 0 1 2370
box -8 -3 16 105
use FILL  FILL_779
timestamp 1713400504
transform 1 0 2288 0 1 2370
box -8 -3 16 105
use FILL  FILL_780
timestamp 1713400504
transform 1 0 2280 0 1 2370
box -8 -3 16 105
use FILL  FILL_781
timestamp 1713400504
transform 1 0 2272 0 1 2370
box -8 -3 16 105
use FILL  FILL_782
timestamp 1713400504
transform 1 0 2264 0 1 2370
box -8 -3 16 105
use FILL  FILL_783
timestamp 1713400504
transform 1 0 2232 0 1 2370
box -8 -3 16 105
use FILL  FILL_784
timestamp 1713400504
transform 1 0 2224 0 1 2370
box -8 -3 16 105
use FILL  FILL_785
timestamp 1713400504
transform 1 0 2216 0 1 2370
box -8 -3 16 105
use FILL  FILL_786
timestamp 1713400504
transform 1 0 2208 0 1 2370
box -8 -3 16 105
use FILL  FILL_787
timestamp 1713400504
transform 1 0 2176 0 1 2370
box -8 -3 16 105
use FILL  FILL_788
timestamp 1713400504
transform 1 0 2168 0 1 2370
box -8 -3 16 105
use FILL  FILL_789
timestamp 1713400504
transform 1 0 2160 0 1 2370
box -8 -3 16 105
use FILL  FILL_790
timestamp 1713400504
transform 1 0 2152 0 1 2370
box -8 -3 16 105
use FILL  FILL_791
timestamp 1713400504
transform 1 0 2144 0 1 2370
box -8 -3 16 105
use FILL  FILL_792
timestamp 1713400504
transform 1 0 2136 0 1 2370
box -8 -3 16 105
use FILL  FILL_793
timestamp 1713400504
transform 1 0 2096 0 1 2370
box -8 -3 16 105
use FILL  FILL_794
timestamp 1713400504
transform 1 0 2088 0 1 2370
box -8 -3 16 105
use FILL  FILL_795
timestamp 1713400504
transform 1 0 2080 0 1 2370
box -8 -3 16 105
use FILL  FILL_796
timestamp 1713400504
transform 1 0 2072 0 1 2370
box -8 -3 16 105
use FILL  FILL_797
timestamp 1713400504
transform 1 0 2040 0 1 2370
box -8 -3 16 105
use FILL  FILL_798
timestamp 1713400504
transform 1 0 2032 0 1 2370
box -8 -3 16 105
use FILL  FILL_799
timestamp 1713400504
transform 1 0 2024 0 1 2370
box -8 -3 16 105
use FILL  FILL_800
timestamp 1713400504
transform 1 0 2016 0 1 2370
box -8 -3 16 105
use FILL  FILL_801
timestamp 1713400504
transform 1 0 1984 0 1 2370
box -8 -3 16 105
use FILL  FILL_802
timestamp 1713400504
transform 1 0 1976 0 1 2370
box -8 -3 16 105
use FILL  FILL_803
timestamp 1713400504
transform 1 0 1968 0 1 2370
box -8 -3 16 105
use FILL  FILL_804
timestamp 1713400504
transform 1 0 1960 0 1 2370
box -8 -3 16 105
use FILL  FILL_805
timestamp 1713400504
transform 1 0 1928 0 1 2370
box -8 -3 16 105
use FILL  FILL_806
timestamp 1713400504
transform 1 0 1920 0 1 2370
box -8 -3 16 105
use FILL  FILL_807
timestamp 1713400504
transform 1 0 1912 0 1 2370
box -8 -3 16 105
use FILL  FILL_808
timestamp 1713400504
transform 1 0 1904 0 1 2370
box -8 -3 16 105
use FILL  FILL_809
timestamp 1713400504
transform 1 0 1872 0 1 2370
box -8 -3 16 105
use FILL  FILL_810
timestamp 1713400504
transform 1 0 1864 0 1 2370
box -8 -3 16 105
use FILL  FILL_811
timestamp 1713400504
transform 1 0 1856 0 1 2370
box -8 -3 16 105
use FILL  FILL_812
timestamp 1713400504
transform 1 0 1848 0 1 2370
box -8 -3 16 105
use FILL  FILL_813
timestamp 1713400504
transform 1 0 1808 0 1 2370
box -8 -3 16 105
use FILL  FILL_814
timestamp 1713400504
transform 1 0 1800 0 1 2370
box -8 -3 16 105
use FILL  FILL_815
timestamp 1713400504
transform 1 0 1792 0 1 2370
box -8 -3 16 105
use FILL  FILL_816
timestamp 1713400504
transform 1 0 1688 0 1 2370
box -8 -3 16 105
use FILL  FILL_817
timestamp 1713400504
transform 1 0 1680 0 1 2370
box -8 -3 16 105
use FILL  FILL_818
timestamp 1713400504
transform 1 0 1672 0 1 2370
box -8 -3 16 105
use FILL  FILL_819
timestamp 1713400504
transform 1 0 1648 0 1 2370
box -8 -3 16 105
use FILL  FILL_820
timestamp 1713400504
transform 1 0 1640 0 1 2370
box -8 -3 16 105
use FILL  FILL_821
timestamp 1713400504
transform 1 0 1632 0 1 2370
box -8 -3 16 105
use FILL  FILL_822
timestamp 1713400504
transform 1 0 1592 0 1 2370
box -8 -3 16 105
use FILL  FILL_823
timestamp 1713400504
transform 1 0 1584 0 1 2370
box -8 -3 16 105
use FILL  FILL_824
timestamp 1713400504
transform 1 0 1576 0 1 2370
box -8 -3 16 105
use FILL  FILL_825
timestamp 1713400504
transform 1 0 1568 0 1 2370
box -8 -3 16 105
use FILL  FILL_826
timestamp 1713400504
transform 1 0 1560 0 1 2370
box -8 -3 16 105
use FILL  FILL_827
timestamp 1713400504
transform 1 0 1528 0 1 2370
box -8 -3 16 105
use FILL  FILL_828
timestamp 1713400504
transform 1 0 1520 0 1 2370
box -8 -3 16 105
use FILL  FILL_829
timestamp 1713400504
transform 1 0 1512 0 1 2370
box -8 -3 16 105
use FILL  FILL_830
timestamp 1713400504
transform 1 0 1504 0 1 2370
box -8 -3 16 105
use FILL  FILL_831
timestamp 1713400504
transform 1 0 1496 0 1 2370
box -8 -3 16 105
use FILL  FILL_832
timestamp 1713400504
transform 1 0 1488 0 1 2370
box -8 -3 16 105
use FILL  FILL_833
timestamp 1713400504
transform 1 0 1440 0 1 2370
box -8 -3 16 105
use FILL  FILL_834
timestamp 1713400504
transform 1 0 1432 0 1 2370
box -8 -3 16 105
use FILL  FILL_835
timestamp 1713400504
transform 1 0 1424 0 1 2370
box -8 -3 16 105
use FILL  FILL_836
timestamp 1713400504
transform 1 0 1416 0 1 2370
box -8 -3 16 105
use FILL  FILL_837
timestamp 1713400504
transform 1 0 1408 0 1 2370
box -8 -3 16 105
use FILL  FILL_838
timestamp 1713400504
transform 1 0 1400 0 1 2370
box -8 -3 16 105
use FILL  FILL_839
timestamp 1713400504
transform 1 0 1392 0 1 2370
box -8 -3 16 105
use FILL  FILL_840
timestamp 1713400504
transform 1 0 1344 0 1 2370
box -8 -3 16 105
use FILL  FILL_841
timestamp 1713400504
transform 1 0 1336 0 1 2370
box -8 -3 16 105
use FILL  FILL_842
timestamp 1713400504
transform 1 0 1328 0 1 2370
box -8 -3 16 105
use FILL  FILL_843
timestamp 1713400504
transform 1 0 1320 0 1 2370
box -8 -3 16 105
use FILL  FILL_844
timestamp 1713400504
transform 1 0 1312 0 1 2370
box -8 -3 16 105
use FILL  FILL_845
timestamp 1713400504
transform 1 0 1304 0 1 2370
box -8 -3 16 105
use FILL  FILL_846
timestamp 1713400504
transform 1 0 1296 0 1 2370
box -8 -3 16 105
use FILL  FILL_847
timestamp 1713400504
transform 1 0 1288 0 1 2370
box -8 -3 16 105
use FILL  FILL_848
timestamp 1713400504
transform 1 0 1248 0 1 2370
box -8 -3 16 105
use FILL  FILL_849
timestamp 1713400504
transform 1 0 1240 0 1 2370
box -8 -3 16 105
use FILL  FILL_850
timestamp 1713400504
transform 1 0 1232 0 1 2370
box -8 -3 16 105
use FILL  FILL_851
timestamp 1713400504
transform 1 0 1224 0 1 2370
box -8 -3 16 105
use FILL  FILL_852
timestamp 1713400504
transform 1 0 1216 0 1 2370
box -8 -3 16 105
use FILL  FILL_853
timestamp 1713400504
transform 1 0 1208 0 1 2370
box -8 -3 16 105
use FILL  FILL_854
timestamp 1713400504
transform 1 0 1200 0 1 2370
box -8 -3 16 105
use FILL  FILL_855
timestamp 1713400504
transform 1 0 1160 0 1 2370
box -8 -3 16 105
use FILL  FILL_856
timestamp 1713400504
transform 1 0 1152 0 1 2370
box -8 -3 16 105
use FILL  FILL_857
timestamp 1713400504
transform 1 0 1144 0 1 2370
box -8 -3 16 105
use FILL  FILL_858
timestamp 1713400504
transform 1 0 1136 0 1 2370
box -8 -3 16 105
use FILL  FILL_859
timestamp 1713400504
transform 1 0 1128 0 1 2370
box -8 -3 16 105
use FILL  FILL_860
timestamp 1713400504
transform 1 0 1120 0 1 2370
box -8 -3 16 105
use FILL  FILL_861
timestamp 1713400504
transform 1 0 1112 0 1 2370
box -8 -3 16 105
use FILL  FILL_862
timestamp 1713400504
transform 1 0 1104 0 1 2370
box -8 -3 16 105
use FILL  FILL_863
timestamp 1713400504
transform 1 0 1096 0 1 2370
box -8 -3 16 105
use FILL  FILL_864
timestamp 1713400504
transform 1 0 1056 0 1 2370
box -8 -3 16 105
use FILL  FILL_865
timestamp 1713400504
transform 1 0 1048 0 1 2370
box -8 -3 16 105
use FILL  FILL_866
timestamp 1713400504
transform 1 0 1040 0 1 2370
box -8 -3 16 105
use FILL  FILL_867
timestamp 1713400504
transform 1 0 1032 0 1 2370
box -8 -3 16 105
use FILL  FILL_868
timestamp 1713400504
transform 1 0 1024 0 1 2370
box -8 -3 16 105
use FILL  FILL_869
timestamp 1713400504
transform 1 0 1016 0 1 2370
box -8 -3 16 105
use FILL  FILL_870
timestamp 1713400504
transform 1 0 1008 0 1 2370
box -8 -3 16 105
use FILL  FILL_871
timestamp 1713400504
transform 1 0 1000 0 1 2370
box -8 -3 16 105
use FILL  FILL_872
timestamp 1713400504
transform 1 0 992 0 1 2370
box -8 -3 16 105
use FILL  FILL_873
timestamp 1713400504
transform 1 0 944 0 1 2370
box -8 -3 16 105
use FILL  FILL_874
timestamp 1713400504
transform 1 0 936 0 1 2370
box -8 -3 16 105
use FILL  FILL_875
timestamp 1713400504
transform 1 0 928 0 1 2370
box -8 -3 16 105
use FILL  FILL_876
timestamp 1713400504
transform 1 0 920 0 1 2370
box -8 -3 16 105
use FILL  FILL_877
timestamp 1713400504
transform 1 0 912 0 1 2370
box -8 -3 16 105
use FILL  FILL_878
timestamp 1713400504
transform 1 0 904 0 1 2370
box -8 -3 16 105
use FILL  FILL_879
timestamp 1713400504
transform 1 0 896 0 1 2370
box -8 -3 16 105
use FILL  FILL_880
timestamp 1713400504
transform 1 0 888 0 1 2370
box -8 -3 16 105
use FILL  FILL_881
timestamp 1713400504
transform 1 0 848 0 1 2370
box -8 -3 16 105
use FILL  FILL_882
timestamp 1713400504
transform 1 0 840 0 1 2370
box -8 -3 16 105
use FILL  FILL_883
timestamp 1713400504
transform 1 0 832 0 1 2370
box -8 -3 16 105
use FILL  FILL_884
timestamp 1713400504
transform 1 0 824 0 1 2370
box -8 -3 16 105
use FILL  FILL_885
timestamp 1713400504
transform 1 0 816 0 1 2370
box -8 -3 16 105
use FILL  FILL_886
timestamp 1713400504
transform 1 0 808 0 1 2370
box -8 -3 16 105
use FILL  FILL_887
timestamp 1713400504
transform 1 0 800 0 1 2370
box -8 -3 16 105
use FILL  FILL_888
timestamp 1713400504
transform 1 0 672 0 1 2370
box -8 -3 16 105
use FILL  FILL_889
timestamp 1713400504
transform 1 0 664 0 1 2370
box -8 -3 16 105
use FILL  FILL_890
timestamp 1713400504
transform 1 0 656 0 1 2370
box -8 -3 16 105
use FILL  FILL_891
timestamp 1713400504
transform 1 0 648 0 1 2370
box -8 -3 16 105
use FILL  FILL_892
timestamp 1713400504
transform 1 0 520 0 1 2370
box -8 -3 16 105
use FILL  FILL_893
timestamp 1713400504
transform 1 0 512 0 1 2370
box -8 -3 16 105
use FILL  FILL_894
timestamp 1713400504
transform 1 0 504 0 1 2370
box -8 -3 16 105
use FILL  FILL_895
timestamp 1713400504
transform 1 0 496 0 1 2370
box -8 -3 16 105
use FILL  FILL_896
timestamp 1713400504
transform 1 0 488 0 1 2370
box -8 -3 16 105
use FILL  FILL_897
timestamp 1713400504
transform 1 0 480 0 1 2370
box -8 -3 16 105
use FILL  FILL_898
timestamp 1713400504
transform 1 0 472 0 1 2370
box -8 -3 16 105
use FILL  FILL_899
timestamp 1713400504
transform 1 0 464 0 1 2370
box -8 -3 16 105
use FILL  FILL_900
timestamp 1713400504
transform 1 0 456 0 1 2370
box -8 -3 16 105
use FILL  FILL_901
timestamp 1713400504
transform 1 0 448 0 1 2370
box -8 -3 16 105
use FILL  FILL_902
timestamp 1713400504
transform 1 0 440 0 1 2370
box -8 -3 16 105
use FILL  FILL_903
timestamp 1713400504
transform 1 0 432 0 1 2370
box -8 -3 16 105
use FILL  FILL_904
timestamp 1713400504
transform 1 0 304 0 1 2370
box -8 -3 16 105
use FILL  FILL_905
timestamp 1713400504
transform 1 0 296 0 1 2370
box -8 -3 16 105
use FILL  FILL_906
timestamp 1713400504
transform 1 0 288 0 1 2370
box -8 -3 16 105
use FILL  FILL_907
timestamp 1713400504
transform 1 0 280 0 1 2370
box -8 -3 16 105
use FILL  FILL_908
timestamp 1713400504
transform 1 0 272 0 1 2370
box -8 -3 16 105
use FILL  FILL_909
timestamp 1713400504
transform 1 0 208 0 1 2370
box -8 -3 16 105
use FILL  FILL_910
timestamp 1713400504
transform 1 0 200 0 1 2370
box -8 -3 16 105
use FILL  FILL_911
timestamp 1713400504
transform 1 0 192 0 1 2370
box -8 -3 16 105
use FILL  FILL_912
timestamp 1713400504
transform 1 0 184 0 1 2370
box -8 -3 16 105
use FILL  FILL_913
timestamp 1713400504
transform 1 0 128 0 1 2370
box -8 -3 16 105
use FILL  FILL_914
timestamp 1713400504
transform 1 0 120 0 1 2370
box -8 -3 16 105
use FILL  FILL_915
timestamp 1713400504
transform 1 0 112 0 1 2370
box -8 -3 16 105
use FILL  FILL_916
timestamp 1713400504
transform 1 0 104 0 1 2370
box -8 -3 16 105
use FILL  FILL_917
timestamp 1713400504
transform 1 0 96 0 1 2370
box -8 -3 16 105
use FILL  FILL_918
timestamp 1713400504
transform 1 0 88 0 1 2370
box -8 -3 16 105
use FILL  FILL_919
timestamp 1713400504
transform 1 0 80 0 1 2370
box -8 -3 16 105
use FILL  FILL_920
timestamp 1713400504
transform 1 0 72 0 1 2370
box -8 -3 16 105
use FILL  FILL_921
timestamp 1713400504
transform 1 0 2896 0 -1 2370
box -8 -3 16 105
use FILL  FILL_922
timestamp 1713400504
transform 1 0 2888 0 -1 2370
box -8 -3 16 105
use FILL  FILL_923
timestamp 1713400504
transform 1 0 2880 0 -1 2370
box -8 -3 16 105
use FILL  FILL_924
timestamp 1713400504
transform 1 0 2832 0 -1 2370
box -8 -3 16 105
use FILL  FILL_925
timestamp 1713400504
transform 1 0 2824 0 -1 2370
box -8 -3 16 105
use FILL  FILL_926
timestamp 1713400504
transform 1 0 2816 0 -1 2370
box -8 -3 16 105
use FILL  FILL_927
timestamp 1713400504
transform 1 0 2808 0 -1 2370
box -8 -3 16 105
use FILL  FILL_928
timestamp 1713400504
transform 1 0 2784 0 -1 2370
box -8 -3 16 105
use FILL  FILL_929
timestamp 1713400504
transform 1 0 2776 0 -1 2370
box -8 -3 16 105
use FILL  FILL_930
timestamp 1713400504
transform 1 0 2768 0 -1 2370
box -8 -3 16 105
use FILL  FILL_931
timestamp 1713400504
transform 1 0 2760 0 -1 2370
box -8 -3 16 105
use FILL  FILL_932
timestamp 1713400504
transform 1 0 2712 0 -1 2370
box -8 -3 16 105
use FILL  FILL_933
timestamp 1713400504
transform 1 0 2704 0 -1 2370
box -8 -3 16 105
use FILL  FILL_934
timestamp 1713400504
transform 1 0 2696 0 -1 2370
box -8 -3 16 105
use FILL  FILL_935
timestamp 1713400504
transform 1 0 2688 0 -1 2370
box -8 -3 16 105
use FILL  FILL_936
timestamp 1713400504
transform 1 0 2680 0 -1 2370
box -8 -3 16 105
use FILL  FILL_937
timestamp 1713400504
transform 1 0 2672 0 -1 2370
box -8 -3 16 105
use FILL  FILL_938
timestamp 1713400504
transform 1 0 2632 0 -1 2370
box -8 -3 16 105
use FILL  FILL_939
timestamp 1713400504
transform 1 0 2608 0 -1 2370
box -8 -3 16 105
use FILL  FILL_940
timestamp 1713400504
transform 1 0 2600 0 -1 2370
box -8 -3 16 105
use FILL  FILL_941
timestamp 1713400504
transform 1 0 2592 0 -1 2370
box -8 -3 16 105
use FILL  FILL_942
timestamp 1713400504
transform 1 0 2584 0 -1 2370
box -8 -3 16 105
use FILL  FILL_943
timestamp 1713400504
transform 1 0 2576 0 -1 2370
box -8 -3 16 105
use FILL  FILL_944
timestamp 1713400504
transform 1 0 2512 0 -1 2370
box -8 -3 16 105
use FILL  FILL_945
timestamp 1713400504
transform 1 0 2504 0 -1 2370
box -8 -3 16 105
use FILL  FILL_946
timestamp 1713400504
transform 1 0 2496 0 -1 2370
box -8 -3 16 105
use FILL  FILL_947
timestamp 1713400504
transform 1 0 2488 0 -1 2370
box -8 -3 16 105
use FILL  FILL_948
timestamp 1713400504
transform 1 0 2480 0 -1 2370
box -8 -3 16 105
use FILL  FILL_949
timestamp 1713400504
transform 1 0 2472 0 -1 2370
box -8 -3 16 105
use FILL  FILL_950
timestamp 1713400504
transform 1 0 2464 0 -1 2370
box -8 -3 16 105
use FILL  FILL_951
timestamp 1713400504
transform 1 0 2408 0 -1 2370
box -8 -3 16 105
use FILL  FILL_952
timestamp 1713400504
transform 1 0 2400 0 -1 2370
box -8 -3 16 105
use FILL  FILL_953
timestamp 1713400504
transform 1 0 2392 0 -1 2370
box -8 -3 16 105
use FILL  FILL_954
timestamp 1713400504
transform 1 0 2384 0 -1 2370
box -8 -3 16 105
use FILL  FILL_955
timestamp 1713400504
transform 1 0 2376 0 -1 2370
box -8 -3 16 105
use FILL  FILL_956
timestamp 1713400504
transform 1 0 2368 0 -1 2370
box -8 -3 16 105
use FILL  FILL_957
timestamp 1713400504
transform 1 0 2336 0 -1 2370
box -8 -3 16 105
use FILL  FILL_958
timestamp 1713400504
transform 1 0 2328 0 -1 2370
box -8 -3 16 105
use FILL  FILL_959
timestamp 1713400504
transform 1 0 2288 0 -1 2370
box -8 -3 16 105
use FILL  FILL_960
timestamp 1713400504
transform 1 0 2280 0 -1 2370
box -8 -3 16 105
use FILL  FILL_961
timestamp 1713400504
transform 1 0 2272 0 -1 2370
box -8 -3 16 105
use FILL  FILL_962
timestamp 1713400504
transform 1 0 2264 0 -1 2370
box -8 -3 16 105
use FILL  FILL_963
timestamp 1713400504
transform 1 0 2256 0 -1 2370
box -8 -3 16 105
use FILL  FILL_964
timestamp 1713400504
transform 1 0 2224 0 -1 2370
box -8 -3 16 105
use FILL  FILL_965
timestamp 1713400504
transform 1 0 2216 0 -1 2370
box -8 -3 16 105
use FILL  FILL_966
timestamp 1713400504
transform 1 0 2208 0 -1 2370
box -8 -3 16 105
use FILL  FILL_967
timestamp 1713400504
transform 1 0 2184 0 -1 2370
box -8 -3 16 105
use FILL  FILL_968
timestamp 1713400504
transform 1 0 2176 0 -1 2370
box -8 -3 16 105
use FILL  FILL_969
timestamp 1713400504
transform 1 0 2168 0 -1 2370
box -8 -3 16 105
use FILL  FILL_970
timestamp 1713400504
transform 1 0 2064 0 -1 2370
box -8 -3 16 105
use FILL  FILL_971
timestamp 1713400504
transform 1 0 2056 0 -1 2370
box -8 -3 16 105
use FILL  FILL_972
timestamp 1713400504
transform 1 0 2048 0 -1 2370
box -8 -3 16 105
use FILL  FILL_973
timestamp 1713400504
transform 1 0 2040 0 -1 2370
box -8 -3 16 105
use FILL  FILL_974
timestamp 1713400504
transform 1 0 2008 0 -1 2370
box -8 -3 16 105
use FILL  FILL_975
timestamp 1713400504
transform 1 0 2000 0 -1 2370
box -8 -3 16 105
use FILL  FILL_976
timestamp 1713400504
transform 1 0 1992 0 -1 2370
box -8 -3 16 105
use FILL  FILL_977
timestamp 1713400504
transform 1 0 1984 0 -1 2370
box -8 -3 16 105
use FILL  FILL_978
timestamp 1713400504
transform 1 0 1952 0 -1 2370
box -8 -3 16 105
use FILL  FILL_979
timestamp 1713400504
transform 1 0 1944 0 -1 2370
box -8 -3 16 105
use FILL  FILL_980
timestamp 1713400504
transform 1 0 1936 0 -1 2370
box -8 -3 16 105
use FILL  FILL_981
timestamp 1713400504
transform 1 0 1928 0 -1 2370
box -8 -3 16 105
use FILL  FILL_982
timestamp 1713400504
transform 1 0 1920 0 -1 2370
box -8 -3 16 105
use FILL  FILL_983
timestamp 1713400504
transform 1 0 1912 0 -1 2370
box -8 -3 16 105
use FILL  FILL_984
timestamp 1713400504
transform 1 0 1880 0 -1 2370
box -8 -3 16 105
use FILL  FILL_985
timestamp 1713400504
transform 1 0 1872 0 -1 2370
box -8 -3 16 105
use FILL  FILL_986
timestamp 1713400504
transform 1 0 1864 0 -1 2370
box -8 -3 16 105
use FILL  FILL_987
timestamp 1713400504
transform 1 0 1832 0 -1 2370
box -8 -3 16 105
use FILL  FILL_988
timestamp 1713400504
transform 1 0 1824 0 -1 2370
box -8 -3 16 105
use FILL  FILL_989
timestamp 1713400504
transform 1 0 1816 0 -1 2370
box -8 -3 16 105
use FILL  FILL_990
timestamp 1713400504
transform 1 0 1808 0 -1 2370
box -8 -3 16 105
use FILL  FILL_991
timestamp 1713400504
transform 1 0 1800 0 -1 2370
box -8 -3 16 105
use FILL  FILL_992
timestamp 1713400504
transform 1 0 1696 0 -1 2370
box -8 -3 16 105
use FILL  FILL_993
timestamp 1713400504
transform 1 0 1592 0 -1 2370
box -8 -3 16 105
use FILL  FILL_994
timestamp 1713400504
transform 1 0 1584 0 -1 2370
box -8 -3 16 105
use FILL  FILL_995
timestamp 1713400504
transform 1 0 1576 0 -1 2370
box -8 -3 16 105
use FILL  FILL_996
timestamp 1713400504
transform 1 0 1568 0 -1 2370
box -8 -3 16 105
use FILL  FILL_997
timestamp 1713400504
transform 1 0 1560 0 -1 2370
box -8 -3 16 105
use FILL  FILL_998
timestamp 1713400504
transform 1 0 1520 0 -1 2370
box -8 -3 16 105
use FILL  FILL_999
timestamp 1713400504
transform 1 0 1512 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1000
timestamp 1713400504
transform 1 0 1504 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1001
timestamp 1713400504
transform 1 0 1496 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1002
timestamp 1713400504
transform 1 0 1488 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1003
timestamp 1713400504
transform 1 0 1480 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1004
timestamp 1713400504
transform 1 0 1472 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1005
timestamp 1713400504
transform 1 0 1424 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1006
timestamp 1713400504
transform 1 0 1416 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1007
timestamp 1713400504
transform 1 0 1408 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1008
timestamp 1713400504
transform 1 0 1400 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1009
timestamp 1713400504
transform 1 0 1392 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1010
timestamp 1713400504
transform 1 0 1384 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1011
timestamp 1713400504
transform 1 0 1376 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1012
timestamp 1713400504
transform 1 0 1344 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1013
timestamp 1713400504
transform 1 0 1336 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1014
timestamp 1713400504
transform 1 0 1328 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1015
timestamp 1713400504
transform 1 0 1304 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1016
timestamp 1713400504
transform 1 0 1296 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1017
timestamp 1713400504
transform 1 0 1288 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1018
timestamp 1713400504
transform 1 0 1280 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1019
timestamp 1713400504
transform 1 0 1272 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1020
timestamp 1713400504
transform 1 0 1264 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1021
timestamp 1713400504
transform 1 0 1256 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1022
timestamp 1713400504
transform 1 0 1248 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1023
timestamp 1713400504
transform 1 0 1208 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1024
timestamp 1713400504
transform 1 0 1200 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1025
timestamp 1713400504
transform 1 0 1192 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1026
timestamp 1713400504
transform 1 0 1184 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1027
timestamp 1713400504
transform 1 0 1176 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1028
timestamp 1713400504
transform 1 0 1168 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1029
timestamp 1713400504
transform 1 0 1160 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1030
timestamp 1713400504
transform 1 0 1152 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1031
timestamp 1713400504
transform 1 0 1112 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1032
timestamp 1713400504
transform 1 0 1104 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1033
timestamp 1713400504
transform 1 0 1096 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1034
timestamp 1713400504
transform 1 0 1088 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1035
timestamp 1713400504
transform 1 0 1080 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1036
timestamp 1713400504
transform 1 0 1072 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1037
timestamp 1713400504
transform 1 0 1064 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1038
timestamp 1713400504
transform 1 0 1056 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1039
timestamp 1713400504
transform 1 0 1048 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1040
timestamp 1713400504
transform 1 0 1000 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1041
timestamp 1713400504
transform 1 0 992 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1042
timestamp 1713400504
transform 1 0 984 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1043
timestamp 1713400504
transform 1 0 976 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1044
timestamp 1713400504
transform 1 0 968 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1045
timestamp 1713400504
transform 1 0 960 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1046
timestamp 1713400504
transform 1 0 952 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1047
timestamp 1713400504
transform 1 0 928 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1048
timestamp 1713400504
transform 1 0 920 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1049
timestamp 1713400504
transform 1 0 912 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1050
timestamp 1713400504
transform 1 0 904 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1051
timestamp 1713400504
transform 1 0 896 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1052
timestamp 1713400504
transform 1 0 888 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1053
timestamp 1713400504
transform 1 0 840 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1054
timestamp 1713400504
transform 1 0 832 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1055
timestamp 1713400504
transform 1 0 824 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1056
timestamp 1713400504
transform 1 0 816 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1057
timestamp 1713400504
transform 1 0 808 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1058
timestamp 1713400504
transform 1 0 800 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1059
timestamp 1713400504
transform 1 0 712 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1060
timestamp 1713400504
transform 1 0 704 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1061
timestamp 1713400504
transform 1 0 696 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1062
timestamp 1713400504
transform 1 0 688 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1063
timestamp 1713400504
transform 1 0 656 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1064
timestamp 1713400504
transform 1 0 648 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1065
timestamp 1713400504
transform 1 0 640 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1066
timestamp 1713400504
transform 1 0 632 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1067
timestamp 1713400504
transform 1 0 504 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1068
timestamp 1713400504
transform 1 0 496 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1069
timestamp 1713400504
transform 1 0 488 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1070
timestamp 1713400504
transform 1 0 360 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1071
timestamp 1713400504
transform 1 0 352 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1072
timestamp 1713400504
transform 1 0 344 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1073
timestamp 1713400504
transform 1 0 336 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1074
timestamp 1713400504
transform 1 0 304 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1075
timestamp 1713400504
transform 1 0 296 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1076
timestamp 1713400504
transform 1 0 288 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1077
timestamp 1713400504
transform 1 0 280 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1078
timestamp 1713400504
transform 1 0 256 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1079
timestamp 1713400504
transform 1 0 248 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1080
timestamp 1713400504
transform 1 0 240 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1081
timestamp 1713400504
transform 1 0 232 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1082
timestamp 1713400504
transform 1 0 224 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1083
timestamp 1713400504
transform 1 0 168 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1084
timestamp 1713400504
transform 1 0 160 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1085
timestamp 1713400504
transform 1 0 152 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1086
timestamp 1713400504
transform 1 0 144 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1087
timestamp 1713400504
transform 1 0 136 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1088
timestamp 1713400504
transform 1 0 96 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1089
timestamp 1713400504
transform 1 0 88 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1090
timestamp 1713400504
transform 1 0 80 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1091
timestamp 1713400504
transform 1 0 72 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1092
timestamp 1713400504
transform 1 0 3008 0 1 2170
box -8 -3 16 105
use FILL  FILL_1093
timestamp 1713400504
transform 1 0 2904 0 1 2170
box -8 -3 16 105
use FILL  FILL_1094
timestamp 1713400504
transform 1 0 2896 0 1 2170
box -8 -3 16 105
use FILL  FILL_1095
timestamp 1713400504
transform 1 0 2888 0 1 2170
box -8 -3 16 105
use FILL  FILL_1096
timestamp 1713400504
transform 1 0 2880 0 1 2170
box -8 -3 16 105
use FILL  FILL_1097
timestamp 1713400504
transform 1 0 2856 0 1 2170
box -8 -3 16 105
use FILL  FILL_1098
timestamp 1713400504
transform 1 0 2848 0 1 2170
box -8 -3 16 105
use FILL  FILL_1099
timestamp 1713400504
transform 1 0 2744 0 1 2170
box -8 -3 16 105
use FILL  FILL_1100
timestamp 1713400504
transform 1 0 2736 0 1 2170
box -8 -3 16 105
use FILL  FILL_1101
timestamp 1713400504
transform 1 0 2728 0 1 2170
box -8 -3 16 105
use FILL  FILL_1102
timestamp 1713400504
transform 1 0 2720 0 1 2170
box -8 -3 16 105
use FILL  FILL_1103
timestamp 1713400504
transform 1 0 2680 0 1 2170
box -8 -3 16 105
use FILL  FILL_1104
timestamp 1713400504
transform 1 0 2672 0 1 2170
box -8 -3 16 105
use FILL  FILL_1105
timestamp 1713400504
transform 1 0 2664 0 1 2170
box -8 -3 16 105
use FILL  FILL_1106
timestamp 1713400504
transform 1 0 2656 0 1 2170
box -8 -3 16 105
use FILL  FILL_1107
timestamp 1713400504
transform 1 0 2624 0 1 2170
box -8 -3 16 105
use FILL  FILL_1108
timestamp 1713400504
transform 1 0 2616 0 1 2170
box -8 -3 16 105
use FILL  FILL_1109
timestamp 1713400504
transform 1 0 2608 0 1 2170
box -8 -3 16 105
use FILL  FILL_1110
timestamp 1713400504
transform 1 0 2600 0 1 2170
box -8 -3 16 105
use FILL  FILL_1111
timestamp 1713400504
transform 1 0 2560 0 1 2170
box -8 -3 16 105
use FILL  FILL_1112
timestamp 1713400504
transform 1 0 2552 0 1 2170
box -8 -3 16 105
use FILL  FILL_1113
timestamp 1713400504
transform 1 0 2544 0 1 2170
box -8 -3 16 105
use FILL  FILL_1114
timestamp 1713400504
transform 1 0 2512 0 1 2170
box -8 -3 16 105
use FILL  FILL_1115
timestamp 1713400504
transform 1 0 2504 0 1 2170
box -8 -3 16 105
use FILL  FILL_1116
timestamp 1713400504
transform 1 0 2496 0 1 2170
box -8 -3 16 105
use FILL  FILL_1117
timestamp 1713400504
transform 1 0 2464 0 1 2170
box -8 -3 16 105
use FILL  FILL_1118
timestamp 1713400504
transform 1 0 2456 0 1 2170
box -8 -3 16 105
use FILL  FILL_1119
timestamp 1713400504
transform 1 0 2448 0 1 2170
box -8 -3 16 105
use FILL  FILL_1120
timestamp 1713400504
transform 1 0 2440 0 1 2170
box -8 -3 16 105
use FILL  FILL_1121
timestamp 1713400504
transform 1 0 2416 0 1 2170
box -8 -3 16 105
use FILL  FILL_1122
timestamp 1713400504
transform 1 0 2408 0 1 2170
box -8 -3 16 105
use FILL  FILL_1123
timestamp 1713400504
transform 1 0 2400 0 1 2170
box -8 -3 16 105
use FILL  FILL_1124
timestamp 1713400504
transform 1 0 2368 0 1 2170
box -8 -3 16 105
use FILL  FILL_1125
timestamp 1713400504
transform 1 0 2360 0 1 2170
box -8 -3 16 105
use FILL  FILL_1126
timestamp 1713400504
transform 1 0 2352 0 1 2170
box -8 -3 16 105
use FILL  FILL_1127
timestamp 1713400504
transform 1 0 2344 0 1 2170
box -8 -3 16 105
use FILL  FILL_1128
timestamp 1713400504
transform 1 0 2336 0 1 2170
box -8 -3 16 105
use FILL  FILL_1129
timestamp 1713400504
transform 1 0 2296 0 1 2170
box -8 -3 16 105
use FILL  FILL_1130
timestamp 1713400504
transform 1 0 2288 0 1 2170
box -8 -3 16 105
use FILL  FILL_1131
timestamp 1713400504
transform 1 0 2280 0 1 2170
box -8 -3 16 105
use FILL  FILL_1132
timestamp 1713400504
transform 1 0 2272 0 1 2170
box -8 -3 16 105
use FILL  FILL_1133
timestamp 1713400504
transform 1 0 2264 0 1 2170
box -8 -3 16 105
use FILL  FILL_1134
timestamp 1713400504
transform 1 0 2232 0 1 2170
box -8 -3 16 105
use FILL  FILL_1135
timestamp 1713400504
transform 1 0 2224 0 1 2170
box -8 -3 16 105
use FILL  FILL_1136
timestamp 1713400504
transform 1 0 2216 0 1 2170
box -8 -3 16 105
use FILL  FILL_1137
timestamp 1713400504
transform 1 0 2184 0 1 2170
box -8 -3 16 105
use FILL  FILL_1138
timestamp 1713400504
transform 1 0 2152 0 1 2170
box -8 -3 16 105
use FILL  FILL_1139
timestamp 1713400504
transform 1 0 2144 0 1 2170
box -8 -3 16 105
use FILL  FILL_1140
timestamp 1713400504
transform 1 0 2136 0 1 2170
box -8 -3 16 105
use FILL  FILL_1141
timestamp 1713400504
transform 1 0 2128 0 1 2170
box -8 -3 16 105
use FILL  FILL_1142
timestamp 1713400504
transform 1 0 2104 0 1 2170
box -8 -3 16 105
use FILL  FILL_1143
timestamp 1713400504
transform 1 0 2096 0 1 2170
box -8 -3 16 105
use FILL  FILL_1144
timestamp 1713400504
transform 1 0 2088 0 1 2170
box -8 -3 16 105
use FILL  FILL_1145
timestamp 1713400504
transform 1 0 2080 0 1 2170
box -8 -3 16 105
use FILL  FILL_1146
timestamp 1713400504
transform 1 0 2040 0 1 2170
box -8 -3 16 105
use FILL  FILL_1147
timestamp 1713400504
transform 1 0 2032 0 1 2170
box -8 -3 16 105
use FILL  FILL_1148
timestamp 1713400504
transform 1 0 2024 0 1 2170
box -8 -3 16 105
use FILL  FILL_1149
timestamp 1713400504
transform 1 0 2016 0 1 2170
box -8 -3 16 105
use FILL  FILL_1150
timestamp 1713400504
transform 1 0 2008 0 1 2170
box -8 -3 16 105
use FILL  FILL_1151
timestamp 1713400504
transform 1 0 2000 0 1 2170
box -8 -3 16 105
use FILL  FILL_1152
timestamp 1713400504
transform 1 0 1960 0 1 2170
box -8 -3 16 105
use FILL  FILL_1153
timestamp 1713400504
transform 1 0 1952 0 1 2170
box -8 -3 16 105
use FILL  FILL_1154
timestamp 1713400504
transform 1 0 1944 0 1 2170
box -8 -3 16 105
use FILL  FILL_1155
timestamp 1713400504
transform 1 0 1936 0 1 2170
box -8 -3 16 105
use FILL  FILL_1156
timestamp 1713400504
transform 1 0 1928 0 1 2170
box -8 -3 16 105
use FILL  FILL_1157
timestamp 1713400504
transform 1 0 1896 0 1 2170
box -8 -3 16 105
use FILL  FILL_1158
timestamp 1713400504
transform 1 0 1888 0 1 2170
box -8 -3 16 105
use FILL  FILL_1159
timestamp 1713400504
transform 1 0 1880 0 1 2170
box -8 -3 16 105
use FILL  FILL_1160
timestamp 1713400504
transform 1 0 1848 0 1 2170
box -8 -3 16 105
use FILL  FILL_1161
timestamp 1713400504
transform 1 0 1840 0 1 2170
box -8 -3 16 105
use FILL  FILL_1162
timestamp 1713400504
transform 1 0 1832 0 1 2170
box -8 -3 16 105
use FILL  FILL_1163
timestamp 1713400504
transform 1 0 1824 0 1 2170
box -8 -3 16 105
use FILL  FILL_1164
timestamp 1713400504
transform 1 0 1816 0 1 2170
box -8 -3 16 105
use FILL  FILL_1165
timestamp 1713400504
transform 1 0 1808 0 1 2170
box -8 -3 16 105
use FILL  FILL_1166
timestamp 1713400504
transform 1 0 1768 0 1 2170
box -8 -3 16 105
use FILL  FILL_1167
timestamp 1713400504
transform 1 0 1760 0 1 2170
box -8 -3 16 105
use FILL  FILL_1168
timestamp 1713400504
transform 1 0 1752 0 1 2170
box -8 -3 16 105
use FILL  FILL_1169
timestamp 1713400504
transform 1 0 1728 0 1 2170
box -8 -3 16 105
use FILL  FILL_1170
timestamp 1713400504
transform 1 0 1720 0 1 2170
box -8 -3 16 105
use FILL  FILL_1171
timestamp 1713400504
transform 1 0 1712 0 1 2170
box -8 -3 16 105
use FILL  FILL_1172
timestamp 1713400504
transform 1 0 1704 0 1 2170
box -8 -3 16 105
use FILL  FILL_1173
timestamp 1713400504
transform 1 0 1696 0 1 2170
box -8 -3 16 105
use FILL  FILL_1174
timestamp 1713400504
transform 1 0 1688 0 1 2170
box -8 -3 16 105
use FILL  FILL_1175
timestamp 1713400504
transform 1 0 1640 0 1 2170
box -8 -3 16 105
use FILL  FILL_1176
timestamp 1713400504
transform 1 0 1632 0 1 2170
box -8 -3 16 105
use FILL  FILL_1177
timestamp 1713400504
transform 1 0 1624 0 1 2170
box -8 -3 16 105
use FILL  FILL_1178
timestamp 1713400504
transform 1 0 1616 0 1 2170
box -8 -3 16 105
use FILL  FILL_1179
timestamp 1713400504
transform 1 0 1608 0 1 2170
box -8 -3 16 105
use FILL  FILL_1180
timestamp 1713400504
transform 1 0 1600 0 1 2170
box -8 -3 16 105
use FILL  FILL_1181
timestamp 1713400504
transform 1 0 1568 0 1 2170
box -8 -3 16 105
use FILL  FILL_1182
timestamp 1713400504
transform 1 0 1544 0 1 2170
box -8 -3 16 105
use FILL  FILL_1183
timestamp 1713400504
transform 1 0 1536 0 1 2170
box -8 -3 16 105
use FILL  FILL_1184
timestamp 1713400504
transform 1 0 1528 0 1 2170
box -8 -3 16 105
use FILL  FILL_1185
timestamp 1713400504
transform 1 0 1520 0 1 2170
box -8 -3 16 105
use FILL  FILL_1186
timestamp 1713400504
transform 1 0 1512 0 1 2170
box -8 -3 16 105
use FILL  FILL_1187
timestamp 1713400504
transform 1 0 1480 0 1 2170
box -8 -3 16 105
use FILL  FILL_1188
timestamp 1713400504
transform 1 0 1472 0 1 2170
box -8 -3 16 105
use FILL  FILL_1189
timestamp 1713400504
transform 1 0 1464 0 1 2170
box -8 -3 16 105
use FILL  FILL_1190
timestamp 1713400504
transform 1 0 1456 0 1 2170
box -8 -3 16 105
use FILL  FILL_1191
timestamp 1713400504
transform 1 0 1352 0 1 2170
box -8 -3 16 105
use FILL  FILL_1192
timestamp 1713400504
transform 1 0 1344 0 1 2170
box -8 -3 16 105
use FILL  FILL_1193
timestamp 1713400504
transform 1 0 1336 0 1 2170
box -8 -3 16 105
use FILL  FILL_1194
timestamp 1713400504
transform 1 0 1328 0 1 2170
box -8 -3 16 105
use FILL  FILL_1195
timestamp 1713400504
transform 1 0 1320 0 1 2170
box -8 -3 16 105
use FILL  FILL_1196
timestamp 1713400504
transform 1 0 1312 0 1 2170
box -8 -3 16 105
use FILL  FILL_1197
timestamp 1713400504
transform 1 0 1264 0 1 2170
box -8 -3 16 105
use FILL  FILL_1198
timestamp 1713400504
transform 1 0 1256 0 1 2170
box -8 -3 16 105
use FILL  FILL_1199
timestamp 1713400504
transform 1 0 1248 0 1 2170
box -8 -3 16 105
use FILL  FILL_1200
timestamp 1713400504
transform 1 0 1240 0 1 2170
box -8 -3 16 105
use FILL  FILL_1201
timestamp 1713400504
transform 1 0 1232 0 1 2170
box -8 -3 16 105
use FILL  FILL_1202
timestamp 1713400504
transform 1 0 1224 0 1 2170
box -8 -3 16 105
use FILL  FILL_1203
timestamp 1713400504
transform 1 0 1216 0 1 2170
box -8 -3 16 105
use FILL  FILL_1204
timestamp 1713400504
transform 1 0 1208 0 1 2170
box -8 -3 16 105
use FILL  FILL_1205
timestamp 1713400504
transform 1 0 1200 0 1 2170
box -8 -3 16 105
use FILL  FILL_1206
timestamp 1713400504
transform 1 0 1176 0 1 2170
box -8 -3 16 105
use FILL  FILL_1207
timestamp 1713400504
transform 1 0 1168 0 1 2170
box -8 -3 16 105
use FILL  FILL_1208
timestamp 1713400504
transform 1 0 1160 0 1 2170
box -8 -3 16 105
use FILL  FILL_1209
timestamp 1713400504
transform 1 0 1152 0 1 2170
box -8 -3 16 105
use FILL  FILL_1210
timestamp 1713400504
transform 1 0 1144 0 1 2170
box -8 -3 16 105
use FILL  FILL_1211
timestamp 1713400504
transform 1 0 1136 0 1 2170
box -8 -3 16 105
use FILL  FILL_1212
timestamp 1713400504
transform 1 0 1128 0 1 2170
box -8 -3 16 105
use FILL  FILL_1213
timestamp 1713400504
transform 1 0 1120 0 1 2170
box -8 -3 16 105
use FILL  FILL_1214
timestamp 1713400504
transform 1 0 1112 0 1 2170
box -8 -3 16 105
use FILL  FILL_1215
timestamp 1713400504
transform 1 0 1104 0 1 2170
box -8 -3 16 105
use FILL  FILL_1216
timestamp 1713400504
transform 1 0 1064 0 1 2170
box -8 -3 16 105
use FILL  FILL_1217
timestamp 1713400504
transform 1 0 1056 0 1 2170
box -8 -3 16 105
use FILL  FILL_1218
timestamp 1713400504
transform 1 0 1048 0 1 2170
box -8 -3 16 105
use FILL  FILL_1219
timestamp 1713400504
transform 1 0 1040 0 1 2170
box -8 -3 16 105
use FILL  FILL_1220
timestamp 1713400504
transform 1 0 1032 0 1 2170
box -8 -3 16 105
use FILL  FILL_1221
timestamp 1713400504
transform 1 0 1024 0 1 2170
box -8 -3 16 105
use FILL  FILL_1222
timestamp 1713400504
transform 1 0 1016 0 1 2170
box -8 -3 16 105
use FILL  FILL_1223
timestamp 1713400504
transform 1 0 1008 0 1 2170
box -8 -3 16 105
use FILL  FILL_1224
timestamp 1713400504
transform 1 0 1000 0 1 2170
box -8 -3 16 105
use FILL  FILL_1225
timestamp 1713400504
transform 1 0 992 0 1 2170
box -8 -3 16 105
use FILL  FILL_1226
timestamp 1713400504
transform 1 0 984 0 1 2170
box -8 -3 16 105
use FILL  FILL_1227
timestamp 1713400504
transform 1 0 936 0 1 2170
box -8 -3 16 105
use FILL  FILL_1228
timestamp 1713400504
transform 1 0 928 0 1 2170
box -8 -3 16 105
use FILL  FILL_1229
timestamp 1713400504
transform 1 0 920 0 1 2170
box -8 -3 16 105
use FILL  FILL_1230
timestamp 1713400504
transform 1 0 912 0 1 2170
box -8 -3 16 105
use FILL  FILL_1231
timestamp 1713400504
transform 1 0 904 0 1 2170
box -8 -3 16 105
use FILL  FILL_1232
timestamp 1713400504
transform 1 0 896 0 1 2170
box -8 -3 16 105
use FILL  FILL_1233
timestamp 1713400504
transform 1 0 888 0 1 2170
box -8 -3 16 105
use FILL  FILL_1234
timestamp 1713400504
transform 1 0 880 0 1 2170
box -8 -3 16 105
use FILL  FILL_1235
timestamp 1713400504
transform 1 0 872 0 1 2170
box -8 -3 16 105
use FILL  FILL_1236
timestamp 1713400504
transform 1 0 840 0 1 2170
box -8 -3 16 105
use FILL  FILL_1237
timestamp 1713400504
transform 1 0 832 0 1 2170
box -8 -3 16 105
use FILL  FILL_1238
timestamp 1713400504
transform 1 0 824 0 1 2170
box -8 -3 16 105
use FILL  FILL_1239
timestamp 1713400504
transform 1 0 816 0 1 2170
box -8 -3 16 105
use FILL  FILL_1240
timestamp 1713400504
transform 1 0 808 0 1 2170
box -8 -3 16 105
use FILL  FILL_1241
timestamp 1713400504
transform 1 0 800 0 1 2170
box -8 -3 16 105
use FILL  FILL_1242
timestamp 1713400504
transform 1 0 792 0 1 2170
box -8 -3 16 105
use FILL  FILL_1243
timestamp 1713400504
transform 1 0 784 0 1 2170
box -8 -3 16 105
use FILL  FILL_1244
timestamp 1713400504
transform 1 0 776 0 1 2170
box -8 -3 16 105
use FILL  FILL_1245
timestamp 1713400504
transform 1 0 744 0 1 2170
box -8 -3 16 105
use FILL  FILL_1246
timestamp 1713400504
transform 1 0 736 0 1 2170
box -8 -3 16 105
use FILL  FILL_1247
timestamp 1713400504
transform 1 0 728 0 1 2170
box -8 -3 16 105
use FILL  FILL_1248
timestamp 1713400504
transform 1 0 720 0 1 2170
box -8 -3 16 105
use FILL  FILL_1249
timestamp 1713400504
transform 1 0 712 0 1 2170
box -8 -3 16 105
use FILL  FILL_1250
timestamp 1713400504
transform 1 0 704 0 1 2170
box -8 -3 16 105
use FILL  FILL_1251
timestamp 1713400504
transform 1 0 672 0 1 2170
box -8 -3 16 105
use FILL  FILL_1252
timestamp 1713400504
transform 1 0 664 0 1 2170
box -8 -3 16 105
use FILL  FILL_1253
timestamp 1713400504
transform 1 0 656 0 1 2170
box -8 -3 16 105
use FILL  FILL_1254
timestamp 1713400504
transform 1 0 648 0 1 2170
box -8 -3 16 105
use FILL  FILL_1255
timestamp 1713400504
transform 1 0 640 0 1 2170
box -8 -3 16 105
use FILL  FILL_1256
timestamp 1713400504
transform 1 0 512 0 1 2170
box -8 -3 16 105
use FILL  FILL_1257
timestamp 1713400504
transform 1 0 504 0 1 2170
box -8 -3 16 105
use FILL  FILL_1258
timestamp 1713400504
transform 1 0 416 0 1 2170
box -8 -3 16 105
use FILL  FILL_1259
timestamp 1713400504
transform 1 0 408 0 1 2170
box -8 -3 16 105
use FILL  FILL_1260
timestamp 1713400504
transform 1 0 400 0 1 2170
box -8 -3 16 105
use FILL  FILL_1261
timestamp 1713400504
transform 1 0 392 0 1 2170
box -8 -3 16 105
use FILL  FILL_1262
timestamp 1713400504
transform 1 0 360 0 1 2170
box -8 -3 16 105
use FILL  FILL_1263
timestamp 1713400504
transform 1 0 352 0 1 2170
box -8 -3 16 105
use FILL  FILL_1264
timestamp 1713400504
transform 1 0 344 0 1 2170
box -8 -3 16 105
use FILL  FILL_1265
timestamp 1713400504
transform 1 0 216 0 1 2170
box -8 -3 16 105
use FILL  FILL_1266
timestamp 1713400504
transform 1 0 208 0 1 2170
box -8 -3 16 105
use FILL  FILL_1267
timestamp 1713400504
transform 1 0 184 0 1 2170
box -8 -3 16 105
use FILL  FILL_1268
timestamp 1713400504
transform 1 0 176 0 1 2170
box -8 -3 16 105
use FILL  FILL_1269
timestamp 1713400504
transform 1 0 168 0 1 2170
box -8 -3 16 105
use FILL  FILL_1270
timestamp 1713400504
transform 1 0 160 0 1 2170
box -8 -3 16 105
use FILL  FILL_1271
timestamp 1713400504
transform 1 0 152 0 1 2170
box -8 -3 16 105
use FILL  FILL_1272
timestamp 1713400504
transform 1 0 128 0 1 2170
box -8 -3 16 105
use FILL  FILL_1273
timestamp 1713400504
transform 1 0 120 0 1 2170
box -8 -3 16 105
use FILL  FILL_1274
timestamp 1713400504
transform 1 0 80 0 1 2170
box -8 -3 16 105
use FILL  FILL_1275
timestamp 1713400504
transform 1 0 72 0 1 2170
box -8 -3 16 105
use FILL  FILL_1276
timestamp 1713400504
transform 1 0 3008 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1277
timestamp 1713400504
transform 1 0 2984 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1278
timestamp 1713400504
transform 1 0 2976 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1279
timestamp 1713400504
transform 1 0 2968 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1280
timestamp 1713400504
transform 1 0 2960 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1281
timestamp 1713400504
transform 1 0 2952 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1282
timestamp 1713400504
transform 1 0 2944 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1283
timestamp 1713400504
transform 1 0 2936 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1284
timestamp 1713400504
transform 1 0 2888 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1285
timestamp 1713400504
transform 1 0 2880 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1286
timestamp 1713400504
transform 1 0 2872 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1287
timestamp 1713400504
transform 1 0 2864 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1288
timestamp 1713400504
transform 1 0 2760 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1289
timestamp 1713400504
transform 1 0 2752 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1290
timestamp 1713400504
transform 1 0 2744 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1291
timestamp 1713400504
transform 1 0 2736 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1292
timestamp 1713400504
transform 1 0 2696 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1293
timestamp 1713400504
transform 1 0 2688 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1294
timestamp 1713400504
transform 1 0 2680 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1295
timestamp 1713400504
transform 1 0 2672 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1296
timestamp 1713400504
transform 1 0 2664 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1297
timestamp 1713400504
transform 1 0 2656 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1298
timestamp 1713400504
transform 1 0 2616 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1299
timestamp 1713400504
transform 1 0 2608 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1300
timestamp 1713400504
transform 1 0 2600 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1301
timestamp 1713400504
transform 1 0 2592 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1302
timestamp 1713400504
transform 1 0 2568 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1303
timestamp 1713400504
transform 1 0 2560 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1304
timestamp 1713400504
transform 1 0 2552 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1305
timestamp 1713400504
transform 1 0 2544 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1306
timestamp 1713400504
transform 1 0 2440 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1307
timestamp 1713400504
transform 1 0 2432 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1308
timestamp 1713400504
transform 1 0 2424 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1309
timestamp 1713400504
transform 1 0 2416 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1310
timestamp 1713400504
transform 1 0 2384 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1311
timestamp 1713400504
transform 1 0 2376 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1312
timestamp 1713400504
transform 1 0 2368 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1313
timestamp 1713400504
transform 1 0 2360 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1314
timestamp 1713400504
transform 1 0 2328 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1315
timestamp 1713400504
transform 1 0 2320 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1316
timestamp 1713400504
transform 1 0 2312 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1317
timestamp 1713400504
transform 1 0 2304 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1318
timestamp 1713400504
transform 1 0 2200 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1319
timestamp 1713400504
transform 1 0 2192 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1320
timestamp 1713400504
transform 1 0 2184 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1321
timestamp 1713400504
transform 1 0 2136 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1322
timestamp 1713400504
transform 1 0 2128 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1323
timestamp 1713400504
transform 1 0 2120 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1324
timestamp 1713400504
transform 1 0 2112 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1325
timestamp 1713400504
transform 1 0 2104 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1326
timestamp 1713400504
transform 1 0 2080 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1327
timestamp 1713400504
transform 1 0 2072 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1328
timestamp 1713400504
transform 1 0 2064 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1329
timestamp 1713400504
transform 1 0 2032 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1330
timestamp 1713400504
transform 1 0 2024 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1331
timestamp 1713400504
transform 1 0 2016 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1332
timestamp 1713400504
transform 1 0 2008 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1333
timestamp 1713400504
transform 1 0 1976 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1334
timestamp 1713400504
transform 1 0 1968 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1335
timestamp 1713400504
transform 1 0 1960 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1336
timestamp 1713400504
transform 1 0 1952 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1337
timestamp 1713400504
transform 1 0 1912 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1338
timestamp 1713400504
transform 1 0 1904 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1339
timestamp 1713400504
transform 1 0 1896 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1340
timestamp 1713400504
transform 1 0 1792 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1341
timestamp 1713400504
transform 1 0 1784 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1342
timestamp 1713400504
transform 1 0 1776 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1343
timestamp 1713400504
transform 1 0 1728 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1344
timestamp 1713400504
transform 1 0 1720 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1345
timestamp 1713400504
transform 1 0 1712 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1346
timestamp 1713400504
transform 1 0 1704 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1347
timestamp 1713400504
transform 1 0 1664 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1348
timestamp 1713400504
transform 1 0 1656 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1349
timestamp 1713400504
transform 1 0 1648 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1350
timestamp 1713400504
transform 1 0 1640 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1351
timestamp 1713400504
transform 1 0 1632 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1352
timestamp 1713400504
transform 1 0 1592 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1353
timestamp 1713400504
transform 1 0 1584 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1354
timestamp 1713400504
transform 1 0 1576 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1355
timestamp 1713400504
transform 1 0 1568 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1356
timestamp 1713400504
transform 1 0 1528 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1357
timestamp 1713400504
transform 1 0 1520 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1358
timestamp 1713400504
transform 1 0 1512 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1359
timestamp 1713400504
transform 1 0 1504 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1360
timestamp 1713400504
transform 1 0 1496 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1361
timestamp 1713400504
transform 1 0 1488 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1362
timestamp 1713400504
transform 1 0 1440 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1363
timestamp 1713400504
transform 1 0 1432 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1364
timestamp 1713400504
transform 1 0 1424 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1365
timestamp 1713400504
transform 1 0 1416 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1366
timestamp 1713400504
transform 1 0 1392 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1367
timestamp 1713400504
transform 1 0 1384 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1368
timestamp 1713400504
transform 1 0 1376 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1369
timestamp 1713400504
transform 1 0 1368 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1370
timestamp 1713400504
transform 1 0 1360 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1371
timestamp 1713400504
transform 1 0 1320 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1372
timestamp 1713400504
transform 1 0 1312 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1373
timestamp 1713400504
transform 1 0 1304 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1374
timestamp 1713400504
transform 1 0 1296 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1375
timestamp 1713400504
transform 1 0 1288 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1376
timestamp 1713400504
transform 1 0 1280 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1377
timestamp 1713400504
transform 1 0 1272 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1378
timestamp 1713400504
transform 1 0 1232 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1379
timestamp 1713400504
transform 1 0 1224 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1380
timestamp 1713400504
transform 1 0 1216 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1381
timestamp 1713400504
transform 1 0 1208 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1382
timestamp 1713400504
transform 1 0 1200 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1383
timestamp 1713400504
transform 1 0 1192 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1384
timestamp 1713400504
transform 1 0 1152 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1385
timestamp 1713400504
transform 1 0 1144 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1386
timestamp 1713400504
transform 1 0 1136 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1387
timestamp 1713400504
transform 1 0 1128 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1388
timestamp 1713400504
transform 1 0 1120 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1389
timestamp 1713400504
transform 1 0 1112 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1390
timestamp 1713400504
transform 1 0 1104 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1391
timestamp 1713400504
transform 1 0 1096 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1392
timestamp 1713400504
transform 1 0 1048 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1393
timestamp 1713400504
transform 1 0 1040 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1394
timestamp 1713400504
transform 1 0 1032 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1395
timestamp 1713400504
transform 1 0 1024 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1396
timestamp 1713400504
transform 1 0 1016 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1397
timestamp 1713400504
transform 1 0 1008 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1398
timestamp 1713400504
transform 1 0 1000 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1399
timestamp 1713400504
transform 1 0 992 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1400
timestamp 1713400504
transform 1 0 944 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1401
timestamp 1713400504
transform 1 0 936 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1402
timestamp 1713400504
transform 1 0 928 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1403
timestamp 1713400504
transform 1 0 920 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1404
timestamp 1713400504
transform 1 0 912 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1405
timestamp 1713400504
transform 1 0 904 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1406
timestamp 1713400504
transform 1 0 896 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1407
timestamp 1713400504
transform 1 0 856 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1408
timestamp 1713400504
transform 1 0 848 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1409
timestamp 1713400504
transform 1 0 840 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1410
timestamp 1713400504
transform 1 0 832 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1411
timestamp 1713400504
transform 1 0 824 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1412
timestamp 1713400504
transform 1 0 696 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1413
timestamp 1713400504
transform 1 0 688 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1414
timestamp 1713400504
transform 1 0 656 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1415
timestamp 1713400504
transform 1 0 648 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1416
timestamp 1713400504
transform 1 0 640 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1417
timestamp 1713400504
transform 1 0 632 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1418
timestamp 1713400504
transform 1 0 624 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1419
timestamp 1713400504
transform 1 0 592 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1420
timestamp 1713400504
transform 1 0 584 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1421
timestamp 1713400504
transform 1 0 576 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1422
timestamp 1713400504
transform 1 0 568 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1423
timestamp 1713400504
transform 1 0 536 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1424
timestamp 1713400504
transform 1 0 528 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1425
timestamp 1713400504
transform 1 0 520 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1426
timestamp 1713400504
transform 1 0 512 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1427
timestamp 1713400504
transform 1 0 480 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1428
timestamp 1713400504
transform 1 0 472 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1429
timestamp 1713400504
transform 1 0 464 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1430
timestamp 1713400504
transform 1 0 376 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1431
timestamp 1713400504
transform 1 0 368 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1432
timestamp 1713400504
transform 1 0 336 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1433
timestamp 1713400504
transform 1 0 328 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1434
timestamp 1713400504
transform 1 0 320 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1435
timestamp 1713400504
transform 1 0 312 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1436
timestamp 1713400504
transform 1 0 304 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1437
timestamp 1713400504
transform 1 0 264 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1438
timestamp 1713400504
transform 1 0 256 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1439
timestamp 1713400504
transform 1 0 248 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1440
timestamp 1713400504
transform 1 0 240 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1441
timestamp 1713400504
transform 1 0 232 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1442
timestamp 1713400504
transform 1 0 224 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1443
timestamp 1713400504
transform 1 0 168 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1444
timestamp 1713400504
transform 1 0 160 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1445
timestamp 1713400504
transform 1 0 72 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1446
timestamp 1713400504
transform 1 0 3008 0 1 1970
box -8 -3 16 105
use FILL  FILL_1447
timestamp 1713400504
transform 1 0 3000 0 1 1970
box -8 -3 16 105
use FILL  FILL_1448
timestamp 1713400504
transform 1 0 2992 0 1 1970
box -8 -3 16 105
use FILL  FILL_1449
timestamp 1713400504
transform 1 0 2968 0 1 1970
box -8 -3 16 105
use FILL  FILL_1450
timestamp 1713400504
transform 1 0 2960 0 1 1970
box -8 -3 16 105
use FILL  FILL_1451
timestamp 1713400504
transform 1 0 2928 0 1 1970
box -8 -3 16 105
use FILL  FILL_1452
timestamp 1713400504
transform 1 0 2920 0 1 1970
box -8 -3 16 105
use FILL  FILL_1453
timestamp 1713400504
transform 1 0 2912 0 1 1970
box -8 -3 16 105
use FILL  FILL_1454
timestamp 1713400504
transform 1 0 2904 0 1 1970
box -8 -3 16 105
use FILL  FILL_1455
timestamp 1713400504
transform 1 0 2896 0 1 1970
box -8 -3 16 105
use FILL  FILL_1456
timestamp 1713400504
transform 1 0 2856 0 1 1970
box -8 -3 16 105
use FILL  FILL_1457
timestamp 1713400504
transform 1 0 2848 0 1 1970
box -8 -3 16 105
use FILL  FILL_1458
timestamp 1713400504
transform 1 0 2840 0 1 1970
box -8 -3 16 105
use FILL  FILL_1459
timestamp 1713400504
transform 1 0 2832 0 1 1970
box -8 -3 16 105
use FILL  FILL_1460
timestamp 1713400504
transform 1 0 2824 0 1 1970
box -8 -3 16 105
use FILL  FILL_1461
timestamp 1713400504
transform 1 0 2792 0 1 1970
box -8 -3 16 105
use FILL  FILL_1462
timestamp 1713400504
transform 1 0 2784 0 1 1970
box -8 -3 16 105
use FILL  FILL_1463
timestamp 1713400504
transform 1 0 2776 0 1 1970
box -8 -3 16 105
use FILL  FILL_1464
timestamp 1713400504
transform 1 0 2768 0 1 1970
box -8 -3 16 105
use FILL  FILL_1465
timestamp 1713400504
transform 1 0 2728 0 1 1970
box -8 -3 16 105
use FILL  FILL_1466
timestamp 1713400504
transform 1 0 2720 0 1 1970
box -8 -3 16 105
use FILL  FILL_1467
timestamp 1713400504
transform 1 0 2712 0 1 1970
box -8 -3 16 105
use FILL  FILL_1468
timestamp 1713400504
transform 1 0 2608 0 1 1970
box -8 -3 16 105
use FILL  FILL_1469
timestamp 1713400504
transform 1 0 2600 0 1 1970
box -8 -3 16 105
use FILL  FILL_1470
timestamp 1713400504
transform 1 0 2592 0 1 1970
box -8 -3 16 105
use FILL  FILL_1471
timestamp 1713400504
transform 1 0 2568 0 1 1970
box -8 -3 16 105
use FILL  FILL_1472
timestamp 1713400504
transform 1 0 2536 0 1 1970
box -8 -3 16 105
use FILL  FILL_1473
timestamp 1713400504
transform 1 0 2528 0 1 1970
box -8 -3 16 105
use FILL  FILL_1474
timestamp 1713400504
transform 1 0 2520 0 1 1970
box -8 -3 16 105
use FILL  FILL_1475
timestamp 1713400504
transform 1 0 2512 0 1 1970
box -8 -3 16 105
use FILL  FILL_1476
timestamp 1713400504
transform 1 0 2488 0 1 1970
box -8 -3 16 105
use FILL  FILL_1477
timestamp 1713400504
transform 1 0 2480 0 1 1970
box -8 -3 16 105
use FILL  FILL_1478
timestamp 1713400504
transform 1 0 2472 0 1 1970
box -8 -3 16 105
use FILL  FILL_1479
timestamp 1713400504
transform 1 0 2464 0 1 1970
box -8 -3 16 105
use FILL  FILL_1480
timestamp 1713400504
transform 1 0 2456 0 1 1970
box -8 -3 16 105
use FILL  FILL_1481
timestamp 1713400504
transform 1 0 2416 0 1 1970
box -8 -3 16 105
use FILL  FILL_1482
timestamp 1713400504
transform 1 0 2408 0 1 1970
box -8 -3 16 105
use FILL  FILL_1483
timestamp 1713400504
transform 1 0 2400 0 1 1970
box -8 -3 16 105
use FILL  FILL_1484
timestamp 1713400504
transform 1 0 2392 0 1 1970
box -8 -3 16 105
use FILL  FILL_1485
timestamp 1713400504
transform 1 0 2384 0 1 1970
box -8 -3 16 105
use FILL  FILL_1486
timestamp 1713400504
transform 1 0 2376 0 1 1970
box -8 -3 16 105
use FILL  FILL_1487
timestamp 1713400504
transform 1 0 2368 0 1 1970
box -8 -3 16 105
use FILL  FILL_1488
timestamp 1713400504
transform 1 0 2336 0 1 1970
box -8 -3 16 105
use FILL  FILL_1489
timestamp 1713400504
transform 1 0 2328 0 1 1970
box -8 -3 16 105
use FILL  FILL_1490
timestamp 1713400504
transform 1 0 2320 0 1 1970
box -8 -3 16 105
use FILL  FILL_1491
timestamp 1713400504
transform 1 0 2312 0 1 1970
box -8 -3 16 105
use FILL  FILL_1492
timestamp 1713400504
transform 1 0 2304 0 1 1970
box -8 -3 16 105
use FILL  FILL_1493
timestamp 1713400504
transform 1 0 2272 0 1 1970
box -8 -3 16 105
use FILL  FILL_1494
timestamp 1713400504
transform 1 0 2264 0 1 1970
box -8 -3 16 105
use FILL  FILL_1495
timestamp 1713400504
transform 1 0 2256 0 1 1970
box -8 -3 16 105
use FILL  FILL_1496
timestamp 1713400504
transform 1 0 2248 0 1 1970
box -8 -3 16 105
use FILL  FILL_1497
timestamp 1713400504
transform 1 0 2240 0 1 1970
box -8 -3 16 105
use FILL  FILL_1498
timestamp 1713400504
transform 1 0 2232 0 1 1970
box -8 -3 16 105
use FILL  FILL_1499
timestamp 1713400504
transform 1 0 2224 0 1 1970
box -8 -3 16 105
use FILL  FILL_1500
timestamp 1713400504
transform 1 0 2192 0 1 1970
box -8 -3 16 105
use FILL  FILL_1501
timestamp 1713400504
transform 1 0 2184 0 1 1970
box -8 -3 16 105
use FILL  FILL_1502
timestamp 1713400504
transform 1 0 2176 0 1 1970
box -8 -3 16 105
use FILL  FILL_1503
timestamp 1713400504
transform 1 0 2168 0 1 1970
box -8 -3 16 105
use FILL  FILL_1504
timestamp 1713400504
transform 1 0 2160 0 1 1970
box -8 -3 16 105
use FILL  FILL_1505
timestamp 1713400504
transform 1 0 2152 0 1 1970
box -8 -3 16 105
use FILL  FILL_1506
timestamp 1713400504
transform 1 0 2120 0 1 1970
box -8 -3 16 105
use FILL  FILL_1507
timestamp 1713400504
transform 1 0 2112 0 1 1970
box -8 -3 16 105
use FILL  FILL_1508
timestamp 1713400504
transform 1 0 2104 0 1 1970
box -8 -3 16 105
use FILL  FILL_1509
timestamp 1713400504
transform 1 0 2096 0 1 1970
box -8 -3 16 105
use FILL  FILL_1510
timestamp 1713400504
transform 1 0 2088 0 1 1970
box -8 -3 16 105
use FILL  FILL_1511
timestamp 1713400504
transform 1 0 2080 0 1 1970
box -8 -3 16 105
use FILL  FILL_1512
timestamp 1713400504
transform 1 0 2072 0 1 1970
box -8 -3 16 105
use FILL  FILL_1513
timestamp 1713400504
transform 1 0 2064 0 1 1970
box -8 -3 16 105
use FILL  FILL_1514
timestamp 1713400504
transform 1 0 2056 0 1 1970
box -8 -3 16 105
use FILL  FILL_1515
timestamp 1713400504
transform 1 0 2016 0 1 1970
box -8 -3 16 105
use FILL  FILL_1516
timestamp 1713400504
transform 1 0 2008 0 1 1970
box -8 -3 16 105
use FILL  FILL_1517
timestamp 1713400504
transform 1 0 2000 0 1 1970
box -8 -3 16 105
use FILL  FILL_1518
timestamp 1713400504
transform 1 0 1992 0 1 1970
box -8 -3 16 105
use FILL  FILL_1519
timestamp 1713400504
transform 1 0 1984 0 1 1970
box -8 -3 16 105
use FILL  FILL_1520
timestamp 1713400504
transform 1 0 1976 0 1 1970
box -8 -3 16 105
use FILL  FILL_1521
timestamp 1713400504
transform 1 0 1944 0 1 1970
box -8 -3 16 105
use FILL  FILL_1522
timestamp 1713400504
transform 1 0 1936 0 1 1970
box -8 -3 16 105
use FILL  FILL_1523
timestamp 1713400504
transform 1 0 1928 0 1 1970
box -8 -3 16 105
use FILL  FILL_1524
timestamp 1713400504
transform 1 0 1920 0 1 1970
box -8 -3 16 105
use FILL  FILL_1525
timestamp 1713400504
transform 1 0 1912 0 1 1970
box -8 -3 16 105
use FILL  FILL_1526
timestamp 1713400504
transform 1 0 1872 0 1 1970
box -8 -3 16 105
use FILL  FILL_1527
timestamp 1713400504
transform 1 0 1864 0 1 1970
box -8 -3 16 105
use FILL  FILL_1528
timestamp 1713400504
transform 1 0 1856 0 1 1970
box -8 -3 16 105
use FILL  FILL_1529
timestamp 1713400504
transform 1 0 1848 0 1 1970
box -8 -3 16 105
use FILL  FILL_1530
timestamp 1713400504
transform 1 0 1840 0 1 1970
box -8 -3 16 105
use FILL  FILL_1531
timestamp 1713400504
transform 1 0 1808 0 1 1970
box -8 -3 16 105
use FILL  FILL_1532
timestamp 1713400504
transform 1 0 1800 0 1 1970
box -8 -3 16 105
use FILL  FILL_1533
timestamp 1713400504
transform 1 0 1792 0 1 1970
box -8 -3 16 105
use FILL  FILL_1534
timestamp 1713400504
transform 1 0 1784 0 1 1970
box -8 -3 16 105
use FILL  FILL_1535
timestamp 1713400504
transform 1 0 1776 0 1 1970
box -8 -3 16 105
use FILL  FILL_1536
timestamp 1713400504
transform 1 0 1768 0 1 1970
box -8 -3 16 105
use FILL  FILL_1537
timestamp 1713400504
transform 1 0 1760 0 1 1970
box -8 -3 16 105
use FILL  FILL_1538
timestamp 1713400504
transform 1 0 1712 0 1 1970
box -8 -3 16 105
use FILL  FILL_1539
timestamp 1713400504
transform 1 0 1704 0 1 1970
box -8 -3 16 105
use FILL  FILL_1540
timestamp 1713400504
transform 1 0 1696 0 1 1970
box -8 -3 16 105
use FILL  FILL_1541
timestamp 1713400504
transform 1 0 1688 0 1 1970
box -8 -3 16 105
use FILL  FILL_1542
timestamp 1713400504
transform 1 0 1680 0 1 1970
box -8 -3 16 105
use FILL  FILL_1543
timestamp 1713400504
transform 1 0 1672 0 1 1970
box -8 -3 16 105
use FILL  FILL_1544
timestamp 1713400504
transform 1 0 1664 0 1 1970
box -8 -3 16 105
use FILL  FILL_1545
timestamp 1713400504
transform 1 0 1656 0 1 1970
box -8 -3 16 105
use FILL  FILL_1546
timestamp 1713400504
transform 1 0 1608 0 1 1970
box -8 -3 16 105
use FILL  FILL_1547
timestamp 1713400504
transform 1 0 1600 0 1 1970
box -8 -3 16 105
use FILL  FILL_1548
timestamp 1713400504
transform 1 0 1592 0 1 1970
box -8 -3 16 105
use FILL  FILL_1549
timestamp 1713400504
transform 1 0 1584 0 1 1970
box -8 -3 16 105
use FILL  FILL_1550
timestamp 1713400504
transform 1 0 1576 0 1 1970
box -8 -3 16 105
use FILL  FILL_1551
timestamp 1713400504
transform 1 0 1568 0 1 1970
box -8 -3 16 105
use FILL  FILL_1552
timestamp 1713400504
transform 1 0 1560 0 1 1970
box -8 -3 16 105
use FILL  FILL_1553
timestamp 1713400504
transform 1 0 1552 0 1 1970
box -8 -3 16 105
use FILL  FILL_1554
timestamp 1713400504
transform 1 0 1512 0 1 1970
box -8 -3 16 105
use FILL  FILL_1555
timestamp 1713400504
transform 1 0 1504 0 1 1970
box -8 -3 16 105
use FILL  FILL_1556
timestamp 1713400504
transform 1 0 1496 0 1 1970
box -8 -3 16 105
use FILL  FILL_1557
timestamp 1713400504
transform 1 0 1488 0 1 1970
box -8 -3 16 105
use FILL  FILL_1558
timestamp 1713400504
transform 1 0 1480 0 1 1970
box -8 -3 16 105
use FILL  FILL_1559
timestamp 1713400504
transform 1 0 1440 0 1 1970
box -8 -3 16 105
use FILL  FILL_1560
timestamp 1713400504
transform 1 0 1432 0 1 1970
box -8 -3 16 105
use FILL  FILL_1561
timestamp 1713400504
transform 1 0 1424 0 1 1970
box -8 -3 16 105
use FILL  FILL_1562
timestamp 1713400504
transform 1 0 1416 0 1 1970
box -8 -3 16 105
use FILL  FILL_1563
timestamp 1713400504
transform 1 0 1408 0 1 1970
box -8 -3 16 105
use FILL  FILL_1564
timestamp 1713400504
transform 1 0 1400 0 1 1970
box -8 -3 16 105
use FILL  FILL_1565
timestamp 1713400504
transform 1 0 1360 0 1 1970
box -8 -3 16 105
use FILL  FILL_1566
timestamp 1713400504
transform 1 0 1352 0 1 1970
box -8 -3 16 105
use FILL  FILL_1567
timestamp 1713400504
transform 1 0 1344 0 1 1970
box -8 -3 16 105
use FILL  FILL_1568
timestamp 1713400504
transform 1 0 1336 0 1 1970
box -8 -3 16 105
use FILL  FILL_1569
timestamp 1713400504
transform 1 0 1272 0 1 1970
box -8 -3 16 105
use FILL  FILL_1570
timestamp 1713400504
transform 1 0 1264 0 1 1970
box -8 -3 16 105
use FILL  FILL_1571
timestamp 1713400504
transform 1 0 1256 0 1 1970
box -8 -3 16 105
use FILL  FILL_1572
timestamp 1713400504
transform 1 0 1248 0 1 1970
box -8 -3 16 105
use FILL  FILL_1573
timestamp 1713400504
transform 1 0 1208 0 1 1970
box -8 -3 16 105
use FILL  FILL_1574
timestamp 1713400504
transform 1 0 1200 0 1 1970
box -8 -3 16 105
use FILL  FILL_1575
timestamp 1713400504
transform 1 0 1192 0 1 1970
box -8 -3 16 105
use FILL  FILL_1576
timestamp 1713400504
transform 1 0 1184 0 1 1970
box -8 -3 16 105
use FILL  FILL_1577
timestamp 1713400504
transform 1 0 1176 0 1 1970
box -8 -3 16 105
use FILL  FILL_1578
timestamp 1713400504
transform 1 0 1168 0 1 1970
box -8 -3 16 105
use FILL  FILL_1579
timestamp 1713400504
transform 1 0 1160 0 1 1970
box -8 -3 16 105
use FILL  FILL_1580
timestamp 1713400504
transform 1 0 1128 0 1 1970
box -8 -3 16 105
use FILL  FILL_1581
timestamp 1713400504
transform 1 0 1120 0 1 1970
box -8 -3 16 105
use FILL  FILL_1582
timestamp 1713400504
transform 1 0 1112 0 1 1970
box -8 -3 16 105
use FILL  FILL_1583
timestamp 1713400504
transform 1 0 1088 0 1 1970
box -8 -3 16 105
use FILL  FILL_1584
timestamp 1713400504
transform 1 0 1080 0 1 1970
box -8 -3 16 105
use FILL  FILL_1585
timestamp 1713400504
transform 1 0 1072 0 1 1970
box -8 -3 16 105
use FILL  FILL_1586
timestamp 1713400504
transform 1 0 1064 0 1 1970
box -8 -3 16 105
use FILL  FILL_1587
timestamp 1713400504
transform 1 0 1056 0 1 1970
box -8 -3 16 105
use FILL  FILL_1588
timestamp 1713400504
transform 1 0 1024 0 1 1970
box -8 -3 16 105
use FILL  FILL_1589
timestamp 1713400504
transform 1 0 1016 0 1 1970
box -8 -3 16 105
use FILL  FILL_1590
timestamp 1713400504
transform 1 0 1008 0 1 1970
box -8 -3 16 105
use FILL  FILL_1591
timestamp 1713400504
transform 1 0 1000 0 1 1970
box -8 -3 16 105
use FILL  FILL_1592
timestamp 1713400504
transform 1 0 992 0 1 1970
box -8 -3 16 105
use FILL  FILL_1593
timestamp 1713400504
transform 1 0 984 0 1 1970
box -8 -3 16 105
use FILL  FILL_1594
timestamp 1713400504
transform 1 0 976 0 1 1970
box -8 -3 16 105
use FILL  FILL_1595
timestamp 1713400504
transform 1 0 928 0 1 1970
box -8 -3 16 105
use FILL  FILL_1596
timestamp 1713400504
transform 1 0 920 0 1 1970
box -8 -3 16 105
use FILL  FILL_1597
timestamp 1713400504
transform 1 0 912 0 1 1970
box -8 -3 16 105
use FILL  FILL_1598
timestamp 1713400504
transform 1 0 904 0 1 1970
box -8 -3 16 105
use FILL  FILL_1599
timestamp 1713400504
transform 1 0 896 0 1 1970
box -8 -3 16 105
use FILL  FILL_1600
timestamp 1713400504
transform 1 0 888 0 1 1970
box -8 -3 16 105
use FILL  FILL_1601
timestamp 1713400504
transform 1 0 880 0 1 1970
box -8 -3 16 105
use FILL  FILL_1602
timestamp 1713400504
transform 1 0 872 0 1 1970
box -8 -3 16 105
use FILL  FILL_1603
timestamp 1713400504
transform 1 0 864 0 1 1970
box -8 -3 16 105
use FILL  FILL_1604
timestamp 1713400504
transform 1 0 824 0 1 1970
box -8 -3 16 105
use FILL  FILL_1605
timestamp 1713400504
transform 1 0 816 0 1 1970
box -8 -3 16 105
use FILL  FILL_1606
timestamp 1713400504
transform 1 0 808 0 1 1970
box -8 -3 16 105
use FILL  FILL_1607
timestamp 1713400504
transform 1 0 800 0 1 1970
box -8 -3 16 105
use FILL  FILL_1608
timestamp 1713400504
transform 1 0 792 0 1 1970
box -8 -3 16 105
use FILL  FILL_1609
timestamp 1713400504
transform 1 0 784 0 1 1970
box -8 -3 16 105
use FILL  FILL_1610
timestamp 1713400504
transform 1 0 776 0 1 1970
box -8 -3 16 105
use FILL  FILL_1611
timestamp 1713400504
transform 1 0 768 0 1 1970
box -8 -3 16 105
use FILL  FILL_1612
timestamp 1713400504
transform 1 0 760 0 1 1970
box -8 -3 16 105
use FILL  FILL_1613
timestamp 1713400504
transform 1 0 712 0 1 1970
box -8 -3 16 105
use FILL  FILL_1614
timestamp 1713400504
transform 1 0 704 0 1 1970
box -8 -3 16 105
use FILL  FILL_1615
timestamp 1713400504
transform 1 0 696 0 1 1970
box -8 -3 16 105
use FILL  FILL_1616
timestamp 1713400504
transform 1 0 688 0 1 1970
box -8 -3 16 105
use FILL  FILL_1617
timestamp 1713400504
transform 1 0 680 0 1 1970
box -8 -3 16 105
use FILL  FILL_1618
timestamp 1713400504
transform 1 0 672 0 1 1970
box -8 -3 16 105
use FILL  FILL_1619
timestamp 1713400504
transform 1 0 664 0 1 1970
box -8 -3 16 105
use FILL  FILL_1620
timestamp 1713400504
transform 1 0 632 0 1 1970
box -8 -3 16 105
use FILL  FILL_1621
timestamp 1713400504
transform 1 0 624 0 1 1970
box -8 -3 16 105
use FILL  FILL_1622
timestamp 1713400504
transform 1 0 616 0 1 1970
box -8 -3 16 105
use FILL  FILL_1623
timestamp 1713400504
transform 1 0 608 0 1 1970
box -8 -3 16 105
use FILL  FILL_1624
timestamp 1713400504
transform 1 0 600 0 1 1970
box -8 -3 16 105
use FILL  FILL_1625
timestamp 1713400504
transform 1 0 568 0 1 1970
box -8 -3 16 105
use FILL  FILL_1626
timestamp 1713400504
transform 1 0 560 0 1 1970
box -8 -3 16 105
use FILL  FILL_1627
timestamp 1713400504
transform 1 0 552 0 1 1970
box -8 -3 16 105
use FILL  FILL_1628
timestamp 1713400504
transform 1 0 544 0 1 1970
box -8 -3 16 105
use FILL  FILL_1629
timestamp 1713400504
transform 1 0 536 0 1 1970
box -8 -3 16 105
use FILL  FILL_1630
timestamp 1713400504
transform 1 0 528 0 1 1970
box -8 -3 16 105
use FILL  FILL_1631
timestamp 1713400504
transform 1 0 496 0 1 1970
box -8 -3 16 105
use FILL  FILL_1632
timestamp 1713400504
transform 1 0 488 0 1 1970
box -8 -3 16 105
use FILL  FILL_1633
timestamp 1713400504
transform 1 0 480 0 1 1970
box -8 -3 16 105
use FILL  FILL_1634
timestamp 1713400504
transform 1 0 472 0 1 1970
box -8 -3 16 105
use FILL  FILL_1635
timestamp 1713400504
transform 1 0 440 0 1 1970
box -8 -3 16 105
use FILL  FILL_1636
timestamp 1713400504
transform 1 0 432 0 1 1970
box -8 -3 16 105
use FILL  FILL_1637
timestamp 1713400504
transform 1 0 424 0 1 1970
box -8 -3 16 105
use FILL  FILL_1638
timestamp 1713400504
transform 1 0 416 0 1 1970
box -8 -3 16 105
use FILL  FILL_1639
timestamp 1713400504
transform 1 0 408 0 1 1970
box -8 -3 16 105
use FILL  FILL_1640
timestamp 1713400504
transform 1 0 400 0 1 1970
box -8 -3 16 105
use FILL  FILL_1641
timestamp 1713400504
transform 1 0 368 0 1 1970
box -8 -3 16 105
use FILL  FILL_1642
timestamp 1713400504
transform 1 0 360 0 1 1970
box -8 -3 16 105
use FILL  FILL_1643
timestamp 1713400504
transform 1 0 352 0 1 1970
box -8 -3 16 105
use FILL  FILL_1644
timestamp 1713400504
transform 1 0 344 0 1 1970
box -8 -3 16 105
use FILL  FILL_1645
timestamp 1713400504
transform 1 0 336 0 1 1970
box -8 -3 16 105
use FILL  FILL_1646
timestamp 1713400504
transform 1 0 312 0 1 1970
box -8 -3 16 105
use FILL  FILL_1647
timestamp 1713400504
transform 1 0 304 0 1 1970
box -8 -3 16 105
use FILL  FILL_1648
timestamp 1713400504
transform 1 0 264 0 1 1970
box -8 -3 16 105
use FILL  FILL_1649
timestamp 1713400504
transform 1 0 256 0 1 1970
box -8 -3 16 105
use FILL  FILL_1650
timestamp 1713400504
transform 1 0 248 0 1 1970
box -8 -3 16 105
use FILL  FILL_1651
timestamp 1713400504
transform 1 0 240 0 1 1970
box -8 -3 16 105
use FILL  FILL_1652
timestamp 1713400504
transform 1 0 232 0 1 1970
box -8 -3 16 105
use FILL  FILL_1653
timestamp 1713400504
transform 1 0 176 0 1 1970
box -8 -3 16 105
use FILL  FILL_1654
timestamp 1713400504
transform 1 0 168 0 1 1970
box -8 -3 16 105
use FILL  FILL_1655
timestamp 1713400504
transform 1 0 160 0 1 1970
box -8 -3 16 105
use FILL  FILL_1656
timestamp 1713400504
transform 1 0 72 0 1 1970
box -8 -3 16 105
use FILL  FILL_1657
timestamp 1713400504
transform 1 0 3008 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1658
timestamp 1713400504
transform 1 0 3000 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1659
timestamp 1713400504
transform 1 0 2992 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1660
timestamp 1713400504
transform 1 0 2984 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1661
timestamp 1713400504
transform 1 0 2976 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1662
timestamp 1713400504
transform 1 0 2968 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1663
timestamp 1713400504
transform 1 0 2944 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1664
timestamp 1713400504
transform 1 0 2936 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1665
timestamp 1713400504
transform 1 0 2928 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1666
timestamp 1713400504
transform 1 0 2888 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1667
timestamp 1713400504
transform 1 0 2880 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1668
timestamp 1713400504
transform 1 0 2872 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1669
timestamp 1713400504
transform 1 0 2864 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1670
timestamp 1713400504
transform 1 0 2760 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1671
timestamp 1713400504
transform 1 0 2752 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1672
timestamp 1713400504
transform 1 0 2712 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1673
timestamp 1713400504
transform 1 0 2704 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1674
timestamp 1713400504
transform 1 0 2696 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1675
timestamp 1713400504
transform 1 0 2688 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1676
timestamp 1713400504
transform 1 0 2680 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1677
timestamp 1713400504
transform 1 0 2672 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1678
timestamp 1713400504
transform 1 0 2624 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1679
timestamp 1713400504
transform 1 0 2616 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1680
timestamp 1713400504
transform 1 0 2608 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1681
timestamp 1713400504
transform 1 0 2600 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1682
timestamp 1713400504
transform 1 0 2592 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1683
timestamp 1713400504
transform 1 0 2552 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1684
timestamp 1713400504
transform 1 0 2544 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1685
timestamp 1713400504
transform 1 0 2536 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1686
timestamp 1713400504
transform 1 0 2528 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1687
timestamp 1713400504
transform 1 0 2488 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1688
timestamp 1713400504
transform 1 0 2480 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1689
timestamp 1713400504
transform 1 0 2472 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1690
timestamp 1713400504
transform 1 0 2464 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1691
timestamp 1713400504
transform 1 0 2432 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1692
timestamp 1713400504
transform 1 0 2424 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1693
timestamp 1713400504
transform 1 0 2416 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1694
timestamp 1713400504
transform 1 0 2384 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1695
timestamp 1713400504
transform 1 0 2376 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1696
timestamp 1713400504
transform 1 0 2368 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1697
timestamp 1713400504
transform 1 0 2360 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1698
timestamp 1713400504
transform 1 0 2352 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1699
timestamp 1713400504
transform 1 0 2320 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1700
timestamp 1713400504
transform 1 0 2312 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1701
timestamp 1713400504
transform 1 0 2304 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1702
timestamp 1713400504
transform 1 0 2272 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1703
timestamp 1713400504
transform 1 0 2264 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1704
timestamp 1713400504
transform 1 0 2256 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1705
timestamp 1713400504
transform 1 0 2248 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1706
timestamp 1713400504
transform 1 0 2144 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1707
timestamp 1713400504
transform 1 0 2136 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1708
timestamp 1713400504
transform 1 0 2128 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1709
timestamp 1713400504
transform 1 0 2120 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1710
timestamp 1713400504
transform 1 0 2072 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1711
timestamp 1713400504
transform 1 0 2064 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1712
timestamp 1713400504
transform 1 0 2056 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1713
timestamp 1713400504
transform 1 0 2048 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1714
timestamp 1713400504
transform 1 0 2040 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1715
timestamp 1713400504
transform 1 0 2032 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1716
timestamp 1713400504
transform 1 0 2024 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1717
timestamp 1713400504
transform 1 0 1984 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1718
timestamp 1713400504
transform 1 0 1976 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1719
timestamp 1713400504
transform 1 0 1968 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1720
timestamp 1713400504
transform 1 0 1960 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1721
timestamp 1713400504
transform 1 0 1952 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1722
timestamp 1713400504
transform 1 0 1944 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1723
timestamp 1713400504
transform 1 0 1912 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1724
timestamp 1713400504
transform 1 0 1904 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1725
timestamp 1713400504
transform 1 0 1896 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1726
timestamp 1713400504
transform 1 0 1888 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1727
timestamp 1713400504
transform 1 0 1864 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1728
timestamp 1713400504
transform 1 0 1856 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1729
timestamp 1713400504
transform 1 0 1848 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1730
timestamp 1713400504
transform 1 0 1816 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1731
timestamp 1713400504
transform 1 0 1808 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1732
timestamp 1713400504
transform 1 0 1800 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1733
timestamp 1713400504
transform 1 0 1792 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1734
timestamp 1713400504
transform 1 0 1784 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1735
timestamp 1713400504
transform 1 0 1776 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1736
timestamp 1713400504
transform 1 0 1728 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1737
timestamp 1713400504
transform 1 0 1720 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1738
timestamp 1713400504
transform 1 0 1712 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1739
timestamp 1713400504
transform 1 0 1704 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1740
timestamp 1713400504
transform 1 0 1696 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1741
timestamp 1713400504
transform 1 0 1688 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1742
timestamp 1713400504
transform 1 0 1680 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1743
timestamp 1713400504
transform 1 0 1672 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1744
timestamp 1713400504
transform 1 0 1632 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1745
timestamp 1713400504
transform 1 0 1624 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1746
timestamp 1713400504
transform 1 0 1616 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1747
timestamp 1713400504
transform 1 0 1608 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1748
timestamp 1713400504
transform 1 0 1600 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1749
timestamp 1713400504
transform 1 0 1576 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1750
timestamp 1713400504
transform 1 0 1568 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1751
timestamp 1713400504
transform 1 0 1560 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1752
timestamp 1713400504
transform 1 0 1552 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1753
timestamp 1713400504
transform 1 0 1544 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1754
timestamp 1713400504
transform 1 0 1496 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1755
timestamp 1713400504
transform 1 0 1488 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1756
timestamp 1713400504
transform 1 0 1480 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1757
timestamp 1713400504
transform 1 0 1472 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1758
timestamp 1713400504
transform 1 0 1464 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1759
timestamp 1713400504
transform 1 0 1456 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1760
timestamp 1713400504
transform 1 0 1432 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1761
timestamp 1713400504
transform 1 0 1424 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1762
timestamp 1713400504
transform 1 0 1416 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1763
timestamp 1713400504
transform 1 0 1352 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1764
timestamp 1713400504
transform 1 0 1344 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1765
timestamp 1713400504
transform 1 0 1336 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1766
timestamp 1713400504
transform 1 0 1304 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1767
timestamp 1713400504
transform 1 0 1296 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1768
timestamp 1713400504
transform 1 0 1288 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1769
timestamp 1713400504
transform 1 0 1280 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1770
timestamp 1713400504
transform 1 0 1272 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1771
timestamp 1713400504
transform 1 0 1264 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1772
timestamp 1713400504
transform 1 0 1232 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1773
timestamp 1713400504
transform 1 0 1224 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1774
timestamp 1713400504
transform 1 0 1216 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1775
timestamp 1713400504
transform 1 0 1208 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1776
timestamp 1713400504
transform 1 0 1176 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1777
timestamp 1713400504
transform 1 0 1168 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1778
timestamp 1713400504
transform 1 0 1160 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1779
timestamp 1713400504
transform 1 0 1152 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1780
timestamp 1713400504
transform 1 0 1144 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1781
timestamp 1713400504
transform 1 0 1136 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1782
timestamp 1713400504
transform 1 0 1128 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1783
timestamp 1713400504
transform 1 0 1088 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1784
timestamp 1713400504
transform 1 0 1080 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1785
timestamp 1713400504
transform 1 0 1072 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1786
timestamp 1713400504
transform 1 0 1064 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1787
timestamp 1713400504
transform 1 0 1056 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1788
timestamp 1713400504
transform 1 0 1048 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1789
timestamp 1713400504
transform 1 0 1040 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1790
timestamp 1713400504
transform 1 0 1008 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1791
timestamp 1713400504
transform 1 0 1000 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1792
timestamp 1713400504
transform 1 0 992 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1793
timestamp 1713400504
transform 1 0 984 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1794
timestamp 1713400504
transform 1 0 976 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1795
timestamp 1713400504
transform 1 0 968 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1796
timestamp 1713400504
transform 1 0 936 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1797
timestamp 1713400504
transform 1 0 928 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1798
timestamp 1713400504
transform 1 0 920 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1799
timestamp 1713400504
transform 1 0 912 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1800
timestamp 1713400504
transform 1 0 904 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1801
timestamp 1713400504
transform 1 0 896 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1802
timestamp 1713400504
transform 1 0 888 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1803
timestamp 1713400504
transform 1 0 880 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1804
timestamp 1713400504
transform 1 0 832 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1805
timestamp 1713400504
transform 1 0 824 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1806
timestamp 1713400504
transform 1 0 816 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1807
timestamp 1713400504
transform 1 0 808 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1808
timestamp 1713400504
transform 1 0 800 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1809
timestamp 1713400504
transform 1 0 792 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1810
timestamp 1713400504
transform 1 0 784 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1811
timestamp 1713400504
transform 1 0 776 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1812
timestamp 1713400504
transform 1 0 768 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1813
timestamp 1713400504
transform 1 0 720 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1814
timestamp 1713400504
transform 1 0 712 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1815
timestamp 1713400504
transform 1 0 704 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1816
timestamp 1713400504
transform 1 0 696 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1817
timestamp 1713400504
transform 1 0 688 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1818
timestamp 1713400504
transform 1 0 680 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1819
timestamp 1713400504
transform 1 0 672 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1820
timestamp 1713400504
transform 1 0 664 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1821
timestamp 1713400504
transform 1 0 656 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1822
timestamp 1713400504
transform 1 0 648 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1823
timestamp 1713400504
transform 1 0 640 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1824
timestamp 1713400504
transform 1 0 632 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1825
timestamp 1713400504
transform 1 0 624 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1826
timestamp 1713400504
transform 1 0 616 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1827
timestamp 1713400504
transform 1 0 608 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1828
timestamp 1713400504
transform 1 0 600 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1829
timestamp 1713400504
transform 1 0 592 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1830
timestamp 1713400504
transform 1 0 584 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1831
timestamp 1713400504
transform 1 0 576 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1832
timestamp 1713400504
transform 1 0 568 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1833
timestamp 1713400504
transform 1 0 544 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1834
timestamp 1713400504
transform 1 0 536 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1835
timestamp 1713400504
transform 1 0 528 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1836
timestamp 1713400504
transform 1 0 520 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1837
timestamp 1713400504
transform 1 0 512 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1838
timestamp 1713400504
transform 1 0 504 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1839
timestamp 1713400504
transform 1 0 480 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1840
timestamp 1713400504
transform 1 0 472 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1841
timestamp 1713400504
transform 1 0 464 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1842
timestamp 1713400504
transform 1 0 456 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1843
timestamp 1713400504
transform 1 0 448 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1844
timestamp 1713400504
transform 1 0 424 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1845
timestamp 1713400504
transform 1 0 416 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1846
timestamp 1713400504
transform 1 0 408 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1847
timestamp 1713400504
transform 1 0 400 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1848
timestamp 1713400504
transform 1 0 376 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1849
timestamp 1713400504
transform 1 0 368 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1850
timestamp 1713400504
transform 1 0 360 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1851
timestamp 1713400504
transform 1 0 352 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1852
timestamp 1713400504
transform 1 0 288 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1853
timestamp 1713400504
transform 1 0 280 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1854
timestamp 1713400504
transform 1 0 272 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1855
timestamp 1713400504
transform 1 0 264 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1856
timestamp 1713400504
transform 1 0 256 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1857
timestamp 1713400504
transform 1 0 224 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1858
timestamp 1713400504
transform 1 0 216 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1859
timestamp 1713400504
transform 1 0 208 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1860
timestamp 1713400504
transform 1 0 144 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1861
timestamp 1713400504
transform 1 0 136 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1862
timestamp 1713400504
transform 1 0 128 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1863
timestamp 1713400504
transform 1 0 120 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1864
timestamp 1713400504
transform 1 0 88 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1865
timestamp 1713400504
transform 1 0 80 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1866
timestamp 1713400504
transform 1 0 72 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1867
timestamp 1713400504
transform 1 0 3008 0 1 1770
box -8 -3 16 105
use FILL  FILL_1868
timestamp 1713400504
transform 1 0 3000 0 1 1770
box -8 -3 16 105
use FILL  FILL_1869
timestamp 1713400504
transform 1 0 2976 0 1 1770
box -8 -3 16 105
use FILL  FILL_1870
timestamp 1713400504
transform 1 0 2968 0 1 1770
box -8 -3 16 105
use FILL  FILL_1871
timestamp 1713400504
transform 1 0 2960 0 1 1770
box -8 -3 16 105
use FILL  FILL_1872
timestamp 1713400504
transform 1 0 2912 0 1 1770
box -8 -3 16 105
use FILL  FILL_1873
timestamp 1713400504
transform 1 0 2904 0 1 1770
box -8 -3 16 105
use FILL  FILL_1874
timestamp 1713400504
transform 1 0 2896 0 1 1770
box -8 -3 16 105
use FILL  FILL_1875
timestamp 1713400504
transform 1 0 2888 0 1 1770
box -8 -3 16 105
use FILL  FILL_1876
timestamp 1713400504
transform 1 0 2880 0 1 1770
box -8 -3 16 105
use FILL  FILL_1877
timestamp 1713400504
transform 1 0 2872 0 1 1770
box -8 -3 16 105
use FILL  FILL_1878
timestamp 1713400504
transform 1 0 2824 0 1 1770
box -8 -3 16 105
use FILL  FILL_1879
timestamp 1713400504
transform 1 0 2816 0 1 1770
box -8 -3 16 105
use FILL  FILL_1880
timestamp 1713400504
transform 1 0 2808 0 1 1770
box -8 -3 16 105
use FILL  FILL_1881
timestamp 1713400504
transform 1 0 2800 0 1 1770
box -8 -3 16 105
use FILL  FILL_1882
timestamp 1713400504
transform 1 0 2792 0 1 1770
box -8 -3 16 105
use FILL  FILL_1883
timestamp 1713400504
transform 1 0 2784 0 1 1770
box -8 -3 16 105
use FILL  FILL_1884
timestamp 1713400504
transform 1 0 2736 0 1 1770
box -8 -3 16 105
use FILL  FILL_1885
timestamp 1713400504
transform 1 0 2728 0 1 1770
box -8 -3 16 105
use FILL  FILL_1886
timestamp 1713400504
transform 1 0 2720 0 1 1770
box -8 -3 16 105
use FILL  FILL_1887
timestamp 1713400504
transform 1 0 2712 0 1 1770
box -8 -3 16 105
use FILL  FILL_1888
timestamp 1713400504
transform 1 0 2704 0 1 1770
box -8 -3 16 105
use FILL  FILL_1889
timestamp 1713400504
transform 1 0 2664 0 1 1770
box -8 -3 16 105
use FILL  FILL_1890
timestamp 1713400504
transform 1 0 2656 0 1 1770
box -8 -3 16 105
use FILL  FILL_1891
timestamp 1713400504
transform 1 0 2648 0 1 1770
box -8 -3 16 105
use FILL  FILL_1892
timestamp 1713400504
transform 1 0 2616 0 1 1770
box -8 -3 16 105
use FILL  FILL_1893
timestamp 1713400504
transform 1 0 2608 0 1 1770
box -8 -3 16 105
use FILL  FILL_1894
timestamp 1713400504
transform 1 0 2600 0 1 1770
box -8 -3 16 105
use FILL  FILL_1895
timestamp 1713400504
transform 1 0 2560 0 1 1770
box -8 -3 16 105
use FILL  FILL_1896
timestamp 1713400504
transform 1 0 2552 0 1 1770
box -8 -3 16 105
use FILL  FILL_1897
timestamp 1713400504
transform 1 0 2544 0 1 1770
box -8 -3 16 105
use FILL  FILL_1898
timestamp 1713400504
transform 1 0 2504 0 1 1770
box -8 -3 16 105
use FILL  FILL_1899
timestamp 1713400504
transform 1 0 2496 0 1 1770
box -8 -3 16 105
use FILL  FILL_1900
timestamp 1713400504
transform 1 0 2392 0 1 1770
box -8 -3 16 105
use FILL  FILL_1901
timestamp 1713400504
transform 1 0 2384 0 1 1770
box -8 -3 16 105
use FILL  FILL_1902
timestamp 1713400504
transform 1 0 2344 0 1 1770
box -8 -3 16 105
use FILL  FILL_1903
timestamp 1713400504
transform 1 0 2336 0 1 1770
box -8 -3 16 105
use FILL  FILL_1904
timestamp 1713400504
transform 1 0 2328 0 1 1770
box -8 -3 16 105
use FILL  FILL_1905
timestamp 1713400504
transform 1 0 2320 0 1 1770
box -8 -3 16 105
use FILL  FILL_1906
timestamp 1713400504
transform 1 0 2288 0 1 1770
box -8 -3 16 105
use FILL  FILL_1907
timestamp 1713400504
transform 1 0 2280 0 1 1770
box -8 -3 16 105
use FILL  FILL_1908
timestamp 1713400504
transform 1 0 2272 0 1 1770
box -8 -3 16 105
use FILL  FILL_1909
timestamp 1713400504
transform 1 0 2240 0 1 1770
box -8 -3 16 105
use FILL  FILL_1910
timestamp 1713400504
transform 1 0 2232 0 1 1770
box -8 -3 16 105
use FILL  FILL_1911
timestamp 1713400504
transform 1 0 2224 0 1 1770
box -8 -3 16 105
use FILL  FILL_1912
timestamp 1713400504
transform 1 0 2192 0 1 1770
box -8 -3 16 105
use FILL  FILL_1913
timestamp 1713400504
transform 1 0 2160 0 1 1770
box -8 -3 16 105
use FILL  FILL_1914
timestamp 1713400504
transform 1 0 2152 0 1 1770
box -8 -3 16 105
use FILL  FILL_1915
timestamp 1713400504
transform 1 0 2144 0 1 1770
box -8 -3 16 105
use FILL  FILL_1916
timestamp 1713400504
transform 1 0 2112 0 1 1770
box -8 -3 16 105
use FILL  FILL_1917
timestamp 1713400504
transform 1 0 2104 0 1 1770
box -8 -3 16 105
use FILL  FILL_1918
timestamp 1713400504
transform 1 0 2096 0 1 1770
box -8 -3 16 105
use FILL  FILL_1919
timestamp 1713400504
transform 1 0 2072 0 1 1770
box -8 -3 16 105
use FILL  FILL_1920
timestamp 1713400504
transform 1 0 2064 0 1 1770
box -8 -3 16 105
use FILL  FILL_1921
timestamp 1713400504
transform 1 0 2056 0 1 1770
box -8 -3 16 105
use FILL  FILL_1922
timestamp 1713400504
transform 1 0 2048 0 1 1770
box -8 -3 16 105
use FILL  FILL_1923
timestamp 1713400504
transform 1 0 2008 0 1 1770
box -8 -3 16 105
use FILL  FILL_1924
timestamp 1713400504
transform 1 0 2000 0 1 1770
box -8 -3 16 105
use FILL  FILL_1925
timestamp 1713400504
transform 1 0 1992 0 1 1770
box -8 -3 16 105
use FILL  FILL_1926
timestamp 1713400504
transform 1 0 1984 0 1 1770
box -8 -3 16 105
use FILL  FILL_1927
timestamp 1713400504
transform 1 0 1944 0 1 1770
box -8 -3 16 105
use FILL  FILL_1928
timestamp 1713400504
transform 1 0 1936 0 1 1770
box -8 -3 16 105
use FILL  FILL_1929
timestamp 1713400504
transform 1 0 1928 0 1 1770
box -8 -3 16 105
use FILL  FILL_1930
timestamp 1713400504
transform 1 0 1920 0 1 1770
box -8 -3 16 105
use FILL  FILL_1931
timestamp 1713400504
transform 1 0 1912 0 1 1770
box -8 -3 16 105
use FILL  FILL_1932
timestamp 1713400504
transform 1 0 1872 0 1 1770
box -8 -3 16 105
use FILL  FILL_1933
timestamp 1713400504
transform 1 0 1864 0 1 1770
box -8 -3 16 105
use FILL  FILL_1934
timestamp 1713400504
transform 1 0 1856 0 1 1770
box -8 -3 16 105
use FILL  FILL_1935
timestamp 1713400504
transform 1 0 1848 0 1 1770
box -8 -3 16 105
use FILL  FILL_1936
timestamp 1713400504
transform 1 0 1808 0 1 1770
box -8 -3 16 105
use FILL  FILL_1937
timestamp 1713400504
transform 1 0 1800 0 1 1770
box -8 -3 16 105
use FILL  FILL_1938
timestamp 1713400504
transform 1 0 1792 0 1 1770
box -8 -3 16 105
use FILL  FILL_1939
timestamp 1713400504
transform 1 0 1768 0 1 1770
box -8 -3 16 105
use FILL  FILL_1940
timestamp 1713400504
transform 1 0 1760 0 1 1770
box -8 -3 16 105
use FILL  FILL_1941
timestamp 1713400504
transform 1 0 1752 0 1 1770
box -8 -3 16 105
use FILL  FILL_1942
timestamp 1713400504
transform 1 0 1744 0 1 1770
box -8 -3 16 105
use FILL  FILL_1943
timestamp 1713400504
transform 1 0 1736 0 1 1770
box -8 -3 16 105
use FILL  FILL_1944
timestamp 1713400504
transform 1 0 1728 0 1 1770
box -8 -3 16 105
use FILL  FILL_1945
timestamp 1713400504
transform 1 0 1680 0 1 1770
box -8 -3 16 105
use FILL  FILL_1946
timestamp 1713400504
transform 1 0 1672 0 1 1770
box -8 -3 16 105
use FILL  FILL_1947
timestamp 1713400504
transform 1 0 1664 0 1 1770
box -8 -3 16 105
use FILL  FILL_1948
timestamp 1713400504
transform 1 0 1656 0 1 1770
box -8 -3 16 105
use FILL  FILL_1949
timestamp 1713400504
transform 1 0 1648 0 1 1770
box -8 -3 16 105
use FILL  FILL_1950
timestamp 1713400504
transform 1 0 1640 0 1 1770
box -8 -3 16 105
use FILL  FILL_1951
timestamp 1713400504
transform 1 0 1632 0 1 1770
box -8 -3 16 105
use FILL  FILL_1952
timestamp 1713400504
transform 1 0 1624 0 1 1770
box -8 -3 16 105
use FILL  FILL_1953
timestamp 1713400504
transform 1 0 1576 0 1 1770
box -8 -3 16 105
use FILL  FILL_1954
timestamp 1713400504
transform 1 0 1568 0 1 1770
box -8 -3 16 105
use FILL  FILL_1955
timestamp 1713400504
transform 1 0 1560 0 1 1770
box -8 -3 16 105
use FILL  FILL_1956
timestamp 1713400504
transform 1 0 1552 0 1 1770
box -8 -3 16 105
use FILL  FILL_1957
timestamp 1713400504
transform 1 0 1544 0 1 1770
box -8 -3 16 105
use FILL  FILL_1958
timestamp 1713400504
transform 1 0 1520 0 1 1770
box -8 -3 16 105
use FILL  FILL_1959
timestamp 1713400504
transform 1 0 1512 0 1 1770
box -8 -3 16 105
use FILL  FILL_1960
timestamp 1713400504
transform 1 0 1504 0 1 1770
box -8 -3 16 105
use FILL  FILL_1961
timestamp 1713400504
transform 1 0 1496 0 1 1770
box -8 -3 16 105
use FILL  FILL_1962
timestamp 1713400504
transform 1 0 1456 0 1 1770
box -8 -3 16 105
use FILL  FILL_1963
timestamp 1713400504
transform 1 0 1448 0 1 1770
box -8 -3 16 105
use FILL  FILL_1964
timestamp 1713400504
transform 1 0 1440 0 1 1770
box -8 -3 16 105
use FILL  FILL_1965
timestamp 1713400504
transform 1 0 1432 0 1 1770
box -8 -3 16 105
use FILL  FILL_1966
timestamp 1713400504
transform 1 0 1424 0 1 1770
box -8 -3 16 105
use FILL  FILL_1967
timestamp 1713400504
transform 1 0 1416 0 1 1770
box -8 -3 16 105
use FILL  FILL_1968
timestamp 1713400504
transform 1 0 1392 0 1 1770
box -8 -3 16 105
use FILL  FILL_1969
timestamp 1713400504
transform 1 0 1368 0 1 1770
box -8 -3 16 105
use FILL  FILL_1970
timestamp 1713400504
transform 1 0 1360 0 1 1770
box -8 -3 16 105
use FILL  FILL_1971
timestamp 1713400504
transform 1 0 1352 0 1 1770
box -8 -3 16 105
use FILL  FILL_1972
timestamp 1713400504
transform 1 0 1344 0 1 1770
box -8 -3 16 105
use FILL  FILL_1973
timestamp 1713400504
transform 1 0 1304 0 1 1770
box -8 -3 16 105
use FILL  FILL_1974
timestamp 1713400504
transform 1 0 1296 0 1 1770
box -8 -3 16 105
use FILL  FILL_1975
timestamp 1713400504
transform 1 0 1288 0 1 1770
box -8 -3 16 105
use FILL  FILL_1976
timestamp 1713400504
transform 1 0 1264 0 1 1770
box -8 -3 16 105
use FILL  FILL_1977
timestamp 1713400504
transform 1 0 1200 0 1 1770
box -8 -3 16 105
use FILL  FILL_1978
timestamp 1713400504
transform 1 0 1192 0 1 1770
box -8 -3 16 105
use FILL  FILL_1979
timestamp 1713400504
transform 1 0 1184 0 1 1770
box -8 -3 16 105
use FILL  FILL_1980
timestamp 1713400504
transform 1 0 1176 0 1 1770
box -8 -3 16 105
use FILL  FILL_1981
timestamp 1713400504
transform 1 0 1144 0 1 1770
box -8 -3 16 105
use FILL  FILL_1982
timestamp 1713400504
transform 1 0 1136 0 1 1770
box -8 -3 16 105
use FILL  FILL_1983
timestamp 1713400504
transform 1 0 1128 0 1 1770
box -8 -3 16 105
use FILL  FILL_1984
timestamp 1713400504
transform 1 0 1120 0 1 1770
box -8 -3 16 105
use FILL  FILL_1985
timestamp 1713400504
transform 1 0 1112 0 1 1770
box -8 -3 16 105
use FILL  FILL_1986
timestamp 1713400504
transform 1 0 1080 0 1 1770
box -8 -3 16 105
use FILL  FILL_1987
timestamp 1713400504
transform 1 0 1072 0 1 1770
box -8 -3 16 105
use FILL  FILL_1988
timestamp 1713400504
transform 1 0 1064 0 1 1770
box -8 -3 16 105
use FILL  FILL_1989
timestamp 1713400504
transform 1 0 1056 0 1 1770
box -8 -3 16 105
use FILL  FILL_1990
timestamp 1713400504
transform 1 0 1032 0 1 1770
box -8 -3 16 105
use FILL  FILL_1991
timestamp 1713400504
transform 1 0 1024 0 1 1770
box -8 -3 16 105
use FILL  FILL_1992
timestamp 1713400504
transform 1 0 1016 0 1 1770
box -8 -3 16 105
use FILL  FILL_1993
timestamp 1713400504
transform 1 0 1008 0 1 1770
box -8 -3 16 105
use FILL  FILL_1994
timestamp 1713400504
transform 1 0 976 0 1 1770
box -8 -3 16 105
use FILL  FILL_1995
timestamp 1713400504
transform 1 0 968 0 1 1770
box -8 -3 16 105
use FILL  FILL_1996
timestamp 1713400504
transform 1 0 960 0 1 1770
box -8 -3 16 105
use FILL  FILL_1997
timestamp 1713400504
transform 1 0 952 0 1 1770
box -8 -3 16 105
use FILL  FILL_1998
timestamp 1713400504
transform 1 0 944 0 1 1770
box -8 -3 16 105
use FILL  FILL_1999
timestamp 1713400504
transform 1 0 912 0 1 1770
box -8 -3 16 105
use FILL  FILL_2000
timestamp 1713400504
transform 1 0 904 0 1 1770
box -8 -3 16 105
use FILL  FILL_2001
timestamp 1713400504
transform 1 0 896 0 1 1770
box -8 -3 16 105
use FILL  FILL_2002
timestamp 1713400504
transform 1 0 888 0 1 1770
box -8 -3 16 105
use FILL  FILL_2003
timestamp 1713400504
transform 1 0 880 0 1 1770
box -8 -3 16 105
use FILL  FILL_2004
timestamp 1713400504
transform 1 0 872 0 1 1770
box -8 -3 16 105
use FILL  FILL_2005
timestamp 1713400504
transform 1 0 864 0 1 1770
box -8 -3 16 105
use FILL  FILL_2006
timestamp 1713400504
transform 1 0 816 0 1 1770
box -8 -3 16 105
use FILL  FILL_2007
timestamp 1713400504
transform 1 0 808 0 1 1770
box -8 -3 16 105
use FILL  FILL_2008
timestamp 1713400504
transform 1 0 800 0 1 1770
box -8 -3 16 105
use FILL  FILL_2009
timestamp 1713400504
transform 1 0 792 0 1 1770
box -8 -3 16 105
use FILL  FILL_2010
timestamp 1713400504
transform 1 0 784 0 1 1770
box -8 -3 16 105
use FILL  FILL_2011
timestamp 1713400504
transform 1 0 776 0 1 1770
box -8 -3 16 105
use FILL  FILL_2012
timestamp 1713400504
transform 1 0 768 0 1 1770
box -8 -3 16 105
use FILL  FILL_2013
timestamp 1713400504
transform 1 0 760 0 1 1770
box -8 -3 16 105
use FILL  FILL_2014
timestamp 1713400504
transform 1 0 720 0 1 1770
box -8 -3 16 105
use FILL  FILL_2015
timestamp 1713400504
transform 1 0 712 0 1 1770
box -8 -3 16 105
use FILL  FILL_2016
timestamp 1713400504
transform 1 0 704 0 1 1770
box -8 -3 16 105
use FILL  FILL_2017
timestamp 1713400504
transform 1 0 696 0 1 1770
box -8 -3 16 105
use FILL  FILL_2018
timestamp 1713400504
transform 1 0 688 0 1 1770
box -8 -3 16 105
use FILL  FILL_2019
timestamp 1713400504
transform 1 0 680 0 1 1770
box -8 -3 16 105
use FILL  FILL_2020
timestamp 1713400504
transform 1 0 672 0 1 1770
box -8 -3 16 105
use FILL  FILL_2021
timestamp 1713400504
transform 1 0 624 0 1 1770
box -8 -3 16 105
use FILL  FILL_2022
timestamp 1713400504
transform 1 0 616 0 1 1770
box -8 -3 16 105
use FILL  FILL_2023
timestamp 1713400504
transform 1 0 608 0 1 1770
box -8 -3 16 105
use FILL  FILL_2024
timestamp 1713400504
transform 1 0 600 0 1 1770
box -8 -3 16 105
use FILL  FILL_2025
timestamp 1713400504
transform 1 0 592 0 1 1770
box -8 -3 16 105
use FILL  FILL_2026
timestamp 1713400504
transform 1 0 584 0 1 1770
box -8 -3 16 105
use FILL  FILL_2027
timestamp 1713400504
transform 1 0 576 0 1 1770
box -8 -3 16 105
use FILL  FILL_2028
timestamp 1713400504
transform 1 0 568 0 1 1770
box -8 -3 16 105
use FILL  FILL_2029
timestamp 1713400504
transform 1 0 520 0 1 1770
box -8 -3 16 105
use FILL  FILL_2030
timestamp 1713400504
transform 1 0 512 0 1 1770
box -8 -3 16 105
use FILL  FILL_2031
timestamp 1713400504
transform 1 0 504 0 1 1770
box -8 -3 16 105
use FILL  FILL_2032
timestamp 1713400504
transform 1 0 496 0 1 1770
box -8 -3 16 105
use FILL  FILL_2033
timestamp 1713400504
transform 1 0 488 0 1 1770
box -8 -3 16 105
use FILL  FILL_2034
timestamp 1713400504
transform 1 0 480 0 1 1770
box -8 -3 16 105
use FILL  FILL_2035
timestamp 1713400504
transform 1 0 472 0 1 1770
box -8 -3 16 105
use FILL  FILL_2036
timestamp 1713400504
transform 1 0 448 0 1 1770
box -8 -3 16 105
use FILL  FILL_2037
timestamp 1713400504
transform 1 0 440 0 1 1770
box -8 -3 16 105
use FILL  FILL_2038
timestamp 1713400504
transform 1 0 416 0 1 1770
box -8 -3 16 105
use FILL  FILL_2039
timestamp 1713400504
transform 1 0 408 0 1 1770
box -8 -3 16 105
use FILL  FILL_2040
timestamp 1713400504
transform 1 0 400 0 1 1770
box -8 -3 16 105
use FILL  FILL_2041
timestamp 1713400504
transform 1 0 392 0 1 1770
box -8 -3 16 105
use FILL  FILL_2042
timestamp 1713400504
transform 1 0 336 0 1 1770
box -8 -3 16 105
use FILL  FILL_2043
timestamp 1713400504
transform 1 0 328 0 1 1770
box -8 -3 16 105
use FILL  FILL_2044
timestamp 1713400504
transform 1 0 320 0 1 1770
box -8 -3 16 105
use FILL  FILL_2045
timestamp 1713400504
transform 1 0 312 0 1 1770
box -8 -3 16 105
use FILL  FILL_2046
timestamp 1713400504
transform 1 0 304 0 1 1770
box -8 -3 16 105
use FILL  FILL_2047
timestamp 1713400504
transform 1 0 248 0 1 1770
box -8 -3 16 105
use FILL  FILL_2048
timestamp 1713400504
transform 1 0 184 0 1 1770
box -8 -3 16 105
use FILL  FILL_2049
timestamp 1713400504
transform 1 0 176 0 1 1770
box -8 -3 16 105
use FILL  FILL_2050
timestamp 1713400504
transform 1 0 168 0 1 1770
box -8 -3 16 105
use FILL  FILL_2051
timestamp 1713400504
transform 1 0 112 0 1 1770
box -8 -3 16 105
use FILL  FILL_2052
timestamp 1713400504
transform 1 0 104 0 1 1770
box -8 -3 16 105
use FILL  FILL_2053
timestamp 1713400504
transform 1 0 96 0 1 1770
box -8 -3 16 105
use FILL  FILL_2054
timestamp 1713400504
transform 1 0 72 0 1 1770
box -8 -3 16 105
use FILL  FILL_2055
timestamp 1713400504
transform 1 0 3008 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2056
timestamp 1713400504
transform 1 0 2904 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2057
timestamp 1713400504
transform 1 0 2896 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2058
timestamp 1713400504
transform 1 0 2888 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2059
timestamp 1713400504
transform 1 0 2864 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2060
timestamp 1713400504
transform 1 0 2856 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2061
timestamp 1713400504
transform 1 0 2848 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2062
timestamp 1713400504
transform 1 0 2840 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2063
timestamp 1713400504
transform 1 0 2832 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2064
timestamp 1713400504
transform 1 0 2784 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2065
timestamp 1713400504
transform 1 0 2776 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2066
timestamp 1713400504
transform 1 0 2768 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2067
timestamp 1713400504
transform 1 0 2760 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2068
timestamp 1713400504
transform 1 0 2752 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2069
timestamp 1713400504
transform 1 0 2744 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2070
timestamp 1713400504
transform 1 0 2736 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2071
timestamp 1713400504
transform 1 0 2696 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2072
timestamp 1713400504
transform 1 0 2688 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2073
timestamp 1713400504
transform 1 0 2664 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2074
timestamp 1713400504
transform 1 0 2656 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2075
timestamp 1713400504
transform 1 0 2648 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2076
timestamp 1713400504
transform 1 0 2640 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2077
timestamp 1713400504
transform 1 0 2536 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2078
timestamp 1713400504
transform 1 0 2528 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2079
timestamp 1713400504
transform 1 0 2520 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2080
timestamp 1713400504
transform 1 0 2472 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2081
timestamp 1713400504
transform 1 0 2464 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2082
timestamp 1713400504
transform 1 0 2456 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2083
timestamp 1713400504
transform 1 0 2448 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2084
timestamp 1713400504
transform 1 0 2440 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2085
timestamp 1713400504
transform 1 0 2432 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2086
timestamp 1713400504
transform 1 0 2424 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2087
timestamp 1713400504
transform 1 0 2416 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2088
timestamp 1713400504
transform 1 0 2384 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2089
timestamp 1713400504
transform 1 0 2376 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2090
timestamp 1713400504
transform 1 0 2368 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2091
timestamp 1713400504
transform 1 0 2360 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2092
timestamp 1713400504
transform 1 0 2352 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2093
timestamp 1713400504
transform 1 0 2344 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2094
timestamp 1713400504
transform 1 0 2312 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2095
timestamp 1713400504
transform 1 0 2304 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2096
timestamp 1713400504
transform 1 0 2296 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2097
timestamp 1713400504
transform 1 0 2288 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2098
timestamp 1713400504
transform 1 0 2280 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2099
timestamp 1713400504
transform 1 0 2272 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2100
timestamp 1713400504
transform 1 0 2264 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2101
timestamp 1713400504
transform 1 0 2256 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2102
timestamp 1713400504
transform 1 0 2224 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2103
timestamp 1713400504
transform 1 0 2216 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2104
timestamp 1713400504
transform 1 0 2208 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2105
timestamp 1713400504
transform 1 0 2200 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2106
timestamp 1713400504
transform 1 0 2192 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2107
timestamp 1713400504
transform 1 0 2184 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2108
timestamp 1713400504
transform 1 0 2176 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2109
timestamp 1713400504
transform 1 0 2144 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2110
timestamp 1713400504
transform 1 0 2136 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2111
timestamp 1713400504
transform 1 0 2128 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2112
timestamp 1713400504
transform 1 0 2120 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2113
timestamp 1713400504
transform 1 0 2088 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2114
timestamp 1713400504
transform 1 0 2080 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2115
timestamp 1713400504
transform 1 0 2072 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2116
timestamp 1713400504
transform 1 0 2064 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2117
timestamp 1713400504
transform 1 0 2056 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2118
timestamp 1713400504
transform 1 0 2048 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2119
timestamp 1713400504
transform 1 0 2016 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2120
timestamp 1713400504
transform 1 0 2008 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2121
timestamp 1713400504
transform 1 0 2000 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2122
timestamp 1713400504
transform 1 0 1992 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2123
timestamp 1713400504
transform 1 0 1984 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2124
timestamp 1713400504
transform 1 0 1976 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2125
timestamp 1713400504
transform 1 0 1944 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2126
timestamp 1713400504
transform 1 0 1936 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2127
timestamp 1713400504
transform 1 0 1928 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2128
timestamp 1713400504
transform 1 0 1920 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2129
timestamp 1713400504
transform 1 0 1912 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2130
timestamp 1713400504
transform 1 0 1888 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2131
timestamp 1713400504
transform 1 0 1880 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2132
timestamp 1713400504
transform 1 0 1872 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2133
timestamp 1713400504
transform 1 0 1864 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2134
timestamp 1713400504
transform 1 0 1832 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2135
timestamp 1713400504
transform 1 0 1824 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2136
timestamp 1713400504
transform 1 0 1816 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2137
timestamp 1713400504
transform 1 0 1808 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2138
timestamp 1713400504
transform 1 0 1800 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2139
timestamp 1713400504
transform 1 0 1792 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2140
timestamp 1713400504
transform 1 0 1784 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2141
timestamp 1713400504
transform 1 0 1744 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2142
timestamp 1713400504
transform 1 0 1736 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2143
timestamp 1713400504
transform 1 0 1728 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2144
timestamp 1713400504
transform 1 0 1720 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2145
timestamp 1713400504
transform 1 0 1712 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2146
timestamp 1713400504
transform 1 0 1704 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2147
timestamp 1713400504
transform 1 0 1696 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2148
timestamp 1713400504
transform 1 0 1664 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2149
timestamp 1713400504
transform 1 0 1656 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2150
timestamp 1713400504
transform 1 0 1648 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2151
timestamp 1713400504
transform 1 0 1640 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2152
timestamp 1713400504
transform 1 0 1632 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2153
timestamp 1713400504
transform 1 0 1608 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2154
timestamp 1713400504
transform 1 0 1600 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2155
timestamp 1713400504
transform 1 0 1592 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2156
timestamp 1713400504
transform 1 0 1584 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2157
timestamp 1713400504
transform 1 0 1576 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2158
timestamp 1713400504
transform 1 0 1544 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2159
timestamp 1713400504
transform 1 0 1536 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2160
timestamp 1713400504
transform 1 0 1528 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2161
timestamp 1713400504
transform 1 0 1520 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2162
timestamp 1713400504
transform 1 0 1512 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2163
timestamp 1713400504
transform 1 0 1504 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2164
timestamp 1713400504
transform 1 0 1496 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2165
timestamp 1713400504
transform 1 0 1488 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2166
timestamp 1713400504
transform 1 0 1440 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2167
timestamp 1713400504
transform 1 0 1432 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2168
timestamp 1713400504
transform 1 0 1424 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2169
timestamp 1713400504
transform 1 0 1416 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2170
timestamp 1713400504
transform 1 0 1408 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2171
timestamp 1713400504
transform 1 0 1400 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2172
timestamp 1713400504
transform 1 0 1392 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2173
timestamp 1713400504
transform 1 0 1384 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2174
timestamp 1713400504
transform 1 0 1344 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2175
timestamp 1713400504
transform 1 0 1336 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2176
timestamp 1713400504
transform 1 0 1328 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2177
timestamp 1713400504
transform 1 0 1320 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2178
timestamp 1713400504
transform 1 0 1256 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2179
timestamp 1713400504
transform 1 0 1248 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2180
timestamp 1713400504
transform 1 0 1240 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2181
timestamp 1713400504
transform 1 0 1232 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2182
timestamp 1713400504
transform 1 0 1224 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2183
timestamp 1713400504
transform 1 0 1216 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2184
timestamp 1713400504
transform 1 0 1208 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2185
timestamp 1713400504
transform 1 0 1168 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2186
timestamp 1713400504
transform 1 0 1160 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2187
timestamp 1713400504
transform 1 0 1152 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2188
timestamp 1713400504
transform 1 0 1144 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2189
timestamp 1713400504
transform 1 0 1136 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2190
timestamp 1713400504
transform 1 0 1128 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2191
timestamp 1713400504
transform 1 0 1120 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2192
timestamp 1713400504
transform 1 0 1112 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2193
timestamp 1713400504
transform 1 0 1104 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2194
timestamp 1713400504
transform 1 0 1056 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2195
timestamp 1713400504
transform 1 0 1048 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2196
timestamp 1713400504
transform 1 0 1040 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2197
timestamp 1713400504
transform 1 0 1032 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2198
timestamp 1713400504
transform 1 0 1024 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2199
timestamp 1713400504
transform 1 0 1016 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2200
timestamp 1713400504
transform 1 0 1008 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2201
timestamp 1713400504
transform 1 0 1000 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2202
timestamp 1713400504
transform 1 0 992 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2203
timestamp 1713400504
transform 1 0 984 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2204
timestamp 1713400504
transform 1 0 936 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2205
timestamp 1713400504
transform 1 0 928 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2206
timestamp 1713400504
transform 1 0 920 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2207
timestamp 1713400504
transform 1 0 912 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2208
timestamp 1713400504
transform 1 0 904 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2209
timestamp 1713400504
transform 1 0 896 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2210
timestamp 1713400504
transform 1 0 888 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2211
timestamp 1713400504
transform 1 0 880 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2212
timestamp 1713400504
transform 1 0 872 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2213
timestamp 1713400504
transform 1 0 864 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2214
timestamp 1713400504
transform 1 0 816 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2215
timestamp 1713400504
transform 1 0 808 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2216
timestamp 1713400504
transform 1 0 800 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2217
timestamp 1713400504
transform 1 0 792 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2218
timestamp 1713400504
transform 1 0 784 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2219
timestamp 1713400504
transform 1 0 776 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2220
timestamp 1713400504
transform 1 0 768 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2221
timestamp 1713400504
transform 1 0 760 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2222
timestamp 1713400504
transform 1 0 728 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2223
timestamp 1713400504
transform 1 0 720 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2224
timestamp 1713400504
transform 1 0 712 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2225
timestamp 1713400504
transform 1 0 704 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2226
timestamp 1713400504
transform 1 0 696 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2227
timestamp 1713400504
transform 1 0 688 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2228
timestamp 1713400504
transform 1 0 680 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2229
timestamp 1713400504
transform 1 0 672 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2230
timestamp 1713400504
transform 1 0 632 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2231
timestamp 1713400504
transform 1 0 624 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2232
timestamp 1713400504
transform 1 0 616 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2233
timestamp 1713400504
transform 1 0 608 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2234
timestamp 1713400504
transform 1 0 600 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2235
timestamp 1713400504
transform 1 0 592 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2236
timestamp 1713400504
transform 1 0 584 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2237
timestamp 1713400504
transform 1 0 576 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2238
timestamp 1713400504
transform 1 0 568 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2239
timestamp 1713400504
transform 1 0 560 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2240
timestamp 1713400504
transform 1 0 552 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2241
timestamp 1713400504
transform 1 0 544 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2242
timestamp 1713400504
transform 1 0 536 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2243
timestamp 1713400504
transform 1 0 528 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2244
timestamp 1713400504
transform 1 0 520 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2245
timestamp 1713400504
transform 1 0 512 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2246
timestamp 1713400504
transform 1 0 504 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2247
timestamp 1713400504
transform 1 0 496 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2248
timestamp 1713400504
transform 1 0 488 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2249
timestamp 1713400504
transform 1 0 480 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2250
timestamp 1713400504
transform 1 0 472 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2251
timestamp 1713400504
transform 1 0 464 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2252
timestamp 1713400504
transform 1 0 456 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2253
timestamp 1713400504
transform 1 0 448 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2254
timestamp 1713400504
transform 1 0 440 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2255
timestamp 1713400504
transform 1 0 432 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2256
timestamp 1713400504
transform 1 0 424 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2257
timestamp 1713400504
transform 1 0 416 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2258
timestamp 1713400504
transform 1 0 408 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2259
timestamp 1713400504
transform 1 0 400 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2260
timestamp 1713400504
transform 1 0 392 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2261
timestamp 1713400504
transform 1 0 384 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2262
timestamp 1713400504
transform 1 0 376 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2263
timestamp 1713400504
transform 1 0 368 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2264
timestamp 1713400504
transform 1 0 336 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2265
timestamp 1713400504
transform 1 0 328 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2266
timestamp 1713400504
transform 1 0 320 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2267
timestamp 1713400504
transform 1 0 312 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2268
timestamp 1713400504
transform 1 0 304 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2269
timestamp 1713400504
transform 1 0 296 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2270
timestamp 1713400504
transform 1 0 288 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2271
timestamp 1713400504
transform 1 0 280 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2272
timestamp 1713400504
transform 1 0 272 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2273
timestamp 1713400504
transform 1 0 264 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2274
timestamp 1713400504
transform 1 0 256 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2275
timestamp 1713400504
transform 1 0 248 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2276
timestamp 1713400504
transform 1 0 240 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2277
timestamp 1713400504
transform 1 0 232 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2278
timestamp 1713400504
transform 1 0 200 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2279
timestamp 1713400504
transform 1 0 192 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2280
timestamp 1713400504
transform 1 0 184 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2281
timestamp 1713400504
transform 1 0 176 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2282
timestamp 1713400504
transform 1 0 168 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2283
timestamp 1713400504
transform 1 0 160 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2284
timestamp 1713400504
transform 1 0 152 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2285
timestamp 1713400504
transform 1 0 144 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2286
timestamp 1713400504
transform 1 0 136 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2287
timestamp 1713400504
transform 1 0 128 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2288
timestamp 1713400504
transform 1 0 120 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2289
timestamp 1713400504
transform 1 0 112 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2290
timestamp 1713400504
transform 1 0 104 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2291
timestamp 1713400504
transform 1 0 96 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2292
timestamp 1713400504
transform 1 0 88 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2293
timestamp 1713400504
transform 1 0 80 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2294
timestamp 1713400504
transform 1 0 72 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2295
timestamp 1713400504
transform 1 0 3008 0 1 1570
box -8 -3 16 105
use FILL  FILL_2296
timestamp 1713400504
transform 1 0 3000 0 1 1570
box -8 -3 16 105
use FILL  FILL_2297
timestamp 1713400504
transform 1 0 2992 0 1 1570
box -8 -3 16 105
use FILL  FILL_2298
timestamp 1713400504
transform 1 0 2984 0 1 1570
box -8 -3 16 105
use FILL  FILL_2299
timestamp 1713400504
transform 1 0 2976 0 1 1570
box -8 -3 16 105
use FILL  FILL_2300
timestamp 1713400504
transform 1 0 2968 0 1 1570
box -8 -3 16 105
use FILL  FILL_2301
timestamp 1713400504
transform 1 0 2960 0 1 1570
box -8 -3 16 105
use FILL  FILL_2302
timestamp 1713400504
transform 1 0 2856 0 1 1570
box -8 -3 16 105
use FILL  FILL_2303
timestamp 1713400504
transform 1 0 2848 0 1 1570
box -8 -3 16 105
use FILL  FILL_2304
timestamp 1713400504
transform 1 0 2840 0 1 1570
box -8 -3 16 105
use FILL  FILL_2305
timestamp 1713400504
transform 1 0 2832 0 1 1570
box -8 -3 16 105
use FILL  FILL_2306
timestamp 1713400504
transform 1 0 2824 0 1 1570
box -8 -3 16 105
use FILL  FILL_2307
timestamp 1713400504
transform 1 0 2776 0 1 1570
box -8 -3 16 105
use FILL  FILL_2308
timestamp 1713400504
transform 1 0 2768 0 1 1570
box -8 -3 16 105
use FILL  FILL_2309
timestamp 1713400504
transform 1 0 2760 0 1 1570
box -8 -3 16 105
use FILL  FILL_2310
timestamp 1713400504
transform 1 0 2752 0 1 1570
box -8 -3 16 105
use FILL  FILL_2311
timestamp 1713400504
transform 1 0 2744 0 1 1570
box -8 -3 16 105
use FILL  FILL_2312
timestamp 1713400504
transform 1 0 2736 0 1 1570
box -8 -3 16 105
use FILL  FILL_2313
timestamp 1713400504
transform 1 0 2728 0 1 1570
box -8 -3 16 105
use FILL  FILL_2314
timestamp 1713400504
transform 1 0 2704 0 1 1570
box -8 -3 16 105
use FILL  FILL_2315
timestamp 1713400504
transform 1 0 2696 0 1 1570
box -8 -3 16 105
use FILL  FILL_2316
timestamp 1713400504
transform 1 0 2688 0 1 1570
box -8 -3 16 105
use FILL  FILL_2317
timestamp 1713400504
transform 1 0 2648 0 1 1570
box -8 -3 16 105
use FILL  FILL_2318
timestamp 1713400504
transform 1 0 2640 0 1 1570
box -8 -3 16 105
use FILL  FILL_2319
timestamp 1713400504
transform 1 0 2632 0 1 1570
box -8 -3 16 105
use FILL  FILL_2320
timestamp 1713400504
transform 1 0 2624 0 1 1570
box -8 -3 16 105
use FILL  FILL_2321
timestamp 1713400504
transform 1 0 2616 0 1 1570
box -8 -3 16 105
use FILL  FILL_2322
timestamp 1713400504
transform 1 0 2608 0 1 1570
box -8 -3 16 105
use FILL  FILL_2323
timestamp 1713400504
transform 1 0 2576 0 1 1570
box -8 -3 16 105
use FILL  FILL_2324
timestamp 1713400504
transform 1 0 2568 0 1 1570
box -8 -3 16 105
use FILL  FILL_2325
timestamp 1713400504
transform 1 0 2560 0 1 1570
box -8 -3 16 105
use FILL  FILL_2326
timestamp 1713400504
transform 1 0 2552 0 1 1570
box -8 -3 16 105
use FILL  FILL_2327
timestamp 1713400504
transform 1 0 2544 0 1 1570
box -8 -3 16 105
use FILL  FILL_2328
timestamp 1713400504
transform 1 0 2504 0 1 1570
box -8 -3 16 105
use FILL  FILL_2329
timestamp 1713400504
transform 1 0 2496 0 1 1570
box -8 -3 16 105
use FILL  FILL_2330
timestamp 1713400504
transform 1 0 2488 0 1 1570
box -8 -3 16 105
use FILL  FILL_2331
timestamp 1713400504
transform 1 0 2464 0 1 1570
box -8 -3 16 105
use FILL  FILL_2332
timestamp 1713400504
transform 1 0 2456 0 1 1570
box -8 -3 16 105
use FILL  FILL_2333
timestamp 1713400504
transform 1 0 2448 0 1 1570
box -8 -3 16 105
use FILL  FILL_2334
timestamp 1713400504
transform 1 0 2440 0 1 1570
box -8 -3 16 105
use FILL  FILL_2335
timestamp 1713400504
transform 1 0 2432 0 1 1570
box -8 -3 16 105
use FILL  FILL_2336
timestamp 1713400504
transform 1 0 2392 0 1 1570
box -8 -3 16 105
use FILL  FILL_2337
timestamp 1713400504
transform 1 0 2384 0 1 1570
box -8 -3 16 105
use FILL  FILL_2338
timestamp 1713400504
transform 1 0 2376 0 1 1570
box -8 -3 16 105
use FILL  FILL_2339
timestamp 1713400504
transform 1 0 2368 0 1 1570
box -8 -3 16 105
use FILL  FILL_2340
timestamp 1713400504
transform 1 0 2360 0 1 1570
box -8 -3 16 105
use FILL  FILL_2341
timestamp 1713400504
transform 1 0 2320 0 1 1570
box -8 -3 16 105
use FILL  FILL_2342
timestamp 1713400504
transform 1 0 2312 0 1 1570
box -8 -3 16 105
use FILL  FILL_2343
timestamp 1713400504
transform 1 0 2304 0 1 1570
box -8 -3 16 105
use FILL  FILL_2344
timestamp 1713400504
transform 1 0 2296 0 1 1570
box -8 -3 16 105
use FILL  FILL_2345
timestamp 1713400504
transform 1 0 2192 0 1 1570
box -8 -3 16 105
use FILL  FILL_2346
timestamp 1713400504
transform 1 0 2184 0 1 1570
box -8 -3 16 105
use FILL  FILL_2347
timestamp 1713400504
transform 1 0 2176 0 1 1570
box -8 -3 16 105
use FILL  FILL_2348
timestamp 1713400504
transform 1 0 2136 0 1 1570
box -8 -3 16 105
use FILL  FILL_2349
timestamp 1713400504
transform 1 0 2128 0 1 1570
box -8 -3 16 105
use FILL  FILL_2350
timestamp 1713400504
transform 1 0 2120 0 1 1570
box -8 -3 16 105
use FILL  FILL_2351
timestamp 1713400504
transform 1 0 2088 0 1 1570
box -8 -3 16 105
use FILL  FILL_2352
timestamp 1713400504
transform 1 0 2080 0 1 1570
box -8 -3 16 105
use FILL  FILL_2353
timestamp 1713400504
transform 1 0 2072 0 1 1570
box -8 -3 16 105
use FILL  FILL_2354
timestamp 1713400504
transform 1 0 2064 0 1 1570
box -8 -3 16 105
use FILL  FILL_2355
timestamp 1713400504
transform 1 0 2024 0 1 1570
box -8 -3 16 105
use FILL  FILL_2356
timestamp 1713400504
transform 1 0 2016 0 1 1570
box -8 -3 16 105
use FILL  FILL_2357
timestamp 1713400504
transform 1 0 2008 0 1 1570
box -8 -3 16 105
use FILL  FILL_2358
timestamp 1713400504
transform 1 0 2000 0 1 1570
box -8 -3 16 105
use FILL  FILL_2359
timestamp 1713400504
transform 1 0 1992 0 1 1570
box -8 -3 16 105
use FILL  FILL_2360
timestamp 1713400504
transform 1 0 1984 0 1 1570
box -8 -3 16 105
use FILL  FILL_2361
timestamp 1713400504
transform 1 0 1952 0 1 1570
box -8 -3 16 105
use FILL  FILL_2362
timestamp 1713400504
transform 1 0 1944 0 1 1570
box -8 -3 16 105
use FILL  FILL_2363
timestamp 1713400504
transform 1 0 1936 0 1 1570
box -8 -3 16 105
use FILL  FILL_2364
timestamp 1713400504
transform 1 0 1928 0 1 1570
box -8 -3 16 105
use FILL  FILL_2365
timestamp 1713400504
transform 1 0 1896 0 1 1570
box -8 -3 16 105
use FILL  FILL_2366
timestamp 1713400504
transform 1 0 1888 0 1 1570
box -8 -3 16 105
use FILL  FILL_2367
timestamp 1713400504
transform 1 0 1880 0 1 1570
box -8 -3 16 105
use FILL  FILL_2368
timestamp 1713400504
transform 1 0 1872 0 1 1570
box -8 -3 16 105
use FILL  FILL_2369
timestamp 1713400504
transform 1 0 1864 0 1 1570
box -8 -3 16 105
use FILL  FILL_2370
timestamp 1713400504
transform 1 0 1856 0 1 1570
box -8 -3 16 105
use FILL  FILL_2371
timestamp 1713400504
transform 1 0 1848 0 1 1570
box -8 -3 16 105
use FILL  FILL_2372
timestamp 1713400504
transform 1 0 1816 0 1 1570
box -8 -3 16 105
use FILL  FILL_2373
timestamp 1713400504
transform 1 0 1808 0 1 1570
box -8 -3 16 105
use FILL  FILL_2374
timestamp 1713400504
transform 1 0 1800 0 1 1570
box -8 -3 16 105
use FILL  FILL_2375
timestamp 1713400504
transform 1 0 1776 0 1 1570
box -8 -3 16 105
use FILL  FILL_2376
timestamp 1713400504
transform 1 0 1768 0 1 1570
box -8 -3 16 105
use FILL  FILL_2377
timestamp 1713400504
transform 1 0 1760 0 1 1570
box -8 -3 16 105
use FILL  FILL_2378
timestamp 1713400504
transform 1 0 1752 0 1 1570
box -8 -3 16 105
use FILL  FILL_2379
timestamp 1713400504
transform 1 0 1744 0 1 1570
box -8 -3 16 105
use FILL  FILL_2380
timestamp 1713400504
transform 1 0 1736 0 1 1570
box -8 -3 16 105
use FILL  FILL_2381
timestamp 1713400504
transform 1 0 1688 0 1 1570
box -8 -3 16 105
use FILL  FILL_2382
timestamp 1713400504
transform 1 0 1680 0 1 1570
box -8 -3 16 105
use FILL  FILL_2383
timestamp 1713400504
transform 1 0 1672 0 1 1570
box -8 -3 16 105
use FILL  FILL_2384
timestamp 1713400504
transform 1 0 1664 0 1 1570
box -8 -3 16 105
use FILL  FILL_2385
timestamp 1713400504
transform 1 0 1656 0 1 1570
box -8 -3 16 105
use FILL  FILL_2386
timestamp 1713400504
transform 1 0 1648 0 1 1570
box -8 -3 16 105
use FILL  FILL_2387
timestamp 1713400504
transform 1 0 1640 0 1 1570
box -8 -3 16 105
use FILL  FILL_2388
timestamp 1713400504
transform 1 0 1592 0 1 1570
box -8 -3 16 105
use FILL  FILL_2389
timestamp 1713400504
transform 1 0 1584 0 1 1570
box -8 -3 16 105
use FILL  FILL_2390
timestamp 1713400504
transform 1 0 1576 0 1 1570
box -8 -3 16 105
use FILL  FILL_2391
timestamp 1713400504
transform 1 0 1568 0 1 1570
box -8 -3 16 105
use FILL  FILL_2392
timestamp 1713400504
transform 1 0 1560 0 1 1570
box -8 -3 16 105
use FILL  FILL_2393
timestamp 1713400504
transform 1 0 1552 0 1 1570
box -8 -3 16 105
use FILL  FILL_2394
timestamp 1713400504
transform 1 0 1520 0 1 1570
box -8 -3 16 105
use FILL  FILL_2395
timestamp 1713400504
transform 1 0 1512 0 1 1570
box -8 -3 16 105
use FILL  FILL_2396
timestamp 1713400504
transform 1 0 1504 0 1 1570
box -8 -3 16 105
use FILL  FILL_2397
timestamp 1713400504
transform 1 0 1440 0 1 1570
box -8 -3 16 105
use FILL  FILL_2398
timestamp 1713400504
transform 1 0 1432 0 1 1570
box -8 -3 16 105
use FILL  FILL_2399
timestamp 1713400504
transform 1 0 1392 0 1 1570
box -8 -3 16 105
use FILL  FILL_2400
timestamp 1713400504
transform 1 0 1384 0 1 1570
box -8 -3 16 105
use FILL  FILL_2401
timestamp 1713400504
transform 1 0 1376 0 1 1570
box -8 -3 16 105
use FILL  FILL_2402
timestamp 1713400504
transform 1 0 1312 0 1 1570
box -8 -3 16 105
use FILL  FILL_2403
timestamp 1713400504
transform 1 0 1288 0 1 1570
box -8 -3 16 105
use FILL  FILL_2404
timestamp 1713400504
transform 1 0 1280 0 1 1570
box -8 -3 16 105
use FILL  FILL_2405
timestamp 1713400504
transform 1 0 1272 0 1 1570
box -8 -3 16 105
use FILL  FILL_2406
timestamp 1713400504
transform 1 0 1264 0 1 1570
box -8 -3 16 105
use FILL  FILL_2407
timestamp 1713400504
transform 1 0 1256 0 1 1570
box -8 -3 16 105
use FILL  FILL_2408
timestamp 1713400504
transform 1 0 1216 0 1 1570
box -8 -3 16 105
use FILL  FILL_2409
timestamp 1713400504
transform 1 0 1208 0 1 1570
box -8 -3 16 105
use FILL  FILL_2410
timestamp 1713400504
transform 1 0 1200 0 1 1570
box -8 -3 16 105
use FILL  FILL_2411
timestamp 1713400504
transform 1 0 1192 0 1 1570
box -8 -3 16 105
use FILL  FILL_2412
timestamp 1713400504
transform 1 0 1184 0 1 1570
box -8 -3 16 105
use FILL  FILL_2413
timestamp 1713400504
transform 1 0 1176 0 1 1570
box -8 -3 16 105
use FILL  FILL_2414
timestamp 1713400504
transform 1 0 1168 0 1 1570
box -8 -3 16 105
use FILL  FILL_2415
timestamp 1713400504
transform 1 0 1160 0 1 1570
box -8 -3 16 105
use FILL  FILL_2416
timestamp 1713400504
transform 1 0 1112 0 1 1570
box -8 -3 16 105
use FILL  FILL_2417
timestamp 1713400504
transform 1 0 1104 0 1 1570
box -8 -3 16 105
use FILL  FILL_2418
timestamp 1713400504
transform 1 0 1096 0 1 1570
box -8 -3 16 105
use FILL  FILL_2419
timestamp 1713400504
transform 1 0 1088 0 1 1570
box -8 -3 16 105
use FILL  FILL_2420
timestamp 1713400504
transform 1 0 1080 0 1 1570
box -8 -3 16 105
use FILL  FILL_2421
timestamp 1713400504
transform 1 0 1072 0 1 1570
box -8 -3 16 105
use FILL  FILL_2422
timestamp 1713400504
transform 1 0 1064 0 1 1570
box -8 -3 16 105
use FILL  FILL_2423
timestamp 1713400504
transform 1 0 1024 0 1 1570
box -8 -3 16 105
use FILL  FILL_2424
timestamp 1713400504
transform 1 0 1016 0 1 1570
box -8 -3 16 105
use FILL  FILL_2425
timestamp 1713400504
transform 1 0 1008 0 1 1570
box -8 -3 16 105
use FILL  FILL_2426
timestamp 1713400504
transform 1 0 1000 0 1 1570
box -8 -3 16 105
use FILL  FILL_2427
timestamp 1713400504
transform 1 0 992 0 1 1570
box -8 -3 16 105
use FILL  FILL_2428
timestamp 1713400504
transform 1 0 984 0 1 1570
box -8 -3 16 105
use FILL  FILL_2429
timestamp 1713400504
transform 1 0 976 0 1 1570
box -8 -3 16 105
use FILL  FILL_2430
timestamp 1713400504
transform 1 0 928 0 1 1570
box -8 -3 16 105
use FILL  FILL_2431
timestamp 1713400504
transform 1 0 920 0 1 1570
box -8 -3 16 105
use FILL  FILL_2432
timestamp 1713400504
transform 1 0 912 0 1 1570
box -8 -3 16 105
use FILL  FILL_2433
timestamp 1713400504
transform 1 0 904 0 1 1570
box -8 -3 16 105
use FILL  FILL_2434
timestamp 1713400504
transform 1 0 896 0 1 1570
box -8 -3 16 105
use FILL  FILL_2435
timestamp 1713400504
transform 1 0 888 0 1 1570
box -8 -3 16 105
use FILL  FILL_2436
timestamp 1713400504
transform 1 0 880 0 1 1570
box -8 -3 16 105
use FILL  FILL_2437
timestamp 1713400504
transform 1 0 872 0 1 1570
box -8 -3 16 105
use FILL  FILL_2438
timestamp 1713400504
transform 1 0 832 0 1 1570
box -8 -3 16 105
use FILL  FILL_2439
timestamp 1713400504
transform 1 0 824 0 1 1570
box -8 -3 16 105
use FILL  FILL_2440
timestamp 1713400504
transform 1 0 816 0 1 1570
box -8 -3 16 105
use FILL  FILL_2441
timestamp 1713400504
transform 1 0 792 0 1 1570
box -8 -3 16 105
use FILL  FILL_2442
timestamp 1713400504
transform 1 0 784 0 1 1570
box -8 -3 16 105
use FILL  FILL_2443
timestamp 1713400504
transform 1 0 776 0 1 1570
box -8 -3 16 105
use FILL  FILL_2444
timestamp 1713400504
transform 1 0 768 0 1 1570
box -8 -3 16 105
use FILL  FILL_2445
timestamp 1713400504
transform 1 0 760 0 1 1570
box -8 -3 16 105
use FILL  FILL_2446
timestamp 1713400504
transform 1 0 752 0 1 1570
box -8 -3 16 105
use FILL  FILL_2447
timestamp 1713400504
transform 1 0 704 0 1 1570
box -8 -3 16 105
use FILL  FILL_2448
timestamp 1713400504
transform 1 0 696 0 1 1570
box -8 -3 16 105
use FILL  FILL_2449
timestamp 1713400504
transform 1 0 688 0 1 1570
box -8 -3 16 105
use FILL  FILL_2450
timestamp 1713400504
transform 1 0 680 0 1 1570
box -8 -3 16 105
use FILL  FILL_2451
timestamp 1713400504
transform 1 0 576 0 1 1570
box -8 -3 16 105
use FILL  FILL_2452
timestamp 1713400504
transform 1 0 568 0 1 1570
box -8 -3 16 105
use FILL  FILL_2453
timestamp 1713400504
transform 1 0 560 0 1 1570
box -8 -3 16 105
use FILL  FILL_2454
timestamp 1713400504
transform 1 0 520 0 1 1570
box -8 -3 16 105
use FILL  FILL_2455
timestamp 1713400504
transform 1 0 512 0 1 1570
box -8 -3 16 105
use FILL  FILL_2456
timestamp 1713400504
transform 1 0 480 0 1 1570
box -8 -3 16 105
use FILL  FILL_2457
timestamp 1713400504
transform 1 0 472 0 1 1570
box -8 -3 16 105
use FILL  FILL_2458
timestamp 1713400504
transform 1 0 368 0 1 1570
box -8 -3 16 105
use FILL  FILL_2459
timestamp 1713400504
transform 1 0 328 0 1 1570
box -8 -3 16 105
use FILL  FILL_2460
timestamp 1713400504
transform 1 0 320 0 1 1570
box -8 -3 16 105
use FILL  FILL_2461
timestamp 1713400504
transform 1 0 216 0 1 1570
box -8 -3 16 105
use FILL  FILL_2462
timestamp 1713400504
transform 1 0 208 0 1 1570
box -8 -3 16 105
use FILL  FILL_2463
timestamp 1713400504
transform 1 0 168 0 1 1570
box -8 -3 16 105
use FILL  FILL_2464
timestamp 1713400504
transform 1 0 3008 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2465
timestamp 1713400504
transform 1 0 2904 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2466
timestamp 1713400504
transform 1 0 2896 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2467
timestamp 1713400504
transform 1 0 2888 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2468
timestamp 1713400504
transform 1 0 2864 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2469
timestamp 1713400504
transform 1 0 2856 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2470
timestamp 1713400504
transform 1 0 2752 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2471
timestamp 1713400504
transform 1 0 2744 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2472
timestamp 1713400504
transform 1 0 2720 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2473
timestamp 1713400504
transform 1 0 2712 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2474
timestamp 1713400504
transform 1 0 2704 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2475
timestamp 1713400504
transform 1 0 2696 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2476
timestamp 1713400504
transform 1 0 2648 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2477
timestamp 1713400504
transform 1 0 2640 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2478
timestamp 1713400504
transform 1 0 2632 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2479
timestamp 1713400504
transform 1 0 2624 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2480
timestamp 1713400504
transform 1 0 2616 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2481
timestamp 1713400504
transform 1 0 2608 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2482
timestamp 1713400504
transform 1 0 2560 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2483
timestamp 1713400504
transform 1 0 2552 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2484
timestamp 1713400504
transform 1 0 2544 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2485
timestamp 1713400504
transform 1 0 2536 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2486
timestamp 1713400504
transform 1 0 2528 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2487
timestamp 1713400504
transform 1 0 2520 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2488
timestamp 1713400504
transform 1 0 2512 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2489
timestamp 1713400504
transform 1 0 2504 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2490
timestamp 1713400504
transform 1 0 2464 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2491
timestamp 1713400504
transform 1 0 2456 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2492
timestamp 1713400504
transform 1 0 2448 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2493
timestamp 1713400504
transform 1 0 2440 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2494
timestamp 1713400504
transform 1 0 2432 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2495
timestamp 1713400504
transform 1 0 2392 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2496
timestamp 1713400504
transform 1 0 2384 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2497
timestamp 1713400504
transform 1 0 2376 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2498
timestamp 1713400504
transform 1 0 2368 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2499
timestamp 1713400504
transform 1 0 2360 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2500
timestamp 1713400504
transform 1 0 2328 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2501
timestamp 1713400504
transform 1 0 2320 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2502
timestamp 1713400504
transform 1 0 2312 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2503
timestamp 1713400504
transform 1 0 2304 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2504
timestamp 1713400504
transform 1 0 2272 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2505
timestamp 1713400504
transform 1 0 2264 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2506
timestamp 1713400504
transform 1 0 2256 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2507
timestamp 1713400504
transform 1 0 2248 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2508
timestamp 1713400504
transform 1 0 2240 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2509
timestamp 1713400504
transform 1 0 2232 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2510
timestamp 1713400504
transform 1 0 2208 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2511
timestamp 1713400504
transform 1 0 2200 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2512
timestamp 1713400504
transform 1 0 2192 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2513
timestamp 1713400504
transform 1 0 2184 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2514
timestamp 1713400504
transform 1 0 2152 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2515
timestamp 1713400504
transform 1 0 2144 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2516
timestamp 1713400504
transform 1 0 2136 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2517
timestamp 1713400504
transform 1 0 2128 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2518
timestamp 1713400504
transform 1 0 2104 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2519
timestamp 1713400504
transform 1 0 2096 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2520
timestamp 1713400504
transform 1 0 2088 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2521
timestamp 1713400504
transform 1 0 2080 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2522
timestamp 1713400504
transform 1 0 2072 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2523
timestamp 1713400504
transform 1 0 1968 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2524
timestamp 1713400504
transform 1 0 1960 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2525
timestamp 1713400504
transform 1 0 1952 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2526
timestamp 1713400504
transform 1 0 1944 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2527
timestamp 1713400504
transform 1 0 1936 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2528
timestamp 1713400504
transform 1 0 1888 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2529
timestamp 1713400504
transform 1 0 1880 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2530
timestamp 1713400504
transform 1 0 1872 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2531
timestamp 1713400504
transform 1 0 1864 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2532
timestamp 1713400504
transform 1 0 1856 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2533
timestamp 1713400504
transform 1 0 1848 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2534
timestamp 1713400504
transform 1 0 1840 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2535
timestamp 1713400504
transform 1 0 1832 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2536
timestamp 1713400504
transform 1 0 1784 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2537
timestamp 1713400504
transform 1 0 1776 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2538
timestamp 1713400504
transform 1 0 1768 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2539
timestamp 1713400504
transform 1 0 1760 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2540
timestamp 1713400504
transform 1 0 1752 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2541
timestamp 1713400504
transform 1 0 1744 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2542
timestamp 1713400504
transform 1 0 1736 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2543
timestamp 1713400504
transform 1 0 1696 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2544
timestamp 1713400504
transform 1 0 1688 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2545
timestamp 1713400504
transform 1 0 1680 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2546
timestamp 1713400504
transform 1 0 1672 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2547
timestamp 1713400504
transform 1 0 1664 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2548
timestamp 1713400504
transform 1 0 1632 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2549
timestamp 1713400504
transform 1 0 1624 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2550
timestamp 1713400504
transform 1 0 1616 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2551
timestamp 1713400504
transform 1 0 1608 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2552
timestamp 1713400504
transform 1 0 1600 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2553
timestamp 1713400504
transform 1 0 1592 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2554
timestamp 1713400504
transform 1 0 1584 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2555
timestamp 1713400504
transform 1 0 1544 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2556
timestamp 1713400504
transform 1 0 1536 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2557
timestamp 1713400504
transform 1 0 1528 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2558
timestamp 1713400504
transform 1 0 1520 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2559
timestamp 1713400504
transform 1 0 1512 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2560
timestamp 1713400504
transform 1 0 1504 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2561
timestamp 1713400504
transform 1 0 1496 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2562
timestamp 1713400504
transform 1 0 1488 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2563
timestamp 1713400504
transform 1 0 1448 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2564
timestamp 1713400504
transform 1 0 1440 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2565
timestamp 1713400504
transform 1 0 1432 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2566
timestamp 1713400504
transform 1 0 1424 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2567
timestamp 1713400504
transform 1 0 1416 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2568
timestamp 1713400504
transform 1 0 1408 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2569
timestamp 1713400504
transform 1 0 1400 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2570
timestamp 1713400504
transform 1 0 1392 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2571
timestamp 1713400504
transform 1 0 1352 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2572
timestamp 1713400504
transform 1 0 1344 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2573
timestamp 1713400504
transform 1 0 1336 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2574
timestamp 1713400504
transform 1 0 1328 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2575
timestamp 1713400504
transform 1 0 1320 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2576
timestamp 1713400504
transform 1 0 1312 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2577
timestamp 1713400504
transform 1 0 1304 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2578
timestamp 1713400504
transform 1 0 1296 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2579
timestamp 1713400504
transform 1 0 1248 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2580
timestamp 1713400504
transform 1 0 1240 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2581
timestamp 1713400504
transform 1 0 1232 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2582
timestamp 1713400504
transform 1 0 1224 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2583
timestamp 1713400504
transform 1 0 1216 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2584
timestamp 1713400504
transform 1 0 1208 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2585
timestamp 1713400504
transform 1 0 1200 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2586
timestamp 1713400504
transform 1 0 1192 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2587
timestamp 1713400504
transform 1 0 1184 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2588
timestamp 1713400504
transform 1 0 1144 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2589
timestamp 1713400504
transform 1 0 1136 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2590
timestamp 1713400504
transform 1 0 1128 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2591
timestamp 1713400504
transform 1 0 1120 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2592
timestamp 1713400504
transform 1 0 1112 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2593
timestamp 1713400504
transform 1 0 1104 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2594
timestamp 1713400504
transform 1 0 1096 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2595
timestamp 1713400504
transform 1 0 1088 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2596
timestamp 1713400504
transform 1 0 1080 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2597
timestamp 1713400504
transform 1 0 1032 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2598
timestamp 1713400504
transform 1 0 1024 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2599
timestamp 1713400504
transform 1 0 1016 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2600
timestamp 1713400504
transform 1 0 1008 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2601
timestamp 1713400504
transform 1 0 1000 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2602
timestamp 1713400504
transform 1 0 992 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2603
timestamp 1713400504
transform 1 0 984 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2604
timestamp 1713400504
transform 1 0 976 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2605
timestamp 1713400504
transform 1 0 968 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2606
timestamp 1713400504
transform 1 0 928 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2607
timestamp 1713400504
transform 1 0 920 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2608
timestamp 1713400504
transform 1 0 912 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2609
timestamp 1713400504
transform 1 0 904 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2610
timestamp 1713400504
transform 1 0 896 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2611
timestamp 1713400504
transform 1 0 888 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2612
timestamp 1713400504
transform 1 0 880 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2613
timestamp 1713400504
transform 1 0 872 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2614
timestamp 1713400504
transform 1 0 864 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2615
timestamp 1713400504
transform 1 0 856 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2616
timestamp 1713400504
transform 1 0 808 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2617
timestamp 1713400504
transform 1 0 800 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2618
timestamp 1713400504
transform 1 0 792 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2619
timestamp 1713400504
transform 1 0 784 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2620
timestamp 1713400504
transform 1 0 776 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2621
timestamp 1713400504
transform 1 0 768 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2622
timestamp 1713400504
transform 1 0 760 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2623
timestamp 1713400504
transform 1 0 752 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2624
timestamp 1713400504
transform 1 0 744 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2625
timestamp 1713400504
transform 1 0 696 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2626
timestamp 1713400504
transform 1 0 688 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2627
timestamp 1713400504
transform 1 0 680 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2628
timestamp 1713400504
transform 1 0 672 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2629
timestamp 1713400504
transform 1 0 664 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2630
timestamp 1713400504
transform 1 0 656 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2631
timestamp 1713400504
transform 1 0 648 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2632
timestamp 1713400504
transform 1 0 640 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2633
timestamp 1713400504
transform 1 0 632 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2634
timestamp 1713400504
transform 1 0 624 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2635
timestamp 1713400504
transform 1 0 616 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2636
timestamp 1713400504
transform 1 0 608 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2637
timestamp 1713400504
transform 1 0 600 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2638
timestamp 1713400504
transform 1 0 592 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2639
timestamp 1713400504
transform 1 0 488 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2640
timestamp 1713400504
transform 1 0 480 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2641
timestamp 1713400504
transform 1 0 376 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2642
timestamp 1713400504
transform 1 0 368 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2643
timestamp 1713400504
transform 1 0 360 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2644
timestamp 1713400504
transform 1 0 352 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2645
timestamp 1713400504
transform 1 0 320 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2646
timestamp 1713400504
transform 1 0 312 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2647
timestamp 1713400504
transform 1 0 304 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2648
timestamp 1713400504
transform 1 0 296 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2649
timestamp 1713400504
transform 1 0 288 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2650
timestamp 1713400504
transform 1 0 248 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2651
timestamp 1713400504
transform 1 0 240 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2652
timestamp 1713400504
transform 1 0 232 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2653
timestamp 1713400504
transform 1 0 224 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2654
timestamp 1713400504
transform 1 0 120 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2655
timestamp 1713400504
transform 1 0 112 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2656
timestamp 1713400504
transform 1 0 104 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2657
timestamp 1713400504
transform 1 0 96 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2658
timestamp 1713400504
transform 1 0 88 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2659
timestamp 1713400504
transform 1 0 80 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2660
timestamp 1713400504
transform 1 0 72 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2661
timestamp 1713400504
transform 1 0 3008 0 1 1370
box -8 -3 16 105
use FILL  FILL_2662
timestamp 1713400504
transform 1 0 2904 0 1 1370
box -8 -3 16 105
use FILL  FILL_2663
timestamp 1713400504
transform 1 0 2896 0 1 1370
box -8 -3 16 105
use FILL  FILL_2664
timestamp 1713400504
transform 1 0 2856 0 1 1370
box -8 -3 16 105
use FILL  FILL_2665
timestamp 1713400504
transform 1 0 2848 0 1 1370
box -8 -3 16 105
use FILL  FILL_2666
timestamp 1713400504
transform 1 0 2840 0 1 1370
box -8 -3 16 105
use FILL  FILL_2667
timestamp 1713400504
transform 1 0 2832 0 1 1370
box -8 -3 16 105
use FILL  FILL_2668
timestamp 1713400504
transform 1 0 2824 0 1 1370
box -8 -3 16 105
use FILL  FILL_2669
timestamp 1713400504
transform 1 0 2816 0 1 1370
box -8 -3 16 105
use FILL  FILL_2670
timestamp 1713400504
transform 1 0 2808 0 1 1370
box -8 -3 16 105
use FILL  FILL_2671
timestamp 1713400504
transform 1 0 2760 0 1 1370
box -8 -3 16 105
use FILL  FILL_2672
timestamp 1713400504
transform 1 0 2752 0 1 1370
box -8 -3 16 105
use FILL  FILL_2673
timestamp 1713400504
transform 1 0 2744 0 1 1370
box -8 -3 16 105
use FILL  FILL_2674
timestamp 1713400504
transform 1 0 2736 0 1 1370
box -8 -3 16 105
use FILL  FILL_2675
timestamp 1713400504
transform 1 0 2728 0 1 1370
box -8 -3 16 105
use FILL  FILL_2676
timestamp 1713400504
transform 1 0 2720 0 1 1370
box -8 -3 16 105
use FILL  FILL_2677
timestamp 1713400504
transform 1 0 2712 0 1 1370
box -8 -3 16 105
use FILL  FILL_2678
timestamp 1713400504
transform 1 0 2656 0 1 1370
box -8 -3 16 105
use FILL  FILL_2679
timestamp 1713400504
transform 1 0 2552 0 1 1370
box -8 -3 16 105
use FILL  FILL_2680
timestamp 1713400504
transform 1 0 2544 0 1 1370
box -8 -3 16 105
use FILL  FILL_2681
timestamp 1713400504
transform 1 0 2536 0 1 1370
box -8 -3 16 105
use FILL  FILL_2682
timestamp 1713400504
transform 1 0 2496 0 1 1370
box -8 -3 16 105
use FILL  FILL_2683
timestamp 1713400504
transform 1 0 2488 0 1 1370
box -8 -3 16 105
use FILL  FILL_2684
timestamp 1713400504
transform 1 0 2480 0 1 1370
box -8 -3 16 105
use FILL  FILL_2685
timestamp 1713400504
transform 1 0 2472 0 1 1370
box -8 -3 16 105
use FILL  FILL_2686
timestamp 1713400504
transform 1 0 2464 0 1 1370
box -8 -3 16 105
use FILL  FILL_2687
timestamp 1713400504
transform 1 0 2456 0 1 1370
box -8 -3 16 105
use FILL  FILL_2688
timestamp 1713400504
transform 1 0 2424 0 1 1370
box -8 -3 16 105
use FILL  FILL_2689
timestamp 1713400504
transform 1 0 2416 0 1 1370
box -8 -3 16 105
use FILL  FILL_2690
timestamp 1713400504
transform 1 0 2408 0 1 1370
box -8 -3 16 105
use FILL  FILL_2691
timestamp 1713400504
transform 1 0 2400 0 1 1370
box -8 -3 16 105
use FILL  FILL_2692
timestamp 1713400504
transform 1 0 2376 0 1 1370
box -8 -3 16 105
use FILL  FILL_2693
timestamp 1713400504
transform 1 0 2368 0 1 1370
box -8 -3 16 105
use FILL  FILL_2694
timestamp 1713400504
transform 1 0 2360 0 1 1370
box -8 -3 16 105
use FILL  FILL_2695
timestamp 1713400504
transform 1 0 2352 0 1 1370
box -8 -3 16 105
use FILL  FILL_2696
timestamp 1713400504
transform 1 0 2328 0 1 1370
box -8 -3 16 105
use FILL  FILL_2697
timestamp 1713400504
transform 1 0 2320 0 1 1370
box -8 -3 16 105
use FILL  FILL_2698
timestamp 1713400504
transform 1 0 2312 0 1 1370
box -8 -3 16 105
use FILL  FILL_2699
timestamp 1713400504
transform 1 0 2304 0 1 1370
box -8 -3 16 105
use FILL  FILL_2700
timestamp 1713400504
transform 1 0 2296 0 1 1370
box -8 -3 16 105
use FILL  FILL_2701
timestamp 1713400504
transform 1 0 2264 0 1 1370
box -8 -3 16 105
use FILL  FILL_2702
timestamp 1713400504
transform 1 0 2256 0 1 1370
box -8 -3 16 105
use FILL  FILL_2703
timestamp 1713400504
transform 1 0 2248 0 1 1370
box -8 -3 16 105
use FILL  FILL_2704
timestamp 1713400504
transform 1 0 2240 0 1 1370
box -8 -3 16 105
use FILL  FILL_2705
timestamp 1713400504
transform 1 0 2176 0 1 1370
box -8 -3 16 105
use FILL  FILL_2706
timestamp 1713400504
transform 1 0 2168 0 1 1370
box -8 -3 16 105
use FILL  FILL_2707
timestamp 1713400504
transform 1 0 2104 0 1 1370
box -8 -3 16 105
use FILL  FILL_2708
timestamp 1713400504
transform 1 0 2096 0 1 1370
box -8 -3 16 105
use FILL  FILL_2709
timestamp 1713400504
transform 1 0 2088 0 1 1370
box -8 -3 16 105
use FILL  FILL_2710
timestamp 1713400504
transform 1 0 2080 0 1 1370
box -8 -3 16 105
use FILL  FILL_2711
timestamp 1713400504
transform 1 0 2072 0 1 1370
box -8 -3 16 105
use FILL  FILL_2712
timestamp 1713400504
transform 1 0 2024 0 1 1370
box -8 -3 16 105
use FILL  FILL_2713
timestamp 1713400504
transform 1 0 2016 0 1 1370
box -8 -3 16 105
use FILL  FILL_2714
timestamp 1713400504
transform 1 0 2008 0 1 1370
box -8 -3 16 105
use FILL  FILL_2715
timestamp 1713400504
transform 1 0 2000 0 1 1370
box -8 -3 16 105
use FILL  FILL_2716
timestamp 1713400504
transform 1 0 1992 0 1 1370
box -8 -3 16 105
use FILL  FILL_2717
timestamp 1713400504
transform 1 0 1984 0 1 1370
box -8 -3 16 105
use FILL  FILL_2718
timestamp 1713400504
transform 1 0 1976 0 1 1370
box -8 -3 16 105
use FILL  FILL_2719
timestamp 1713400504
transform 1 0 1968 0 1 1370
box -8 -3 16 105
use FILL  FILL_2720
timestamp 1713400504
transform 1 0 1960 0 1 1370
box -8 -3 16 105
use FILL  FILL_2721
timestamp 1713400504
transform 1 0 1912 0 1 1370
box -8 -3 16 105
use FILL  FILL_2722
timestamp 1713400504
transform 1 0 1904 0 1 1370
box -8 -3 16 105
use FILL  FILL_2723
timestamp 1713400504
transform 1 0 1896 0 1 1370
box -8 -3 16 105
use FILL  FILL_2724
timestamp 1713400504
transform 1 0 1888 0 1 1370
box -8 -3 16 105
use FILL  FILL_2725
timestamp 1713400504
transform 1 0 1880 0 1 1370
box -8 -3 16 105
use FILL  FILL_2726
timestamp 1713400504
transform 1 0 1872 0 1 1370
box -8 -3 16 105
use FILL  FILL_2727
timestamp 1713400504
transform 1 0 1864 0 1 1370
box -8 -3 16 105
use FILL  FILL_2728
timestamp 1713400504
transform 1 0 1840 0 1 1370
box -8 -3 16 105
use FILL  FILL_2729
timestamp 1713400504
transform 1 0 1832 0 1 1370
box -8 -3 16 105
use FILL  FILL_2730
timestamp 1713400504
transform 1 0 1824 0 1 1370
box -8 -3 16 105
use FILL  FILL_2731
timestamp 1713400504
transform 1 0 1816 0 1 1370
box -8 -3 16 105
use FILL  FILL_2732
timestamp 1713400504
transform 1 0 1808 0 1 1370
box -8 -3 16 105
use FILL  FILL_2733
timestamp 1713400504
transform 1 0 1768 0 1 1370
box -8 -3 16 105
use FILL  FILL_2734
timestamp 1713400504
transform 1 0 1760 0 1 1370
box -8 -3 16 105
use FILL  FILL_2735
timestamp 1713400504
transform 1 0 1752 0 1 1370
box -8 -3 16 105
use FILL  FILL_2736
timestamp 1713400504
transform 1 0 1744 0 1 1370
box -8 -3 16 105
use FILL  FILL_2737
timestamp 1713400504
transform 1 0 1736 0 1 1370
box -8 -3 16 105
use FILL  FILL_2738
timestamp 1713400504
transform 1 0 1712 0 1 1370
box -8 -3 16 105
use FILL  FILL_2739
timestamp 1713400504
transform 1 0 1704 0 1 1370
box -8 -3 16 105
use FILL  FILL_2740
timestamp 1713400504
transform 1 0 1696 0 1 1370
box -8 -3 16 105
use FILL  FILL_2741
timestamp 1713400504
transform 1 0 1688 0 1 1370
box -8 -3 16 105
use FILL  FILL_2742
timestamp 1713400504
transform 1 0 1680 0 1 1370
box -8 -3 16 105
use FILL  FILL_2743
timestamp 1713400504
transform 1 0 1640 0 1 1370
box -8 -3 16 105
use FILL  FILL_2744
timestamp 1713400504
transform 1 0 1632 0 1 1370
box -8 -3 16 105
use FILL  FILL_2745
timestamp 1713400504
transform 1 0 1624 0 1 1370
box -8 -3 16 105
use FILL  FILL_2746
timestamp 1713400504
transform 1 0 1616 0 1 1370
box -8 -3 16 105
use FILL  FILL_2747
timestamp 1713400504
transform 1 0 1608 0 1 1370
box -8 -3 16 105
use FILL  FILL_2748
timestamp 1713400504
transform 1 0 1600 0 1 1370
box -8 -3 16 105
use FILL  FILL_2749
timestamp 1713400504
transform 1 0 1592 0 1 1370
box -8 -3 16 105
use FILL  FILL_2750
timestamp 1713400504
transform 1 0 1552 0 1 1370
box -8 -3 16 105
use FILL  FILL_2751
timestamp 1713400504
transform 1 0 1544 0 1 1370
box -8 -3 16 105
use FILL  FILL_2752
timestamp 1713400504
transform 1 0 1536 0 1 1370
box -8 -3 16 105
use FILL  FILL_2753
timestamp 1713400504
transform 1 0 1528 0 1 1370
box -8 -3 16 105
use FILL  FILL_2754
timestamp 1713400504
transform 1 0 1520 0 1 1370
box -8 -3 16 105
use FILL  FILL_2755
timestamp 1713400504
transform 1 0 1512 0 1 1370
box -8 -3 16 105
use FILL  FILL_2756
timestamp 1713400504
transform 1 0 1504 0 1 1370
box -8 -3 16 105
use FILL  FILL_2757
timestamp 1713400504
transform 1 0 1496 0 1 1370
box -8 -3 16 105
use FILL  FILL_2758
timestamp 1713400504
transform 1 0 1448 0 1 1370
box -8 -3 16 105
use FILL  FILL_2759
timestamp 1713400504
transform 1 0 1440 0 1 1370
box -8 -3 16 105
use FILL  FILL_2760
timestamp 1713400504
transform 1 0 1432 0 1 1370
box -8 -3 16 105
use FILL  FILL_2761
timestamp 1713400504
transform 1 0 1424 0 1 1370
box -8 -3 16 105
use FILL  FILL_2762
timestamp 1713400504
transform 1 0 1416 0 1 1370
box -8 -3 16 105
use FILL  FILL_2763
timestamp 1713400504
transform 1 0 1408 0 1 1370
box -8 -3 16 105
use FILL  FILL_2764
timestamp 1713400504
transform 1 0 1400 0 1 1370
box -8 -3 16 105
use FILL  FILL_2765
timestamp 1713400504
transform 1 0 1360 0 1 1370
box -8 -3 16 105
use FILL  FILL_2766
timestamp 1713400504
transform 1 0 1352 0 1 1370
box -8 -3 16 105
use FILL  FILL_2767
timestamp 1713400504
transform 1 0 1344 0 1 1370
box -8 -3 16 105
use FILL  FILL_2768
timestamp 1713400504
transform 1 0 1336 0 1 1370
box -8 -3 16 105
use FILL  FILL_2769
timestamp 1713400504
transform 1 0 1296 0 1 1370
box -8 -3 16 105
use FILL  FILL_2770
timestamp 1713400504
transform 1 0 1288 0 1 1370
box -8 -3 16 105
use FILL  FILL_2771
timestamp 1713400504
transform 1 0 1280 0 1 1370
box -8 -3 16 105
use FILL  FILL_2772
timestamp 1713400504
transform 1 0 1272 0 1 1370
box -8 -3 16 105
use FILL  FILL_2773
timestamp 1713400504
transform 1 0 1208 0 1 1370
box -8 -3 16 105
use FILL  FILL_2774
timestamp 1713400504
transform 1 0 1200 0 1 1370
box -8 -3 16 105
use FILL  FILL_2775
timestamp 1713400504
transform 1 0 1192 0 1 1370
box -8 -3 16 105
use FILL  FILL_2776
timestamp 1713400504
transform 1 0 1184 0 1 1370
box -8 -3 16 105
use FILL  FILL_2777
timestamp 1713400504
transform 1 0 1152 0 1 1370
box -8 -3 16 105
use FILL  FILL_2778
timestamp 1713400504
transform 1 0 1144 0 1 1370
box -8 -3 16 105
use FILL  FILL_2779
timestamp 1713400504
transform 1 0 1136 0 1 1370
box -8 -3 16 105
use FILL  FILL_2780
timestamp 1713400504
transform 1 0 1128 0 1 1370
box -8 -3 16 105
use FILL  FILL_2781
timestamp 1713400504
transform 1 0 1120 0 1 1370
box -8 -3 16 105
use FILL  FILL_2782
timestamp 1713400504
transform 1 0 1112 0 1 1370
box -8 -3 16 105
use FILL  FILL_2783
timestamp 1713400504
transform 1 0 1080 0 1 1370
box -8 -3 16 105
use FILL  FILL_2784
timestamp 1713400504
transform 1 0 1072 0 1 1370
box -8 -3 16 105
use FILL  FILL_2785
timestamp 1713400504
transform 1 0 1064 0 1 1370
box -8 -3 16 105
use FILL  FILL_2786
timestamp 1713400504
transform 1 0 1056 0 1 1370
box -8 -3 16 105
use FILL  FILL_2787
timestamp 1713400504
transform 1 0 1048 0 1 1370
box -8 -3 16 105
use FILL  FILL_2788
timestamp 1713400504
transform 1 0 1040 0 1 1370
box -8 -3 16 105
use FILL  FILL_2789
timestamp 1713400504
transform 1 0 1032 0 1 1370
box -8 -3 16 105
use FILL  FILL_2790
timestamp 1713400504
transform 1 0 1024 0 1 1370
box -8 -3 16 105
use FILL  FILL_2791
timestamp 1713400504
transform 1 0 976 0 1 1370
box -8 -3 16 105
use FILL  FILL_2792
timestamp 1713400504
transform 1 0 968 0 1 1370
box -8 -3 16 105
use FILL  FILL_2793
timestamp 1713400504
transform 1 0 960 0 1 1370
box -8 -3 16 105
use FILL  FILL_2794
timestamp 1713400504
transform 1 0 952 0 1 1370
box -8 -3 16 105
use FILL  FILL_2795
timestamp 1713400504
transform 1 0 944 0 1 1370
box -8 -3 16 105
use FILL  FILL_2796
timestamp 1713400504
transform 1 0 936 0 1 1370
box -8 -3 16 105
use FILL  FILL_2797
timestamp 1713400504
transform 1 0 928 0 1 1370
box -8 -3 16 105
use FILL  FILL_2798
timestamp 1713400504
transform 1 0 920 0 1 1370
box -8 -3 16 105
use FILL  FILL_2799
timestamp 1713400504
transform 1 0 880 0 1 1370
box -8 -3 16 105
use FILL  FILL_2800
timestamp 1713400504
transform 1 0 872 0 1 1370
box -8 -3 16 105
use FILL  FILL_2801
timestamp 1713400504
transform 1 0 864 0 1 1370
box -8 -3 16 105
use FILL  FILL_2802
timestamp 1713400504
transform 1 0 856 0 1 1370
box -8 -3 16 105
use FILL  FILL_2803
timestamp 1713400504
transform 1 0 848 0 1 1370
box -8 -3 16 105
use FILL  FILL_2804
timestamp 1713400504
transform 1 0 840 0 1 1370
box -8 -3 16 105
use FILL  FILL_2805
timestamp 1713400504
transform 1 0 832 0 1 1370
box -8 -3 16 105
use FILL  FILL_2806
timestamp 1713400504
transform 1 0 824 0 1 1370
box -8 -3 16 105
use FILL  FILL_2807
timestamp 1713400504
transform 1 0 776 0 1 1370
box -8 -3 16 105
use FILL  FILL_2808
timestamp 1713400504
transform 1 0 768 0 1 1370
box -8 -3 16 105
use FILL  FILL_2809
timestamp 1713400504
transform 1 0 760 0 1 1370
box -8 -3 16 105
use FILL  FILL_2810
timestamp 1713400504
transform 1 0 752 0 1 1370
box -8 -3 16 105
use FILL  FILL_2811
timestamp 1713400504
transform 1 0 696 0 1 1370
box -8 -3 16 105
use FILL  FILL_2812
timestamp 1713400504
transform 1 0 688 0 1 1370
box -8 -3 16 105
use FILL  FILL_2813
timestamp 1713400504
transform 1 0 680 0 1 1370
box -8 -3 16 105
use FILL  FILL_2814
timestamp 1713400504
transform 1 0 672 0 1 1370
box -8 -3 16 105
use FILL  FILL_2815
timestamp 1713400504
transform 1 0 664 0 1 1370
box -8 -3 16 105
use FILL  FILL_2816
timestamp 1713400504
transform 1 0 656 0 1 1370
box -8 -3 16 105
use FILL  FILL_2817
timestamp 1713400504
transform 1 0 648 0 1 1370
box -8 -3 16 105
use FILL  FILL_2818
timestamp 1713400504
transform 1 0 640 0 1 1370
box -8 -3 16 105
use FILL  FILL_2819
timestamp 1713400504
transform 1 0 632 0 1 1370
box -8 -3 16 105
use FILL  FILL_2820
timestamp 1713400504
transform 1 0 576 0 1 1370
box -8 -3 16 105
use FILL  FILL_2821
timestamp 1713400504
transform 1 0 568 0 1 1370
box -8 -3 16 105
use FILL  FILL_2822
timestamp 1713400504
transform 1 0 560 0 1 1370
box -8 -3 16 105
use FILL  FILL_2823
timestamp 1713400504
transform 1 0 520 0 1 1370
box -8 -3 16 105
use FILL  FILL_2824
timestamp 1713400504
transform 1 0 512 0 1 1370
box -8 -3 16 105
use FILL  FILL_2825
timestamp 1713400504
transform 1 0 504 0 1 1370
box -8 -3 16 105
use FILL  FILL_2826
timestamp 1713400504
transform 1 0 496 0 1 1370
box -8 -3 16 105
use FILL  FILL_2827
timestamp 1713400504
transform 1 0 488 0 1 1370
box -8 -3 16 105
use FILL  FILL_2828
timestamp 1713400504
transform 1 0 480 0 1 1370
box -8 -3 16 105
use FILL  FILL_2829
timestamp 1713400504
transform 1 0 448 0 1 1370
box -8 -3 16 105
use FILL  FILL_2830
timestamp 1713400504
transform 1 0 440 0 1 1370
box -8 -3 16 105
use FILL  FILL_2831
timestamp 1713400504
transform 1 0 432 0 1 1370
box -8 -3 16 105
use FILL  FILL_2832
timestamp 1713400504
transform 1 0 424 0 1 1370
box -8 -3 16 105
use FILL  FILL_2833
timestamp 1713400504
transform 1 0 384 0 1 1370
box -8 -3 16 105
use FILL  FILL_2834
timestamp 1713400504
transform 1 0 376 0 1 1370
box -8 -3 16 105
use FILL  FILL_2835
timestamp 1713400504
transform 1 0 368 0 1 1370
box -8 -3 16 105
use FILL  FILL_2836
timestamp 1713400504
transform 1 0 360 0 1 1370
box -8 -3 16 105
use FILL  FILL_2837
timestamp 1713400504
transform 1 0 352 0 1 1370
box -8 -3 16 105
use FILL  FILL_2838
timestamp 1713400504
transform 1 0 344 0 1 1370
box -8 -3 16 105
use FILL  FILL_2839
timestamp 1713400504
transform 1 0 312 0 1 1370
box -8 -3 16 105
use FILL  FILL_2840
timestamp 1713400504
transform 1 0 304 0 1 1370
box -8 -3 16 105
use FILL  FILL_2841
timestamp 1713400504
transform 1 0 296 0 1 1370
box -8 -3 16 105
use FILL  FILL_2842
timestamp 1713400504
transform 1 0 288 0 1 1370
box -8 -3 16 105
use FILL  FILL_2843
timestamp 1713400504
transform 1 0 280 0 1 1370
box -8 -3 16 105
use FILL  FILL_2844
timestamp 1713400504
transform 1 0 240 0 1 1370
box -8 -3 16 105
use FILL  FILL_2845
timestamp 1713400504
transform 1 0 232 0 1 1370
box -8 -3 16 105
use FILL  FILL_2846
timestamp 1713400504
transform 1 0 224 0 1 1370
box -8 -3 16 105
use FILL  FILL_2847
timestamp 1713400504
transform 1 0 216 0 1 1370
box -8 -3 16 105
use FILL  FILL_2848
timestamp 1713400504
transform 1 0 192 0 1 1370
box -8 -3 16 105
use FILL  FILL_2849
timestamp 1713400504
transform 1 0 184 0 1 1370
box -8 -3 16 105
use FILL  FILL_2850
timestamp 1713400504
transform 1 0 176 0 1 1370
box -8 -3 16 105
use FILL  FILL_2851
timestamp 1713400504
transform 1 0 72 0 1 1370
box -8 -3 16 105
use FILL  FILL_2852
timestamp 1713400504
transform 1 0 2912 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2853
timestamp 1713400504
transform 1 0 2904 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2854
timestamp 1713400504
transform 1 0 2800 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2855
timestamp 1713400504
transform 1 0 2792 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2856
timestamp 1713400504
transform 1 0 2784 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2857
timestamp 1713400504
transform 1 0 2776 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2858
timestamp 1713400504
transform 1 0 2728 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2859
timestamp 1713400504
transform 1 0 2720 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2860
timestamp 1713400504
transform 1 0 2712 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2861
timestamp 1713400504
transform 1 0 2704 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2862
timestamp 1713400504
transform 1 0 2696 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2863
timestamp 1713400504
transform 1 0 2688 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2864
timestamp 1713400504
transform 1 0 2680 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2865
timestamp 1713400504
transform 1 0 2648 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2866
timestamp 1713400504
transform 1 0 2640 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2867
timestamp 1713400504
transform 1 0 2632 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2868
timestamp 1713400504
transform 1 0 2624 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2869
timestamp 1713400504
transform 1 0 2592 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2870
timestamp 1713400504
transform 1 0 2584 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2871
timestamp 1713400504
transform 1 0 2576 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2872
timestamp 1713400504
transform 1 0 2568 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2873
timestamp 1713400504
transform 1 0 2560 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2874
timestamp 1713400504
transform 1 0 2552 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2875
timestamp 1713400504
transform 1 0 2504 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2876
timestamp 1713400504
transform 1 0 2496 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2877
timestamp 1713400504
transform 1 0 2488 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2878
timestamp 1713400504
transform 1 0 2480 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2879
timestamp 1713400504
transform 1 0 2472 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2880
timestamp 1713400504
transform 1 0 2464 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2881
timestamp 1713400504
transform 1 0 2456 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2882
timestamp 1713400504
transform 1 0 2424 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2883
timestamp 1713400504
transform 1 0 2416 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2884
timestamp 1713400504
transform 1 0 2408 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2885
timestamp 1713400504
transform 1 0 2400 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2886
timestamp 1713400504
transform 1 0 2392 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2887
timestamp 1713400504
transform 1 0 2384 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2888
timestamp 1713400504
transform 1 0 2376 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2889
timestamp 1713400504
transform 1 0 2368 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2890
timestamp 1713400504
transform 1 0 2320 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2891
timestamp 1713400504
transform 1 0 2312 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2892
timestamp 1713400504
transform 1 0 2304 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2893
timestamp 1713400504
transform 1 0 2296 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2894
timestamp 1713400504
transform 1 0 2288 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2895
timestamp 1713400504
transform 1 0 2224 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2896
timestamp 1713400504
transform 1 0 2216 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2897
timestamp 1713400504
transform 1 0 2208 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2898
timestamp 1713400504
transform 1 0 2200 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2899
timestamp 1713400504
transform 1 0 2136 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2900
timestamp 1713400504
transform 1 0 2128 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2901
timestamp 1713400504
transform 1 0 2120 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2902
timestamp 1713400504
transform 1 0 2096 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2903
timestamp 1713400504
transform 1 0 2088 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2904
timestamp 1713400504
transform 1 0 2080 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2905
timestamp 1713400504
transform 1 0 2072 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2906
timestamp 1713400504
transform 1 0 2008 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2907
timestamp 1713400504
transform 1 0 2000 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2908
timestamp 1713400504
transform 1 0 1992 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2909
timestamp 1713400504
transform 1 0 1984 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2910
timestamp 1713400504
transform 1 0 1976 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2911
timestamp 1713400504
transform 1 0 1968 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2912
timestamp 1713400504
transform 1 0 1960 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2913
timestamp 1713400504
transform 1 0 1912 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2914
timestamp 1713400504
transform 1 0 1904 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2915
timestamp 1713400504
transform 1 0 1896 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2916
timestamp 1713400504
transform 1 0 1888 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2917
timestamp 1713400504
transform 1 0 1880 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2918
timestamp 1713400504
transform 1 0 1872 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2919
timestamp 1713400504
transform 1 0 1848 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2920
timestamp 1713400504
transform 1 0 1840 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2921
timestamp 1713400504
transform 1 0 1832 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2922
timestamp 1713400504
transform 1 0 1824 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2923
timestamp 1713400504
transform 1 0 1816 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2924
timestamp 1713400504
transform 1 0 1776 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2925
timestamp 1713400504
transform 1 0 1768 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2926
timestamp 1713400504
transform 1 0 1760 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2927
timestamp 1713400504
transform 1 0 1752 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2928
timestamp 1713400504
transform 1 0 1744 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2929
timestamp 1713400504
transform 1 0 1736 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2930
timestamp 1713400504
transform 1 0 1728 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2931
timestamp 1713400504
transform 1 0 1680 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2932
timestamp 1713400504
transform 1 0 1672 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2933
timestamp 1713400504
transform 1 0 1664 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2934
timestamp 1713400504
transform 1 0 1656 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2935
timestamp 1713400504
transform 1 0 1648 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2936
timestamp 1713400504
transform 1 0 1640 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2937
timestamp 1713400504
transform 1 0 1616 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2938
timestamp 1713400504
transform 1 0 1608 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2939
timestamp 1713400504
transform 1 0 1600 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2940
timestamp 1713400504
transform 1 0 1592 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2941
timestamp 1713400504
transform 1 0 1584 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2942
timestamp 1713400504
transform 1 0 1544 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2943
timestamp 1713400504
transform 1 0 1536 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2944
timestamp 1713400504
transform 1 0 1528 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2945
timestamp 1713400504
transform 1 0 1520 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2946
timestamp 1713400504
transform 1 0 1512 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2947
timestamp 1713400504
transform 1 0 1504 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2948
timestamp 1713400504
transform 1 0 1496 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2949
timestamp 1713400504
transform 1 0 1488 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2950
timestamp 1713400504
transform 1 0 1440 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2951
timestamp 1713400504
transform 1 0 1432 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2952
timestamp 1713400504
transform 1 0 1424 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2953
timestamp 1713400504
transform 1 0 1416 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2954
timestamp 1713400504
transform 1 0 1408 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2955
timestamp 1713400504
transform 1 0 1400 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2956
timestamp 1713400504
transform 1 0 1336 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2957
timestamp 1713400504
transform 1 0 1328 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2958
timestamp 1713400504
transform 1 0 1320 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2959
timestamp 1713400504
transform 1 0 1256 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2960
timestamp 1713400504
transform 1 0 1248 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2961
timestamp 1713400504
transform 1 0 1240 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2962
timestamp 1713400504
transform 1 0 1232 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2963
timestamp 1713400504
transform 1 0 1208 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2964
timestamp 1713400504
transform 1 0 1200 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2965
timestamp 1713400504
transform 1 0 1192 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2966
timestamp 1713400504
transform 1 0 1184 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2967
timestamp 1713400504
transform 1 0 1176 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2968
timestamp 1713400504
transform 1 0 1168 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2969
timestamp 1713400504
transform 1 0 1160 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2970
timestamp 1713400504
transform 1 0 1128 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2971
timestamp 1713400504
transform 1 0 1120 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2972
timestamp 1713400504
transform 1 0 1112 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2973
timestamp 1713400504
transform 1 0 1104 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2974
timestamp 1713400504
transform 1 0 1096 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2975
timestamp 1713400504
transform 1 0 1088 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2976
timestamp 1713400504
transform 1 0 1080 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2977
timestamp 1713400504
transform 1 0 1072 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2978
timestamp 1713400504
transform 1 0 1032 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2979
timestamp 1713400504
transform 1 0 1024 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2980
timestamp 1713400504
transform 1 0 1016 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2981
timestamp 1713400504
transform 1 0 1008 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2982
timestamp 1713400504
transform 1 0 1000 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2983
timestamp 1713400504
transform 1 0 992 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2984
timestamp 1713400504
transform 1 0 984 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2985
timestamp 1713400504
transform 1 0 976 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2986
timestamp 1713400504
transform 1 0 968 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2987
timestamp 1713400504
transform 1 0 920 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2988
timestamp 1713400504
transform 1 0 912 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2989
timestamp 1713400504
transform 1 0 904 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2990
timestamp 1713400504
transform 1 0 896 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2991
timestamp 1713400504
transform 1 0 888 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2992
timestamp 1713400504
transform 1 0 880 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2993
timestamp 1713400504
transform 1 0 872 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2994
timestamp 1713400504
transform 1 0 864 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2995
timestamp 1713400504
transform 1 0 856 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2996
timestamp 1713400504
transform 1 0 848 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2997
timestamp 1713400504
transform 1 0 800 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2998
timestamp 1713400504
transform 1 0 792 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2999
timestamp 1713400504
transform 1 0 784 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3000
timestamp 1713400504
transform 1 0 776 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3001
timestamp 1713400504
transform 1 0 768 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3002
timestamp 1713400504
transform 1 0 760 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3003
timestamp 1713400504
transform 1 0 752 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3004
timestamp 1713400504
transform 1 0 744 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3005
timestamp 1713400504
transform 1 0 736 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3006
timestamp 1713400504
transform 1 0 728 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3007
timestamp 1713400504
transform 1 0 720 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3008
timestamp 1713400504
transform 1 0 712 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3009
timestamp 1713400504
transform 1 0 608 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3010
timestamp 1713400504
transform 1 0 600 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3011
timestamp 1713400504
transform 1 0 592 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3012
timestamp 1713400504
transform 1 0 584 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3013
timestamp 1713400504
transform 1 0 576 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3014
timestamp 1713400504
transform 1 0 544 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3015
timestamp 1713400504
transform 1 0 536 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3016
timestamp 1713400504
transform 1 0 528 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3017
timestamp 1713400504
transform 1 0 504 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3018
timestamp 1713400504
transform 1 0 496 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3019
timestamp 1713400504
transform 1 0 488 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3020
timestamp 1713400504
transform 1 0 480 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3021
timestamp 1713400504
transform 1 0 472 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3022
timestamp 1713400504
transform 1 0 448 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3023
timestamp 1713400504
transform 1 0 440 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3024
timestamp 1713400504
transform 1 0 432 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3025
timestamp 1713400504
transform 1 0 400 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3026
timestamp 1713400504
transform 1 0 392 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3027
timestamp 1713400504
transform 1 0 384 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3028
timestamp 1713400504
transform 1 0 376 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3029
timestamp 1713400504
transform 1 0 368 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3030
timestamp 1713400504
transform 1 0 328 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3031
timestamp 1713400504
transform 1 0 320 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3032
timestamp 1713400504
transform 1 0 312 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3033
timestamp 1713400504
transform 1 0 304 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3034
timestamp 1713400504
transform 1 0 296 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3035
timestamp 1713400504
transform 1 0 288 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3036
timestamp 1713400504
transform 1 0 248 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3037
timestamp 1713400504
transform 1 0 240 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3038
timestamp 1713400504
transform 1 0 232 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3039
timestamp 1713400504
transform 1 0 208 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3040
timestamp 1713400504
transform 1 0 200 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3041
timestamp 1713400504
transform 1 0 192 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3042
timestamp 1713400504
transform 1 0 184 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3043
timestamp 1713400504
transform 1 0 144 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3044
timestamp 1713400504
transform 1 0 136 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3045
timestamp 1713400504
transform 1 0 128 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3046
timestamp 1713400504
transform 1 0 120 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3047
timestamp 1713400504
transform 1 0 112 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3048
timestamp 1713400504
transform 1 0 80 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3049
timestamp 1713400504
transform 1 0 72 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3050
timestamp 1713400504
transform 1 0 3008 0 1 1170
box -8 -3 16 105
use FILL  FILL_3051
timestamp 1713400504
transform 1 0 3000 0 1 1170
box -8 -3 16 105
use FILL  FILL_3052
timestamp 1713400504
transform 1 0 2992 0 1 1170
box -8 -3 16 105
use FILL  FILL_3053
timestamp 1713400504
transform 1 0 2904 0 1 1170
box -8 -3 16 105
use FILL  FILL_3054
timestamp 1713400504
transform 1 0 2896 0 1 1170
box -8 -3 16 105
use FILL  FILL_3055
timestamp 1713400504
transform 1 0 2888 0 1 1170
box -8 -3 16 105
use FILL  FILL_3056
timestamp 1713400504
transform 1 0 2880 0 1 1170
box -8 -3 16 105
use FILL  FILL_3057
timestamp 1713400504
transform 1 0 2872 0 1 1170
box -8 -3 16 105
use FILL  FILL_3058
timestamp 1713400504
transform 1 0 2824 0 1 1170
box -8 -3 16 105
use FILL  FILL_3059
timestamp 1713400504
transform 1 0 2816 0 1 1170
box -8 -3 16 105
use FILL  FILL_3060
timestamp 1713400504
transform 1 0 2808 0 1 1170
box -8 -3 16 105
use FILL  FILL_3061
timestamp 1713400504
transform 1 0 2800 0 1 1170
box -8 -3 16 105
use FILL  FILL_3062
timestamp 1713400504
transform 1 0 2776 0 1 1170
box -8 -3 16 105
use FILL  FILL_3063
timestamp 1713400504
transform 1 0 2768 0 1 1170
box -8 -3 16 105
use FILL  FILL_3064
timestamp 1713400504
transform 1 0 2568 0 1 1170
box -8 -3 16 105
use FILL  FILL_3065
timestamp 1713400504
transform 1 0 2560 0 1 1170
box -8 -3 16 105
use FILL  FILL_3066
timestamp 1713400504
transform 1 0 2552 0 1 1170
box -8 -3 16 105
use FILL  FILL_3067
timestamp 1713400504
transform 1 0 2512 0 1 1170
box -8 -3 16 105
use FILL  FILL_3068
timestamp 1713400504
transform 1 0 2504 0 1 1170
box -8 -3 16 105
use FILL  FILL_3069
timestamp 1713400504
transform 1 0 2480 0 1 1170
box -8 -3 16 105
use FILL  FILL_3070
timestamp 1713400504
transform 1 0 2472 0 1 1170
box -8 -3 16 105
use FILL  FILL_3071
timestamp 1713400504
transform 1 0 2464 0 1 1170
box -8 -3 16 105
use FILL  FILL_3072
timestamp 1713400504
transform 1 0 2456 0 1 1170
box -8 -3 16 105
use FILL  FILL_3073
timestamp 1713400504
transform 1 0 2448 0 1 1170
box -8 -3 16 105
use FILL  FILL_3074
timestamp 1713400504
transform 1 0 2440 0 1 1170
box -8 -3 16 105
use FILL  FILL_3075
timestamp 1713400504
transform 1 0 2392 0 1 1170
box -8 -3 16 105
use FILL  FILL_3076
timestamp 1713400504
transform 1 0 2384 0 1 1170
box -8 -3 16 105
use FILL  FILL_3077
timestamp 1713400504
transform 1 0 2376 0 1 1170
box -8 -3 16 105
use FILL  FILL_3078
timestamp 1713400504
transform 1 0 2256 0 1 1170
box -8 -3 16 105
use FILL  FILL_3079
timestamp 1713400504
transform 1 0 2248 0 1 1170
box -8 -3 16 105
use FILL  FILL_3080
timestamp 1713400504
transform 1 0 2240 0 1 1170
box -8 -3 16 105
use FILL  FILL_3081
timestamp 1713400504
transform 1 0 2232 0 1 1170
box -8 -3 16 105
use FILL  FILL_3082
timestamp 1713400504
transform 1 0 2184 0 1 1170
box -8 -3 16 105
use FILL  FILL_3083
timestamp 1713400504
transform 1 0 2176 0 1 1170
box -8 -3 16 105
use FILL  FILL_3084
timestamp 1713400504
transform 1 0 2168 0 1 1170
box -8 -3 16 105
use FILL  FILL_3085
timestamp 1713400504
transform 1 0 2048 0 1 1170
box -8 -3 16 105
use FILL  FILL_3086
timestamp 1713400504
transform 1 0 2040 0 1 1170
box -8 -3 16 105
use FILL  FILL_3087
timestamp 1713400504
transform 1 0 2032 0 1 1170
box -8 -3 16 105
use FILL  FILL_3088
timestamp 1713400504
transform 1 0 1984 0 1 1170
box -8 -3 16 105
use FILL  FILL_3089
timestamp 1713400504
transform 1 0 1976 0 1 1170
box -8 -3 16 105
use FILL  FILL_3090
timestamp 1713400504
transform 1 0 1968 0 1 1170
box -8 -3 16 105
use FILL  FILL_3091
timestamp 1713400504
transform 1 0 1960 0 1 1170
box -8 -3 16 105
use FILL  FILL_3092
timestamp 1713400504
transform 1 0 1952 0 1 1170
box -8 -3 16 105
use FILL  FILL_3093
timestamp 1713400504
transform 1 0 1944 0 1 1170
box -8 -3 16 105
use FILL  FILL_3094
timestamp 1713400504
transform 1 0 1896 0 1 1170
box -8 -3 16 105
use FILL  FILL_3095
timestamp 1713400504
transform 1 0 1888 0 1 1170
box -8 -3 16 105
use FILL  FILL_3096
timestamp 1713400504
transform 1 0 1880 0 1 1170
box -8 -3 16 105
use FILL  FILL_3097
timestamp 1713400504
transform 1 0 1872 0 1 1170
box -8 -3 16 105
use FILL  FILL_3098
timestamp 1713400504
transform 1 0 1864 0 1 1170
box -8 -3 16 105
use FILL  FILL_3099
timestamp 1713400504
transform 1 0 1856 0 1 1170
box -8 -3 16 105
use FILL  FILL_3100
timestamp 1713400504
transform 1 0 1824 0 1 1170
box -8 -3 16 105
use FILL  FILL_3101
timestamp 1713400504
transform 1 0 1816 0 1 1170
box -8 -3 16 105
use FILL  FILL_3102
timestamp 1713400504
transform 1 0 1808 0 1 1170
box -8 -3 16 105
use FILL  FILL_3103
timestamp 1713400504
transform 1 0 1776 0 1 1170
box -8 -3 16 105
use FILL  FILL_3104
timestamp 1713400504
transform 1 0 1768 0 1 1170
box -8 -3 16 105
use FILL  FILL_3105
timestamp 1713400504
transform 1 0 1760 0 1 1170
box -8 -3 16 105
use FILL  FILL_3106
timestamp 1713400504
transform 1 0 1752 0 1 1170
box -8 -3 16 105
use FILL  FILL_3107
timestamp 1713400504
transform 1 0 1728 0 1 1170
box -8 -3 16 105
use FILL  FILL_3108
timestamp 1713400504
transform 1 0 1720 0 1 1170
box -8 -3 16 105
use FILL  FILL_3109
timestamp 1713400504
transform 1 0 1712 0 1 1170
box -8 -3 16 105
use FILL  FILL_3110
timestamp 1713400504
transform 1 0 1704 0 1 1170
box -8 -3 16 105
use FILL  FILL_3111
timestamp 1713400504
transform 1 0 1696 0 1 1170
box -8 -3 16 105
use FILL  FILL_3112
timestamp 1713400504
transform 1 0 1656 0 1 1170
box -8 -3 16 105
use FILL  FILL_3113
timestamp 1713400504
transform 1 0 1648 0 1 1170
box -8 -3 16 105
use FILL  FILL_3114
timestamp 1713400504
transform 1 0 1640 0 1 1170
box -8 -3 16 105
use FILL  FILL_3115
timestamp 1713400504
transform 1 0 1632 0 1 1170
box -8 -3 16 105
use FILL  FILL_3116
timestamp 1713400504
transform 1 0 1624 0 1 1170
box -8 -3 16 105
use FILL  FILL_3117
timestamp 1713400504
transform 1 0 1616 0 1 1170
box -8 -3 16 105
use FILL  FILL_3118
timestamp 1713400504
transform 1 0 1608 0 1 1170
box -8 -3 16 105
use FILL  FILL_3119
timestamp 1713400504
transform 1 0 1560 0 1 1170
box -8 -3 16 105
use FILL  FILL_3120
timestamp 1713400504
transform 1 0 1552 0 1 1170
box -8 -3 16 105
use FILL  FILL_3121
timestamp 1713400504
transform 1 0 1544 0 1 1170
box -8 -3 16 105
use FILL  FILL_3122
timestamp 1713400504
transform 1 0 1536 0 1 1170
box -8 -3 16 105
use FILL  FILL_3123
timestamp 1713400504
transform 1 0 1528 0 1 1170
box -8 -3 16 105
use FILL  FILL_3124
timestamp 1713400504
transform 1 0 1520 0 1 1170
box -8 -3 16 105
use FILL  FILL_3125
timestamp 1713400504
transform 1 0 1512 0 1 1170
box -8 -3 16 105
use FILL  FILL_3126
timestamp 1713400504
transform 1 0 1504 0 1 1170
box -8 -3 16 105
use FILL  FILL_3127
timestamp 1713400504
transform 1 0 1456 0 1 1170
box -8 -3 16 105
use FILL  FILL_3128
timestamp 1713400504
transform 1 0 1448 0 1 1170
box -8 -3 16 105
use FILL  FILL_3129
timestamp 1713400504
transform 1 0 1440 0 1 1170
box -8 -3 16 105
use FILL  FILL_3130
timestamp 1713400504
transform 1 0 1432 0 1 1170
box -8 -3 16 105
use FILL  FILL_3131
timestamp 1713400504
transform 1 0 1424 0 1 1170
box -8 -3 16 105
use FILL  FILL_3132
timestamp 1713400504
transform 1 0 1416 0 1 1170
box -8 -3 16 105
use FILL  FILL_3133
timestamp 1713400504
transform 1 0 1408 0 1 1170
box -8 -3 16 105
use FILL  FILL_3134
timestamp 1713400504
transform 1 0 1368 0 1 1170
box -8 -3 16 105
use FILL  FILL_3135
timestamp 1713400504
transform 1 0 1360 0 1 1170
box -8 -3 16 105
use FILL  FILL_3136
timestamp 1713400504
transform 1 0 1352 0 1 1170
box -8 -3 16 105
use FILL  FILL_3137
timestamp 1713400504
transform 1 0 1344 0 1 1170
box -8 -3 16 105
use FILL  FILL_3138
timestamp 1713400504
transform 1 0 1336 0 1 1170
box -8 -3 16 105
use FILL  FILL_3139
timestamp 1713400504
transform 1 0 1296 0 1 1170
box -8 -3 16 105
use FILL  FILL_3140
timestamp 1713400504
transform 1 0 1288 0 1 1170
box -8 -3 16 105
use FILL  FILL_3141
timestamp 1713400504
transform 1 0 1280 0 1 1170
box -8 -3 16 105
use FILL  FILL_3142
timestamp 1713400504
transform 1 0 1272 0 1 1170
box -8 -3 16 105
use FILL  FILL_3143
timestamp 1713400504
transform 1 0 1264 0 1 1170
box -8 -3 16 105
use FILL  FILL_3144
timestamp 1713400504
transform 1 0 1256 0 1 1170
box -8 -3 16 105
use FILL  FILL_3145
timestamp 1713400504
transform 1 0 1248 0 1 1170
box -8 -3 16 105
use FILL  FILL_3146
timestamp 1713400504
transform 1 0 1200 0 1 1170
box -8 -3 16 105
use FILL  FILL_3147
timestamp 1713400504
transform 1 0 1192 0 1 1170
box -8 -3 16 105
use FILL  FILL_3148
timestamp 1713400504
transform 1 0 1184 0 1 1170
box -8 -3 16 105
use FILL  FILL_3149
timestamp 1713400504
transform 1 0 1176 0 1 1170
box -8 -3 16 105
use FILL  FILL_3150
timestamp 1713400504
transform 1 0 1168 0 1 1170
box -8 -3 16 105
use FILL  FILL_3151
timestamp 1713400504
transform 1 0 1160 0 1 1170
box -8 -3 16 105
use FILL  FILL_3152
timestamp 1713400504
transform 1 0 1152 0 1 1170
box -8 -3 16 105
use FILL  FILL_3153
timestamp 1713400504
transform 1 0 1112 0 1 1170
box -8 -3 16 105
use FILL  FILL_3154
timestamp 1713400504
transform 1 0 1104 0 1 1170
box -8 -3 16 105
use FILL  FILL_3155
timestamp 1713400504
transform 1 0 1096 0 1 1170
box -8 -3 16 105
use FILL  FILL_3156
timestamp 1713400504
transform 1 0 1088 0 1 1170
box -8 -3 16 105
use FILL  FILL_3157
timestamp 1713400504
transform 1 0 1080 0 1 1170
box -8 -3 16 105
use FILL  FILL_3158
timestamp 1713400504
transform 1 0 1072 0 1 1170
box -8 -3 16 105
use FILL  FILL_3159
timestamp 1713400504
transform 1 0 1064 0 1 1170
box -8 -3 16 105
use FILL  FILL_3160
timestamp 1713400504
transform 1 0 1024 0 1 1170
box -8 -3 16 105
use FILL  FILL_3161
timestamp 1713400504
transform 1 0 1016 0 1 1170
box -8 -3 16 105
use FILL  FILL_3162
timestamp 1713400504
transform 1 0 1008 0 1 1170
box -8 -3 16 105
use FILL  FILL_3163
timestamp 1713400504
transform 1 0 1000 0 1 1170
box -8 -3 16 105
use FILL  FILL_3164
timestamp 1713400504
transform 1 0 992 0 1 1170
box -8 -3 16 105
use FILL  FILL_3165
timestamp 1713400504
transform 1 0 984 0 1 1170
box -8 -3 16 105
use FILL  FILL_3166
timestamp 1713400504
transform 1 0 976 0 1 1170
box -8 -3 16 105
use FILL  FILL_3167
timestamp 1713400504
transform 1 0 944 0 1 1170
box -8 -3 16 105
use FILL  FILL_3168
timestamp 1713400504
transform 1 0 936 0 1 1170
box -8 -3 16 105
use FILL  FILL_3169
timestamp 1713400504
transform 1 0 928 0 1 1170
box -8 -3 16 105
use FILL  FILL_3170
timestamp 1713400504
transform 1 0 920 0 1 1170
box -8 -3 16 105
use FILL  FILL_3171
timestamp 1713400504
transform 1 0 912 0 1 1170
box -8 -3 16 105
use FILL  FILL_3172
timestamp 1713400504
transform 1 0 904 0 1 1170
box -8 -3 16 105
use FILL  FILL_3173
timestamp 1713400504
transform 1 0 896 0 1 1170
box -8 -3 16 105
use FILL  FILL_3174
timestamp 1713400504
transform 1 0 848 0 1 1170
box -8 -3 16 105
use FILL  FILL_3175
timestamp 1713400504
transform 1 0 840 0 1 1170
box -8 -3 16 105
use FILL  FILL_3176
timestamp 1713400504
transform 1 0 832 0 1 1170
box -8 -3 16 105
use FILL  FILL_3177
timestamp 1713400504
transform 1 0 824 0 1 1170
box -8 -3 16 105
use FILL  FILL_3178
timestamp 1713400504
transform 1 0 816 0 1 1170
box -8 -3 16 105
use FILL  FILL_3179
timestamp 1713400504
transform 1 0 808 0 1 1170
box -8 -3 16 105
use FILL  FILL_3180
timestamp 1713400504
transform 1 0 800 0 1 1170
box -8 -3 16 105
use FILL  FILL_3181
timestamp 1713400504
transform 1 0 792 0 1 1170
box -8 -3 16 105
use FILL  FILL_3182
timestamp 1713400504
transform 1 0 744 0 1 1170
box -8 -3 16 105
use FILL  FILL_3183
timestamp 1713400504
transform 1 0 736 0 1 1170
box -8 -3 16 105
use FILL  FILL_3184
timestamp 1713400504
transform 1 0 728 0 1 1170
box -8 -3 16 105
use FILL  FILL_3185
timestamp 1713400504
transform 1 0 720 0 1 1170
box -8 -3 16 105
use FILL  FILL_3186
timestamp 1713400504
transform 1 0 712 0 1 1170
box -8 -3 16 105
use FILL  FILL_3187
timestamp 1713400504
transform 1 0 704 0 1 1170
box -8 -3 16 105
use FILL  FILL_3188
timestamp 1713400504
transform 1 0 672 0 1 1170
box -8 -3 16 105
use FILL  FILL_3189
timestamp 1713400504
transform 1 0 664 0 1 1170
box -8 -3 16 105
use FILL  FILL_3190
timestamp 1713400504
transform 1 0 656 0 1 1170
box -8 -3 16 105
use FILL  FILL_3191
timestamp 1713400504
transform 1 0 648 0 1 1170
box -8 -3 16 105
use FILL  FILL_3192
timestamp 1713400504
transform 1 0 608 0 1 1170
box -8 -3 16 105
use FILL  FILL_3193
timestamp 1713400504
transform 1 0 600 0 1 1170
box -8 -3 16 105
use FILL  FILL_3194
timestamp 1713400504
transform 1 0 592 0 1 1170
box -8 -3 16 105
use FILL  FILL_3195
timestamp 1713400504
transform 1 0 584 0 1 1170
box -8 -3 16 105
use FILL  FILL_3196
timestamp 1713400504
transform 1 0 576 0 1 1170
box -8 -3 16 105
use FILL  FILL_3197
timestamp 1713400504
transform 1 0 568 0 1 1170
box -8 -3 16 105
use FILL  FILL_3198
timestamp 1713400504
transform 1 0 544 0 1 1170
box -8 -3 16 105
use FILL  FILL_3199
timestamp 1713400504
transform 1 0 536 0 1 1170
box -8 -3 16 105
use FILL  FILL_3200
timestamp 1713400504
transform 1 0 528 0 1 1170
box -8 -3 16 105
use FILL  FILL_3201
timestamp 1713400504
transform 1 0 488 0 1 1170
box -8 -3 16 105
use FILL  FILL_3202
timestamp 1713400504
transform 1 0 480 0 1 1170
box -8 -3 16 105
use FILL  FILL_3203
timestamp 1713400504
transform 1 0 472 0 1 1170
box -8 -3 16 105
use FILL  FILL_3204
timestamp 1713400504
transform 1 0 464 0 1 1170
box -8 -3 16 105
use FILL  FILL_3205
timestamp 1713400504
transform 1 0 456 0 1 1170
box -8 -3 16 105
use FILL  FILL_3206
timestamp 1713400504
transform 1 0 448 0 1 1170
box -8 -3 16 105
use FILL  FILL_3207
timestamp 1713400504
transform 1 0 408 0 1 1170
box -8 -3 16 105
use FILL  FILL_3208
timestamp 1713400504
transform 1 0 400 0 1 1170
box -8 -3 16 105
use FILL  FILL_3209
timestamp 1713400504
transform 1 0 392 0 1 1170
box -8 -3 16 105
use FILL  FILL_3210
timestamp 1713400504
transform 1 0 384 0 1 1170
box -8 -3 16 105
use FILL  FILL_3211
timestamp 1713400504
transform 1 0 376 0 1 1170
box -8 -3 16 105
use FILL  FILL_3212
timestamp 1713400504
transform 1 0 336 0 1 1170
box -8 -3 16 105
use FILL  FILL_3213
timestamp 1713400504
transform 1 0 328 0 1 1170
box -8 -3 16 105
use FILL  FILL_3214
timestamp 1713400504
transform 1 0 320 0 1 1170
box -8 -3 16 105
use FILL  FILL_3215
timestamp 1713400504
transform 1 0 312 0 1 1170
box -8 -3 16 105
use FILL  FILL_3216
timestamp 1713400504
transform 1 0 304 0 1 1170
box -8 -3 16 105
use FILL  FILL_3217
timestamp 1713400504
transform 1 0 280 0 1 1170
box -8 -3 16 105
use FILL  FILL_3218
timestamp 1713400504
transform 1 0 272 0 1 1170
box -8 -3 16 105
use FILL  FILL_3219
timestamp 1713400504
transform 1 0 264 0 1 1170
box -8 -3 16 105
use FILL  FILL_3220
timestamp 1713400504
transform 1 0 224 0 1 1170
box -8 -3 16 105
use FILL  FILL_3221
timestamp 1713400504
transform 1 0 216 0 1 1170
box -8 -3 16 105
use FILL  FILL_3222
timestamp 1713400504
transform 1 0 208 0 1 1170
box -8 -3 16 105
use FILL  FILL_3223
timestamp 1713400504
transform 1 0 200 0 1 1170
box -8 -3 16 105
use FILL  FILL_3224
timestamp 1713400504
transform 1 0 192 0 1 1170
box -8 -3 16 105
use FILL  FILL_3225
timestamp 1713400504
transform 1 0 168 0 1 1170
box -8 -3 16 105
use FILL  FILL_3226
timestamp 1713400504
transform 1 0 160 0 1 1170
box -8 -3 16 105
use FILL  FILL_3227
timestamp 1713400504
transform 1 0 152 0 1 1170
box -8 -3 16 105
use FILL  FILL_3228
timestamp 1713400504
transform 1 0 144 0 1 1170
box -8 -3 16 105
use FILL  FILL_3229
timestamp 1713400504
transform 1 0 112 0 1 1170
box -8 -3 16 105
use FILL  FILL_3230
timestamp 1713400504
transform 1 0 104 0 1 1170
box -8 -3 16 105
use FILL  FILL_3231
timestamp 1713400504
transform 1 0 96 0 1 1170
box -8 -3 16 105
use FILL  FILL_3232
timestamp 1713400504
transform 1 0 88 0 1 1170
box -8 -3 16 105
use FILL  FILL_3233
timestamp 1713400504
transform 1 0 80 0 1 1170
box -8 -3 16 105
use FILL  FILL_3234
timestamp 1713400504
transform 1 0 72 0 1 1170
box -8 -3 16 105
use FILL  FILL_3235
timestamp 1713400504
transform 1 0 2912 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3236
timestamp 1713400504
transform 1 0 2904 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3237
timestamp 1713400504
transform 1 0 2800 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3238
timestamp 1713400504
transform 1 0 2792 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3239
timestamp 1713400504
transform 1 0 2784 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3240
timestamp 1713400504
transform 1 0 2776 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3241
timestamp 1713400504
transform 1 0 2768 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3242
timestamp 1713400504
transform 1 0 2720 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3243
timestamp 1713400504
transform 1 0 2712 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3244
timestamp 1713400504
transform 1 0 2704 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3245
timestamp 1713400504
transform 1 0 2696 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3246
timestamp 1713400504
transform 1 0 2688 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3247
timestamp 1713400504
transform 1 0 2680 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3248
timestamp 1713400504
transform 1 0 2672 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3249
timestamp 1713400504
transform 1 0 2648 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3250
timestamp 1713400504
transform 1 0 2640 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3251
timestamp 1713400504
transform 1 0 2632 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3252
timestamp 1713400504
transform 1 0 2624 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3253
timestamp 1713400504
transform 1 0 2584 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3254
timestamp 1713400504
transform 1 0 2576 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3255
timestamp 1713400504
transform 1 0 2568 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3256
timestamp 1713400504
transform 1 0 2560 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3257
timestamp 1713400504
transform 1 0 2552 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3258
timestamp 1713400504
transform 1 0 2544 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3259
timestamp 1713400504
transform 1 0 2504 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3260
timestamp 1713400504
transform 1 0 2496 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3261
timestamp 1713400504
transform 1 0 2488 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3262
timestamp 1713400504
transform 1 0 2480 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3263
timestamp 1713400504
transform 1 0 2472 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3264
timestamp 1713400504
transform 1 0 2464 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3265
timestamp 1713400504
transform 1 0 2424 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3266
timestamp 1713400504
transform 1 0 2416 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3267
timestamp 1713400504
transform 1 0 2408 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3268
timestamp 1713400504
transform 1 0 2400 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3269
timestamp 1713400504
transform 1 0 2392 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3270
timestamp 1713400504
transform 1 0 2368 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3271
timestamp 1713400504
transform 1 0 2360 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3272
timestamp 1713400504
transform 1 0 2352 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3273
timestamp 1713400504
transform 1 0 2344 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3274
timestamp 1713400504
transform 1 0 2280 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3275
timestamp 1713400504
transform 1 0 2216 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3276
timestamp 1713400504
transform 1 0 2208 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3277
timestamp 1713400504
transform 1 0 2200 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3278
timestamp 1713400504
transform 1 0 2192 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3279
timestamp 1713400504
transform 1 0 2184 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3280
timestamp 1713400504
transform 1 0 2136 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3281
timestamp 1713400504
transform 1 0 2128 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3282
timestamp 1713400504
transform 1 0 2120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3283
timestamp 1713400504
transform 1 0 2112 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3284
timestamp 1713400504
transform 1 0 2104 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3285
timestamp 1713400504
transform 1 0 1984 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3286
timestamp 1713400504
transform 1 0 1976 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3287
timestamp 1713400504
transform 1 0 1968 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3288
timestamp 1713400504
transform 1 0 1960 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3289
timestamp 1713400504
transform 1 0 1952 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3290
timestamp 1713400504
transform 1 0 1904 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3291
timestamp 1713400504
transform 1 0 1896 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3292
timestamp 1713400504
transform 1 0 1888 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3293
timestamp 1713400504
transform 1 0 1880 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3294
timestamp 1713400504
transform 1 0 1872 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3295
timestamp 1713400504
transform 1 0 1864 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3296
timestamp 1713400504
transform 1 0 1856 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3297
timestamp 1713400504
transform 1 0 1848 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3298
timestamp 1713400504
transform 1 0 1816 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3299
timestamp 1713400504
transform 1 0 1792 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3300
timestamp 1713400504
transform 1 0 1784 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3301
timestamp 1713400504
transform 1 0 1776 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3302
timestamp 1713400504
transform 1 0 1768 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3303
timestamp 1713400504
transform 1 0 1760 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3304
timestamp 1713400504
transform 1 0 1752 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3305
timestamp 1713400504
transform 1 0 1744 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3306
timestamp 1713400504
transform 1 0 1696 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3307
timestamp 1713400504
transform 1 0 1688 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3308
timestamp 1713400504
transform 1 0 1680 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3309
timestamp 1713400504
transform 1 0 1672 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3310
timestamp 1713400504
transform 1 0 1664 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3311
timestamp 1713400504
transform 1 0 1656 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3312
timestamp 1713400504
transform 1 0 1648 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3313
timestamp 1713400504
transform 1 0 1640 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3314
timestamp 1713400504
transform 1 0 1592 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3315
timestamp 1713400504
transform 1 0 1584 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3316
timestamp 1713400504
transform 1 0 1576 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3317
timestamp 1713400504
transform 1 0 1568 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3318
timestamp 1713400504
transform 1 0 1560 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3319
timestamp 1713400504
transform 1 0 1552 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3320
timestamp 1713400504
transform 1 0 1544 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3321
timestamp 1713400504
transform 1 0 1536 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3322
timestamp 1713400504
transform 1 0 1496 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3323
timestamp 1713400504
transform 1 0 1488 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3324
timestamp 1713400504
transform 1 0 1480 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3325
timestamp 1713400504
transform 1 0 1472 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3326
timestamp 1713400504
transform 1 0 1464 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3327
timestamp 1713400504
transform 1 0 1456 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3328
timestamp 1713400504
transform 1 0 1448 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3329
timestamp 1713400504
transform 1 0 1440 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3330
timestamp 1713400504
transform 1 0 1408 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3331
timestamp 1713400504
transform 1 0 1400 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3332
timestamp 1713400504
transform 1 0 1392 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3333
timestamp 1713400504
transform 1 0 1384 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3334
timestamp 1713400504
transform 1 0 1376 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3335
timestamp 1713400504
transform 1 0 1368 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3336
timestamp 1713400504
transform 1 0 1360 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3337
timestamp 1713400504
transform 1 0 1352 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3338
timestamp 1713400504
transform 1 0 1344 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3339
timestamp 1713400504
transform 1 0 1296 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3340
timestamp 1713400504
transform 1 0 1288 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3341
timestamp 1713400504
transform 1 0 1280 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3342
timestamp 1713400504
transform 1 0 1272 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3343
timestamp 1713400504
transform 1 0 1264 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3344
timestamp 1713400504
transform 1 0 1256 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3345
timestamp 1713400504
transform 1 0 1248 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3346
timestamp 1713400504
transform 1 0 1240 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3347
timestamp 1713400504
transform 1 0 1232 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3348
timestamp 1713400504
transform 1 0 1224 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3349
timestamp 1713400504
transform 1 0 1216 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3350
timestamp 1713400504
transform 1 0 1208 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3351
timestamp 1713400504
transform 1 0 1200 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3352
timestamp 1713400504
transform 1 0 1192 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3353
timestamp 1713400504
transform 1 0 1184 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3354
timestamp 1713400504
transform 1 0 1176 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3355
timestamp 1713400504
transform 1 0 1128 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3356
timestamp 1713400504
transform 1 0 1120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3357
timestamp 1713400504
transform 1 0 1112 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3358
timestamp 1713400504
transform 1 0 1104 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3359
timestamp 1713400504
transform 1 0 1096 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3360
timestamp 1713400504
transform 1 0 1088 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3361
timestamp 1713400504
transform 1 0 1080 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3362
timestamp 1713400504
transform 1 0 1072 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3363
timestamp 1713400504
transform 1 0 1064 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3364
timestamp 1713400504
transform 1 0 1040 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3365
timestamp 1713400504
transform 1 0 1032 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3366
timestamp 1713400504
transform 1 0 1024 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3367
timestamp 1713400504
transform 1 0 1016 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3368
timestamp 1713400504
transform 1 0 1008 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3369
timestamp 1713400504
transform 1 0 1000 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3370
timestamp 1713400504
transform 1 0 992 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3371
timestamp 1713400504
transform 1 0 984 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3372
timestamp 1713400504
transform 1 0 976 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3373
timestamp 1713400504
transform 1 0 968 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3374
timestamp 1713400504
transform 1 0 928 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3375
timestamp 1713400504
transform 1 0 920 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3376
timestamp 1713400504
transform 1 0 912 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3377
timestamp 1713400504
transform 1 0 904 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3378
timestamp 1713400504
transform 1 0 896 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3379
timestamp 1713400504
transform 1 0 888 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3380
timestamp 1713400504
transform 1 0 784 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3381
timestamp 1713400504
transform 1 0 776 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3382
timestamp 1713400504
transform 1 0 768 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3383
timestamp 1713400504
transform 1 0 760 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3384
timestamp 1713400504
transform 1 0 720 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3385
timestamp 1713400504
transform 1 0 712 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3386
timestamp 1713400504
transform 1 0 704 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3387
timestamp 1713400504
transform 1 0 696 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3388
timestamp 1713400504
transform 1 0 688 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3389
timestamp 1713400504
transform 1 0 680 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3390
timestamp 1713400504
transform 1 0 672 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3391
timestamp 1713400504
transform 1 0 640 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3392
timestamp 1713400504
transform 1 0 632 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3393
timestamp 1713400504
transform 1 0 624 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3394
timestamp 1713400504
transform 1 0 616 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3395
timestamp 1713400504
transform 1 0 608 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3396
timestamp 1713400504
transform 1 0 584 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3397
timestamp 1713400504
transform 1 0 576 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3398
timestamp 1713400504
transform 1 0 568 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3399
timestamp 1713400504
transform 1 0 544 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3400
timestamp 1713400504
transform 1 0 536 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3401
timestamp 1713400504
transform 1 0 528 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3402
timestamp 1713400504
transform 1 0 520 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3403
timestamp 1713400504
transform 1 0 480 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3404
timestamp 1713400504
transform 1 0 472 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3405
timestamp 1713400504
transform 1 0 464 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3406
timestamp 1713400504
transform 1 0 456 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3407
timestamp 1713400504
transform 1 0 448 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3408
timestamp 1713400504
transform 1 0 440 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3409
timestamp 1713400504
transform 1 0 400 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3410
timestamp 1713400504
transform 1 0 392 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3411
timestamp 1713400504
transform 1 0 384 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3412
timestamp 1713400504
transform 1 0 360 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3413
timestamp 1713400504
transform 1 0 352 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3414
timestamp 1713400504
transform 1 0 344 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3415
timestamp 1713400504
transform 1 0 336 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3416
timestamp 1713400504
transform 1 0 296 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3417
timestamp 1713400504
transform 1 0 288 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3418
timestamp 1713400504
transform 1 0 280 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3419
timestamp 1713400504
transform 1 0 272 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3420
timestamp 1713400504
transform 1 0 264 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3421
timestamp 1713400504
transform 1 0 240 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3422
timestamp 1713400504
transform 1 0 232 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3423
timestamp 1713400504
transform 1 0 224 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3424
timestamp 1713400504
transform 1 0 192 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3425
timestamp 1713400504
transform 1 0 184 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3426
timestamp 1713400504
transform 1 0 176 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3427
timestamp 1713400504
transform 1 0 168 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3428
timestamp 1713400504
transform 1 0 160 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3429
timestamp 1713400504
transform 1 0 152 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3430
timestamp 1713400504
transform 1 0 120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3431
timestamp 1713400504
transform 1 0 112 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3432
timestamp 1713400504
transform 1 0 88 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3433
timestamp 1713400504
transform 1 0 80 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3434
timestamp 1713400504
transform 1 0 72 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3435
timestamp 1713400504
transform 1 0 2912 0 1 970
box -8 -3 16 105
use FILL  FILL_3436
timestamp 1713400504
transform 1 0 2808 0 1 970
box -8 -3 16 105
use FILL  FILL_3437
timestamp 1713400504
transform 1 0 2800 0 1 970
box -8 -3 16 105
use FILL  FILL_3438
timestamp 1713400504
transform 1 0 2792 0 1 970
box -8 -3 16 105
use FILL  FILL_3439
timestamp 1713400504
transform 1 0 2744 0 1 970
box -8 -3 16 105
use FILL  FILL_3440
timestamp 1713400504
transform 1 0 2736 0 1 970
box -8 -3 16 105
use FILL  FILL_3441
timestamp 1713400504
transform 1 0 2520 0 1 970
box -8 -3 16 105
use FILL  FILL_3442
timestamp 1713400504
transform 1 0 2512 0 1 970
box -8 -3 16 105
use FILL  FILL_3443
timestamp 1713400504
transform 1 0 2472 0 1 970
box -8 -3 16 105
use FILL  FILL_3444
timestamp 1713400504
transform 1 0 2464 0 1 970
box -8 -3 16 105
use FILL  FILL_3445
timestamp 1713400504
transform 1 0 2456 0 1 970
box -8 -3 16 105
use FILL  FILL_3446
timestamp 1713400504
transform 1 0 2416 0 1 970
box -8 -3 16 105
use FILL  FILL_3447
timestamp 1713400504
transform 1 0 2408 0 1 970
box -8 -3 16 105
use FILL  FILL_3448
timestamp 1713400504
transform 1 0 2400 0 1 970
box -8 -3 16 105
use FILL  FILL_3449
timestamp 1713400504
transform 1 0 2392 0 1 970
box -8 -3 16 105
use FILL  FILL_3450
timestamp 1713400504
transform 1 0 2384 0 1 970
box -8 -3 16 105
use FILL  FILL_3451
timestamp 1713400504
transform 1 0 2376 0 1 970
box -8 -3 16 105
use FILL  FILL_3452
timestamp 1713400504
transform 1 0 2336 0 1 970
box -8 -3 16 105
use FILL  FILL_3453
timestamp 1713400504
transform 1 0 2328 0 1 970
box -8 -3 16 105
use FILL  FILL_3454
timestamp 1713400504
transform 1 0 2320 0 1 970
box -8 -3 16 105
use FILL  FILL_3455
timestamp 1713400504
transform 1 0 2256 0 1 970
box -8 -3 16 105
use FILL  FILL_3456
timestamp 1713400504
transform 1 0 2248 0 1 970
box -8 -3 16 105
use FILL  FILL_3457
timestamp 1713400504
transform 1 0 2240 0 1 970
box -8 -3 16 105
use FILL  FILL_3458
timestamp 1713400504
transform 1 0 2232 0 1 970
box -8 -3 16 105
use FILL  FILL_3459
timestamp 1713400504
transform 1 0 2208 0 1 970
box -8 -3 16 105
use FILL  FILL_3460
timestamp 1713400504
transform 1 0 2200 0 1 970
box -8 -3 16 105
use FILL  FILL_3461
timestamp 1713400504
transform 1 0 2192 0 1 970
box -8 -3 16 105
use FILL  FILL_3462
timestamp 1713400504
transform 1 0 2168 0 1 970
box -8 -3 16 105
use FILL  FILL_3463
timestamp 1713400504
transform 1 0 2160 0 1 970
box -8 -3 16 105
use FILL  FILL_3464
timestamp 1713400504
transform 1 0 2152 0 1 970
box -8 -3 16 105
use FILL  FILL_3465
timestamp 1713400504
transform 1 0 2144 0 1 970
box -8 -3 16 105
use FILL  FILL_3466
timestamp 1713400504
transform 1 0 2080 0 1 970
box -8 -3 16 105
use FILL  FILL_3467
timestamp 1713400504
transform 1 0 2072 0 1 970
box -8 -3 16 105
use FILL  FILL_3468
timestamp 1713400504
transform 1 0 2064 0 1 970
box -8 -3 16 105
use FILL  FILL_3469
timestamp 1713400504
transform 1 0 2056 0 1 970
box -8 -3 16 105
use FILL  FILL_3470
timestamp 1713400504
transform 1 0 2032 0 1 970
box -8 -3 16 105
use FILL  FILL_3471
timestamp 1713400504
transform 1 0 2024 0 1 970
box -8 -3 16 105
use FILL  FILL_3472
timestamp 1713400504
transform 1 0 2016 0 1 970
box -8 -3 16 105
use FILL  FILL_3473
timestamp 1713400504
transform 1 0 2008 0 1 970
box -8 -3 16 105
use FILL  FILL_3474
timestamp 1713400504
transform 1 0 1944 0 1 970
box -8 -3 16 105
use FILL  FILL_3475
timestamp 1713400504
transform 1 0 1936 0 1 970
box -8 -3 16 105
use FILL  FILL_3476
timestamp 1713400504
transform 1 0 1928 0 1 970
box -8 -3 16 105
use FILL  FILL_3477
timestamp 1713400504
transform 1 0 1920 0 1 970
box -8 -3 16 105
use FILL  FILL_3478
timestamp 1713400504
transform 1 0 1912 0 1 970
box -8 -3 16 105
use FILL  FILL_3479
timestamp 1713400504
transform 1 0 1904 0 1 970
box -8 -3 16 105
use FILL  FILL_3480
timestamp 1713400504
transform 1 0 1856 0 1 970
box -8 -3 16 105
use FILL  FILL_3481
timestamp 1713400504
transform 1 0 1848 0 1 970
box -8 -3 16 105
use FILL  FILL_3482
timestamp 1713400504
transform 1 0 1840 0 1 970
box -8 -3 16 105
use FILL  FILL_3483
timestamp 1713400504
transform 1 0 1832 0 1 970
box -8 -3 16 105
use FILL  FILL_3484
timestamp 1713400504
transform 1 0 1824 0 1 970
box -8 -3 16 105
use FILL  FILL_3485
timestamp 1713400504
transform 1 0 1800 0 1 970
box -8 -3 16 105
use FILL  FILL_3486
timestamp 1713400504
transform 1 0 1792 0 1 970
box -8 -3 16 105
use FILL  FILL_3487
timestamp 1713400504
transform 1 0 1784 0 1 970
box -8 -3 16 105
use FILL  FILL_3488
timestamp 1713400504
transform 1 0 1776 0 1 970
box -8 -3 16 105
use FILL  FILL_3489
timestamp 1713400504
transform 1 0 1768 0 1 970
box -8 -3 16 105
use FILL  FILL_3490
timestamp 1713400504
transform 1 0 1728 0 1 970
box -8 -3 16 105
use FILL  FILL_3491
timestamp 1713400504
transform 1 0 1720 0 1 970
box -8 -3 16 105
use FILL  FILL_3492
timestamp 1713400504
transform 1 0 1712 0 1 970
box -8 -3 16 105
use FILL  FILL_3493
timestamp 1713400504
transform 1 0 1704 0 1 970
box -8 -3 16 105
use FILL  FILL_3494
timestamp 1713400504
transform 1 0 1696 0 1 970
box -8 -3 16 105
use FILL  FILL_3495
timestamp 1713400504
transform 1 0 1656 0 1 970
box -8 -3 16 105
use FILL  FILL_3496
timestamp 1713400504
transform 1 0 1648 0 1 970
box -8 -3 16 105
use FILL  FILL_3497
timestamp 1713400504
transform 1 0 1640 0 1 970
box -8 -3 16 105
use FILL  FILL_3498
timestamp 1713400504
transform 1 0 1632 0 1 970
box -8 -3 16 105
use FILL  FILL_3499
timestamp 1713400504
transform 1 0 1624 0 1 970
box -8 -3 16 105
use FILL  FILL_3500
timestamp 1713400504
transform 1 0 1616 0 1 970
box -8 -3 16 105
use FILL  FILL_3501
timestamp 1713400504
transform 1 0 1568 0 1 970
box -8 -3 16 105
use FILL  FILL_3502
timestamp 1713400504
transform 1 0 1560 0 1 970
box -8 -3 16 105
use FILL  FILL_3503
timestamp 1713400504
transform 1 0 1552 0 1 970
box -8 -3 16 105
use FILL  FILL_3504
timestamp 1713400504
transform 1 0 1544 0 1 970
box -8 -3 16 105
use FILL  FILL_3505
timestamp 1713400504
transform 1 0 1536 0 1 970
box -8 -3 16 105
use FILL  FILL_3506
timestamp 1713400504
transform 1 0 1528 0 1 970
box -8 -3 16 105
use FILL  FILL_3507
timestamp 1713400504
transform 1 0 1520 0 1 970
box -8 -3 16 105
use FILL  FILL_3508
timestamp 1713400504
transform 1 0 1512 0 1 970
box -8 -3 16 105
use FILL  FILL_3509
timestamp 1713400504
transform 1 0 1504 0 1 970
box -8 -3 16 105
use FILL  FILL_3510
timestamp 1713400504
transform 1 0 1456 0 1 970
box -8 -3 16 105
use FILL  FILL_3511
timestamp 1713400504
transform 1 0 1448 0 1 970
box -8 -3 16 105
use FILL  FILL_3512
timestamp 1713400504
transform 1 0 1440 0 1 970
box -8 -3 16 105
use FILL  FILL_3513
timestamp 1713400504
transform 1 0 1432 0 1 970
box -8 -3 16 105
use FILL  FILL_3514
timestamp 1713400504
transform 1 0 1424 0 1 970
box -8 -3 16 105
use FILL  FILL_3515
timestamp 1713400504
transform 1 0 1416 0 1 970
box -8 -3 16 105
use FILL  FILL_3516
timestamp 1713400504
transform 1 0 1408 0 1 970
box -8 -3 16 105
use FILL  FILL_3517
timestamp 1713400504
transform 1 0 1400 0 1 970
box -8 -3 16 105
use FILL  FILL_3518
timestamp 1713400504
transform 1 0 1392 0 1 970
box -8 -3 16 105
use FILL  FILL_3519
timestamp 1713400504
transform 1 0 1344 0 1 970
box -8 -3 16 105
use FILL  FILL_3520
timestamp 1713400504
transform 1 0 1336 0 1 970
box -8 -3 16 105
use FILL  FILL_3521
timestamp 1713400504
transform 1 0 1328 0 1 970
box -8 -3 16 105
use FILL  FILL_3522
timestamp 1713400504
transform 1 0 1320 0 1 970
box -8 -3 16 105
use FILL  FILL_3523
timestamp 1713400504
transform 1 0 1312 0 1 970
box -8 -3 16 105
use FILL  FILL_3524
timestamp 1713400504
transform 1 0 1304 0 1 970
box -8 -3 16 105
use FILL  FILL_3525
timestamp 1713400504
transform 1 0 1296 0 1 970
box -8 -3 16 105
use FILL  FILL_3526
timestamp 1713400504
transform 1 0 1288 0 1 970
box -8 -3 16 105
use FILL  FILL_3527
timestamp 1713400504
transform 1 0 1280 0 1 970
box -8 -3 16 105
use FILL  FILL_3528
timestamp 1713400504
transform 1 0 1232 0 1 970
box -8 -3 16 105
use FILL  FILL_3529
timestamp 1713400504
transform 1 0 1224 0 1 970
box -8 -3 16 105
use FILL  FILL_3530
timestamp 1713400504
transform 1 0 1216 0 1 970
box -8 -3 16 105
use FILL  FILL_3531
timestamp 1713400504
transform 1 0 1208 0 1 970
box -8 -3 16 105
use FILL  FILL_3532
timestamp 1713400504
transform 1 0 1200 0 1 970
box -8 -3 16 105
use FILL  FILL_3533
timestamp 1713400504
transform 1 0 1192 0 1 970
box -8 -3 16 105
use FILL  FILL_3534
timestamp 1713400504
transform 1 0 1184 0 1 970
box -8 -3 16 105
use FILL  FILL_3535
timestamp 1713400504
transform 1 0 1176 0 1 970
box -8 -3 16 105
use FILL  FILL_3536
timestamp 1713400504
transform 1 0 1168 0 1 970
box -8 -3 16 105
use FILL  FILL_3537
timestamp 1713400504
transform 1 0 1128 0 1 970
box -8 -3 16 105
use FILL  FILL_3538
timestamp 1713400504
transform 1 0 1120 0 1 970
box -8 -3 16 105
use FILL  FILL_3539
timestamp 1713400504
transform 1 0 1112 0 1 970
box -8 -3 16 105
use FILL  FILL_3540
timestamp 1713400504
transform 1 0 1104 0 1 970
box -8 -3 16 105
use FILL  FILL_3541
timestamp 1713400504
transform 1 0 1096 0 1 970
box -8 -3 16 105
use FILL  FILL_3542
timestamp 1713400504
transform 1 0 1088 0 1 970
box -8 -3 16 105
use FILL  FILL_3543
timestamp 1713400504
transform 1 0 1080 0 1 970
box -8 -3 16 105
use FILL  FILL_3544
timestamp 1713400504
transform 1 0 1072 0 1 970
box -8 -3 16 105
use FILL  FILL_3545
timestamp 1713400504
transform 1 0 1032 0 1 970
box -8 -3 16 105
use FILL  FILL_3546
timestamp 1713400504
transform 1 0 1024 0 1 970
box -8 -3 16 105
use FILL  FILL_3547
timestamp 1713400504
transform 1 0 1016 0 1 970
box -8 -3 16 105
use FILL  FILL_3548
timestamp 1713400504
transform 1 0 1008 0 1 970
box -8 -3 16 105
use FILL  FILL_3549
timestamp 1713400504
transform 1 0 1000 0 1 970
box -8 -3 16 105
use FILL  FILL_3550
timestamp 1713400504
transform 1 0 992 0 1 970
box -8 -3 16 105
use FILL  FILL_3551
timestamp 1713400504
transform 1 0 984 0 1 970
box -8 -3 16 105
use FILL  FILL_3552
timestamp 1713400504
transform 1 0 976 0 1 970
box -8 -3 16 105
use FILL  FILL_3553
timestamp 1713400504
transform 1 0 936 0 1 970
box -8 -3 16 105
use FILL  FILL_3554
timestamp 1713400504
transform 1 0 928 0 1 970
box -8 -3 16 105
use FILL  FILL_3555
timestamp 1713400504
transform 1 0 920 0 1 970
box -8 -3 16 105
use FILL  FILL_3556
timestamp 1713400504
transform 1 0 912 0 1 970
box -8 -3 16 105
use FILL  FILL_3557
timestamp 1713400504
transform 1 0 904 0 1 970
box -8 -3 16 105
use FILL  FILL_3558
timestamp 1713400504
transform 1 0 896 0 1 970
box -8 -3 16 105
use FILL  FILL_3559
timestamp 1713400504
transform 1 0 888 0 1 970
box -8 -3 16 105
use FILL  FILL_3560
timestamp 1713400504
transform 1 0 840 0 1 970
box -8 -3 16 105
use FILL  FILL_3561
timestamp 1713400504
transform 1 0 832 0 1 970
box -8 -3 16 105
use FILL  FILL_3562
timestamp 1713400504
transform 1 0 824 0 1 970
box -8 -3 16 105
use FILL  FILL_3563
timestamp 1713400504
transform 1 0 816 0 1 970
box -8 -3 16 105
use FILL  FILL_3564
timestamp 1713400504
transform 1 0 808 0 1 970
box -8 -3 16 105
use FILL  FILL_3565
timestamp 1713400504
transform 1 0 800 0 1 970
box -8 -3 16 105
use FILL  FILL_3566
timestamp 1713400504
transform 1 0 792 0 1 970
box -8 -3 16 105
use FILL  FILL_3567
timestamp 1713400504
transform 1 0 784 0 1 970
box -8 -3 16 105
use FILL  FILL_3568
timestamp 1713400504
transform 1 0 736 0 1 970
box -8 -3 16 105
use FILL  FILL_3569
timestamp 1713400504
transform 1 0 728 0 1 970
box -8 -3 16 105
use FILL  FILL_3570
timestamp 1713400504
transform 1 0 720 0 1 970
box -8 -3 16 105
use FILL  FILL_3571
timestamp 1713400504
transform 1 0 712 0 1 970
box -8 -3 16 105
use FILL  FILL_3572
timestamp 1713400504
transform 1 0 704 0 1 970
box -8 -3 16 105
use FILL  FILL_3573
timestamp 1713400504
transform 1 0 696 0 1 970
box -8 -3 16 105
use FILL  FILL_3574
timestamp 1713400504
transform 1 0 592 0 1 970
box -8 -3 16 105
use FILL  FILL_3575
timestamp 1713400504
transform 1 0 584 0 1 970
box -8 -3 16 105
use FILL  FILL_3576
timestamp 1713400504
transform 1 0 576 0 1 970
box -8 -3 16 105
use FILL  FILL_3577
timestamp 1713400504
transform 1 0 544 0 1 970
box -8 -3 16 105
use FILL  FILL_3578
timestamp 1713400504
transform 1 0 536 0 1 970
box -8 -3 16 105
use FILL  FILL_3579
timestamp 1713400504
transform 1 0 528 0 1 970
box -8 -3 16 105
use FILL  FILL_3580
timestamp 1713400504
transform 1 0 520 0 1 970
box -8 -3 16 105
use FILL  FILL_3581
timestamp 1713400504
transform 1 0 512 0 1 970
box -8 -3 16 105
use FILL  FILL_3582
timestamp 1713400504
transform 1 0 472 0 1 970
box -8 -3 16 105
use FILL  FILL_3583
timestamp 1713400504
transform 1 0 464 0 1 970
box -8 -3 16 105
use FILL  FILL_3584
timestamp 1713400504
transform 1 0 456 0 1 970
box -8 -3 16 105
use FILL  FILL_3585
timestamp 1713400504
transform 1 0 448 0 1 970
box -8 -3 16 105
use FILL  FILL_3586
timestamp 1713400504
transform 1 0 440 0 1 970
box -8 -3 16 105
use FILL  FILL_3587
timestamp 1713400504
transform 1 0 432 0 1 970
box -8 -3 16 105
use FILL  FILL_3588
timestamp 1713400504
transform 1 0 408 0 1 970
box -8 -3 16 105
use FILL  FILL_3589
timestamp 1713400504
transform 1 0 400 0 1 970
box -8 -3 16 105
use FILL  FILL_3590
timestamp 1713400504
transform 1 0 392 0 1 970
box -8 -3 16 105
use FILL  FILL_3591
timestamp 1713400504
transform 1 0 384 0 1 970
box -8 -3 16 105
use FILL  FILL_3592
timestamp 1713400504
transform 1 0 344 0 1 970
box -8 -3 16 105
use FILL  FILL_3593
timestamp 1713400504
transform 1 0 336 0 1 970
box -8 -3 16 105
use FILL  FILL_3594
timestamp 1713400504
transform 1 0 328 0 1 970
box -8 -3 16 105
use FILL  FILL_3595
timestamp 1713400504
transform 1 0 320 0 1 970
box -8 -3 16 105
use FILL  FILL_3596
timestamp 1713400504
transform 1 0 312 0 1 970
box -8 -3 16 105
use FILL  FILL_3597
timestamp 1713400504
transform 1 0 304 0 1 970
box -8 -3 16 105
use FILL  FILL_3598
timestamp 1713400504
transform 1 0 296 0 1 970
box -8 -3 16 105
use FILL  FILL_3599
timestamp 1713400504
transform 1 0 256 0 1 970
box -8 -3 16 105
use FILL  FILL_3600
timestamp 1713400504
transform 1 0 248 0 1 970
box -8 -3 16 105
use FILL  FILL_3601
timestamp 1713400504
transform 1 0 240 0 1 970
box -8 -3 16 105
use FILL  FILL_3602
timestamp 1713400504
transform 1 0 232 0 1 970
box -8 -3 16 105
use FILL  FILL_3603
timestamp 1713400504
transform 1 0 224 0 1 970
box -8 -3 16 105
use FILL  FILL_3604
timestamp 1713400504
transform 1 0 192 0 1 970
box -8 -3 16 105
use FILL  FILL_3605
timestamp 1713400504
transform 1 0 184 0 1 970
box -8 -3 16 105
use FILL  FILL_3606
timestamp 1713400504
transform 1 0 176 0 1 970
box -8 -3 16 105
use FILL  FILL_3607
timestamp 1713400504
transform 1 0 168 0 1 970
box -8 -3 16 105
use FILL  FILL_3608
timestamp 1713400504
transform 1 0 3008 0 -1 970
box -8 -3 16 105
use FILL  FILL_3609
timestamp 1713400504
transform 1 0 2944 0 -1 970
box -8 -3 16 105
use FILL  FILL_3610
timestamp 1713400504
transform 1 0 2936 0 -1 970
box -8 -3 16 105
use FILL  FILL_3611
timestamp 1713400504
transform 1 0 2928 0 -1 970
box -8 -3 16 105
use FILL  FILL_3612
timestamp 1713400504
transform 1 0 2920 0 -1 970
box -8 -3 16 105
use FILL  FILL_3613
timestamp 1713400504
transform 1 0 2912 0 -1 970
box -8 -3 16 105
use FILL  FILL_3614
timestamp 1713400504
transform 1 0 2904 0 -1 970
box -8 -3 16 105
use FILL  FILL_3615
timestamp 1713400504
transform 1 0 2856 0 -1 970
box -8 -3 16 105
use FILL  FILL_3616
timestamp 1713400504
transform 1 0 2848 0 -1 970
box -8 -3 16 105
use FILL  FILL_3617
timestamp 1713400504
transform 1 0 2840 0 -1 970
box -8 -3 16 105
use FILL  FILL_3618
timestamp 1713400504
transform 1 0 2832 0 -1 970
box -8 -3 16 105
use FILL  FILL_3619
timestamp 1713400504
transform 1 0 2824 0 -1 970
box -8 -3 16 105
use FILL  FILL_3620
timestamp 1713400504
transform 1 0 2816 0 -1 970
box -8 -3 16 105
use FILL  FILL_3621
timestamp 1713400504
transform 1 0 2808 0 -1 970
box -8 -3 16 105
use FILL  FILL_3622
timestamp 1713400504
transform 1 0 2800 0 -1 970
box -8 -3 16 105
use FILL  FILL_3623
timestamp 1713400504
transform 1 0 2792 0 -1 970
box -8 -3 16 105
use FILL  FILL_3624
timestamp 1713400504
transform 1 0 2784 0 -1 970
box -8 -3 16 105
use FILL  FILL_3625
timestamp 1713400504
transform 1 0 2776 0 -1 970
box -8 -3 16 105
use FILL  FILL_3626
timestamp 1713400504
transform 1 0 2768 0 -1 970
box -8 -3 16 105
use FILL  FILL_3627
timestamp 1713400504
transform 1 0 2760 0 -1 970
box -8 -3 16 105
use FILL  FILL_3628
timestamp 1713400504
transform 1 0 2728 0 -1 970
box -8 -3 16 105
use FILL  FILL_3629
timestamp 1713400504
transform 1 0 2720 0 -1 970
box -8 -3 16 105
use FILL  FILL_3630
timestamp 1713400504
transform 1 0 2712 0 -1 970
box -8 -3 16 105
use FILL  FILL_3631
timestamp 1713400504
transform 1 0 2704 0 -1 970
box -8 -3 16 105
use FILL  FILL_3632
timestamp 1713400504
transform 1 0 2696 0 -1 970
box -8 -3 16 105
use FILL  FILL_3633
timestamp 1713400504
transform 1 0 2688 0 -1 970
box -8 -3 16 105
use FILL  FILL_3634
timestamp 1713400504
transform 1 0 2680 0 -1 970
box -8 -3 16 105
use FILL  FILL_3635
timestamp 1713400504
transform 1 0 2672 0 -1 970
box -8 -3 16 105
use FILL  FILL_3636
timestamp 1713400504
transform 1 0 2664 0 -1 970
box -8 -3 16 105
use FILL  FILL_3637
timestamp 1713400504
transform 1 0 2656 0 -1 970
box -8 -3 16 105
use FILL  FILL_3638
timestamp 1713400504
transform 1 0 2648 0 -1 970
box -8 -3 16 105
use FILL  FILL_3639
timestamp 1713400504
transform 1 0 2640 0 -1 970
box -8 -3 16 105
use FILL  FILL_3640
timestamp 1713400504
transform 1 0 2608 0 -1 970
box -8 -3 16 105
use FILL  FILL_3641
timestamp 1713400504
transform 1 0 2600 0 -1 970
box -8 -3 16 105
use FILL  FILL_3642
timestamp 1713400504
transform 1 0 2592 0 -1 970
box -8 -3 16 105
use FILL  FILL_3643
timestamp 1713400504
transform 1 0 2584 0 -1 970
box -8 -3 16 105
use FILL  FILL_3644
timestamp 1713400504
transform 1 0 2480 0 -1 970
box -8 -3 16 105
use FILL  FILL_3645
timestamp 1713400504
transform 1 0 2472 0 -1 970
box -8 -3 16 105
use FILL  FILL_3646
timestamp 1713400504
transform 1 0 2464 0 -1 970
box -8 -3 16 105
use FILL  FILL_3647
timestamp 1713400504
transform 1 0 2432 0 -1 970
box -8 -3 16 105
use FILL  FILL_3648
timestamp 1713400504
transform 1 0 2424 0 -1 970
box -8 -3 16 105
use FILL  FILL_3649
timestamp 1713400504
transform 1 0 2416 0 -1 970
box -8 -3 16 105
use FILL  FILL_3650
timestamp 1713400504
transform 1 0 2408 0 -1 970
box -8 -3 16 105
use FILL  FILL_3651
timestamp 1713400504
transform 1 0 2344 0 -1 970
box -8 -3 16 105
use FILL  FILL_3652
timestamp 1713400504
transform 1 0 2336 0 -1 970
box -8 -3 16 105
use FILL  FILL_3653
timestamp 1713400504
transform 1 0 2328 0 -1 970
box -8 -3 16 105
use FILL  FILL_3654
timestamp 1713400504
transform 1 0 2320 0 -1 970
box -8 -3 16 105
use FILL  FILL_3655
timestamp 1713400504
transform 1 0 2312 0 -1 970
box -8 -3 16 105
use FILL  FILL_3656
timestamp 1713400504
transform 1 0 2264 0 -1 970
box -8 -3 16 105
use FILL  FILL_3657
timestamp 1713400504
transform 1 0 2256 0 -1 970
box -8 -3 16 105
use FILL  FILL_3658
timestamp 1713400504
transform 1 0 2248 0 -1 970
box -8 -3 16 105
use FILL  FILL_3659
timestamp 1713400504
transform 1 0 2240 0 -1 970
box -8 -3 16 105
use FILL  FILL_3660
timestamp 1713400504
transform 1 0 2232 0 -1 970
box -8 -3 16 105
use FILL  FILL_3661
timestamp 1713400504
transform 1 0 2168 0 -1 970
box -8 -3 16 105
use FILL  FILL_3662
timestamp 1713400504
transform 1 0 2160 0 -1 970
box -8 -3 16 105
use FILL  FILL_3663
timestamp 1713400504
transform 1 0 2152 0 -1 970
box -8 -3 16 105
use FILL  FILL_3664
timestamp 1713400504
transform 1 0 2144 0 -1 970
box -8 -3 16 105
use FILL  FILL_3665
timestamp 1713400504
transform 1 0 2136 0 -1 970
box -8 -3 16 105
use FILL  FILL_3666
timestamp 1713400504
transform 1 0 2088 0 -1 970
box -8 -3 16 105
use FILL  FILL_3667
timestamp 1713400504
transform 1 0 2080 0 -1 970
box -8 -3 16 105
use FILL  FILL_3668
timestamp 1713400504
transform 1 0 2072 0 -1 970
box -8 -3 16 105
use FILL  FILL_3669
timestamp 1713400504
transform 1 0 2064 0 -1 970
box -8 -3 16 105
use FILL  FILL_3670
timestamp 1713400504
transform 1 0 2056 0 -1 970
box -8 -3 16 105
use FILL  FILL_3671
timestamp 1713400504
transform 1 0 2048 0 -1 970
box -8 -3 16 105
use FILL  FILL_3672
timestamp 1713400504
transform 1 0 2040 0 -1 970
box -8 -3 16 105
use FILL  FILL_3673
timestamp 1713400504
transform 1 0 2016 0 -1 970
box -8 -3 16 105
use FILL  FILL_3674
timestamp 1713400504
transform 1 0 1952 0 -1 970
box -8 -3 16 105
use FILL  FILL_3675
timestamp 1713400504
transform 1 0 1944 0 -1 970
box -8 -3 16 105
use FILL  FILL_3676
timestamp 1713400504
transform 1 0 1936 0 -1 970
box -8 -3 16 105
use FILL  FILL_3677
timestamp 1713400504
transform 1 0 1928 0 -1 970
box -8 -3 16 105
use FILL  FILL_3678
timestamp 1713400504
transform 1 0 1888 0 -1 970
box -8 -3 16 105
use FILL  FILL_3679
timestamp 1713400504
transform 1 0 1880 0 -1 970
box -8 -3 16 105
use FILL  FILL_3680
timestamp 1713400504
transform 1 0 1872 0 -1 970
box -8 -3 16 105
use FILL  FILL_3681
timestamp 1713400504
transform 1 0 1864 0 -1 970
box -8 -3 16 105
use FILL  FILL_3682
timestamp 1713400504
transform 1 0 1856 0 -1 970
box -8 -3 16 105
use FILL  FILL_3683
timestamp 1713400504
transform 1 0 1816 0 -1 970
box -8 -3 16 105
use FILL  FILL_3684
timestamp 1713400504
transform 1 0 1808 0 -1 970
box -8 -3 16 105
use FILL  FILL_3685
timestamp 1713400504
transform 1 0 1800 0 -1 970
box -8 -3 16 105
use FILL  FILL_3686
timestamp 1713400504
transform 1 0 1792 0 -1 970
box -8 -3 16 105
use FILL  FILL_3687
timestamp 1713400504
transform 1 0 1784 0 -1 970
box -8 -3 16 105
use FILL  FILL_3688
timestamp 1713400504
transform 1 0 1744 0 -1 970
box -8 -3 16 105
use FILL  FILL_3689
timestamp 1713400504
transform 1 0 1736 0 -1 970
box -8 -3 16 105
use FILL  FILL_3690
timestamp 1713400504
transform 1 0 1728 0 -1 970
box -8 -3 16 105
use FILL  FILL_3691
timestamp 1713400504
transform 1 0 1720 0 -1 970
box -8 -3 16 105
use FILL  FILL_3692
timestamp 1713400504
transform 1 0 1712 0 -1 970
box -8 -3 16 105
use FILL  FILL_3693
timestamp 1713400504
transform 1 0 1704 0 -1 970
box -8 -3 16 105
use FILL  FILL_3694
timestamp 1713400504
transform 1 0 1656 0 -1 970
box -8 -3 16 105
use FILL  FILL_3695
timestamp 1713400504
transform 1 0 1648 0 -1 970
box -8 -3 16 105
use FILL  FILL_3696
timestamp 1713400504
transform 1 0 1640 0 -1 970
box -8 -3 16 105
use FILL  FILL_3697
timestamp 1713400504
transform 1 0 1632 0 -1 970
box -8 -3 16 105
use FILL  FILL_3698
timestamp 1713400504
transform 1 0 1624 0 -1 970
box -8 -3 16 105
use FILL  FILL_3699
timestamp 1713400504
transform 1 0 1616 0 -1 970
box -8 -3 16 105
use FILL  FILL_3700
timestamp 1713400504
transform 1 0 1608 0 -1 970
box -8 -3 16 105
use FILL  FILL_3701
timestamp 1713400504
transform 1 0 1600 0 -1 970
box -8 -3 16 105
use FILL  FILL_3702
timestamp 1713400504
transform 1 0 1552 0 -1 970
box -8 -3 16 105
use FILL  FILL_3703
timestamp 1713400504
transform 1 0 1544 0 -1 970
box -8 -3 16 105
use FILL  FILL_3704
timestamp 1713400504
transform 1 0 1536 0 -1 970
box -8 -3 16 105
use FILL  FILL_3705
timestamp 1713400504
transform 1 0 1528 0 -1 970
box -8 -3 16 105
use FILL  FILL_3706
timestamp 1713400504
transform 1 0 1520 0 -1 970
box -8 -3 16 105
use FILL  FILL_3707
timestamp 1713400504
transform 1 0 1512 0 -1 970
box -8 -3 16 105
use FILL  FILL_3708
timestamp 1713400504
transform 1 0 1480 0 -1 970
box -8 -3 16 105
use FILL  FILL_3709
timestamp 1713400504
transform 1 0 1472 0 -1 970
box -8 -3 16 105
use FILL  FILL_3710
timestamp 1713400504
transform 1 0 1464 0 -1 970
box -8 -3 16 105
use FILL  FILL_3711
timestamp 1713400504
transform 1 0 1456 0 -1 970
box -8 -3 16 105
use FILL  FILL_3712
timestamp 1713400504
transform 1 0 1448 0 -1 970
box -8 -3 16 105
use FILL  FILL_3713
timestamp 1713400504
transform 1 0 1440 0 -1 970
box -8 -3 16 105
use FILL  FILL_3714
timestamp 1713400504
transform 1 0 1392 0 -1 970
box -8 -3 16 105
use FILL  FILL_3715
timestamp 1713400504
transform 1 0 1384 0 -1 970
box -8 -3 16 105
use FILL  FILL_3716
timestamp 1713400504
transform 1 0 1376 0 -1 970
box -8 -3 16 105
use FILL  FILL_3717
timestamp 1713400504
transform 1 0 1368 0 -1 970
box -8 -3 16 105
use FILL  FILL_3718
timestamp 1713400504
transform 1 0 1360 0 -1 970
box -8 -3 16 105
use FILL  FILL_3719
timestamp 1713400504
transform 1 0 1352 0 -1 970
box -8 -3 16 105
use FILL  FILL_3720
timestamp 1713400504
transform 1 0 1344 0 -1 970
box -8 -3 16 105
use FILL  FILL_3721
timestamp 1713400504
transform 1 0 1336 0 -1 970
box -8 -3 16 105
use FILL  FILL_3722
timestamp 1713400504
transform 1 0 1288 0 -1 970
box -8 -3 16 105
use FILL  FILL_3723
timestamp 1713400504
transform 1 0 1280 0 -1 970
box -8 -3 16 105
use FILL  FILL_3724
timestamp 1713400504
transform 1 0 1272 0 -1 970
box -8 -3 16 105
use FILL  FILL_3725
timestamp 1713400504
transform 1 0 1264 0 -1 970
box -8 -3 16 105
use FILL  FILL_3726
timestamp 1713400504
transform 1 0 1256 0 -1 970
box -8 -3 16 105
use FILL  FILL_3727
timestamp 1713400504
transform 1 0 1248 0 -1 970
box -8 -3 16 105
use FILL  FILL_3728
timestamp 1713400504
transform 1 0 1240 0 -1 970
box -8 -3 16 105
use FILL  FILL_3729
timestamp 1713400504
transform 1 0 1232 0 -1 970
box -8 -3 16 105
use FILL  FILL_3730
timestamp 1713400504
transform 1 0 1224 0 -1 970
box -8 -3 16 105
use FILL  FILL_3731
timestamp 1713400504
transform 1 0 1176 0 -1 970
box -8 -3 16 105
use FILL  FILL_3732
timestamp 1713400504
transform 1 0 1168 0 -1 970
box -8 -3 16 105
use FILL  FILL_3733
timestamp 1713400504
transform 1 0 1160 0 -1 970
box -8 -3 16 105
use FILL  FILL_3734
timestamp 1713400504
transform 1 0 1152 0 -1 970
box -8 -3 16 105
use FILL  FILL_3735
timestamp 1713400504
transform 1 0 1144 0 -1 970
box -8 -3 16 105
use FILL  FILL_3736
timestamp 1713400504
transform 1 0 1136 0 -1 970
box -8 -3 16 105
use FILL  FILL_3737
timestamp 1713400504
transform 1 0 1128 0 -1 970
box -8 -3 16 105
use FILL  FILL_3738
timestamp 1713400504
transform 1 0 1120 0 -1 970
box -8 -3 16 105
use FILL  FILL_3739
timestamp 1713400504
transform 1 0 1072 0 -1 970
box -8 -3 16 105
use FILL  FILL_3740
timestamp 1713400504
transform 1 0 1064 0 -1 970
box -8 -3 16 105
use FILL  FILL_3741
timestamp 1713400504
transform 1 0 1056 0 -1 970
box -8 -3 16 105
use FILL  FILL_3742
timestamp 1713400504
transform 1 0 1048 0 -1 970
box -8 -3 16 105
use FILL  FILL_3743
timestamp 1713400504
transform 1 0 1040 0 -1 970
box -8 -3 16 105
use FILL  FILL_3744
timestamp 1713400504
transform 1 0 1032 0 -1 970
box -8 -3 16 105
use FILL  FILL_3745
timestamp 1713400504
transform 1 0 1024 0 -1 970
box -8 -3 16 105
use FILL  FILL_3746
timestamp 1713400504
transform 1 0 1016 0 -1 970
box -8 -3 16 105
use FILL  FILL_3747
timestamp 1713400504
transform 1 0 1008 0 -1 970
box -8 -3 16 105
use FILL  FILL_3748
timestamp 1713400504
transform 1 0 960 0 -1 970
box -8 -3 16 105
use FILL  FILL_3749
timestamp 1713400504
transform 1 0 952 0 -1 970
box -8 -3 16 105
use FILL  FILL_3750
timestamp 1713400504
transform 1 0 944 0 -1 970
box -8 -3 16 105
use FILL  FILL_3751
timestamp 1713400504
transform 1 0 936 0 -1 970
box -8 -3 16 105
use FILL  FILL_3752
timestamp 1713400504
transform 1 0 928 0 -1 970
box -8 -3 16 105
use FILL  FILL_3753
timestamp 1713400504
transform 1 0 920 0 -1 970
box -8 -3 16 105
use FILL  FILL_3754
timestamp 1713400504
transform 1 0 912 0 -1 970
box -8 -3 16 105
use FILL  FILL_3755
timestamp 1713400504
transform 1 0 904 0 -1 970
box -8 -3 16 105
use FILL  FILL_3756
timestamp 1713400504
transform 1 0 896 0 -1 970
box -8 -3 16 105
use FILL  FILL_3757
timestamp 1713400504
transform 1 0 848 0 -1 970
box -8 -3 16 105
use FILL  FILL_3758
timestamp 1713400504
transform 1 0 840 0 -1 970
box -8 -3 16 105
use FILL  FILL_3759
timestamp 1713400504
transform 1 0 832 0 -1 970
box -8 -3 16 105
use FILL  FILL_3760
timestamp 1713400504
transform 1 0 824 0 -1 970
box -8 -3 16 105
use FILL  FILL_3761
timestamp 1713400504
transform 1 0 816 0 -1 970
box -8 -3 16 105
use FILL  FILL_3762
timestamp 1713400504
transform 1 0 808 0 -1 970
box -8 -3 16 105
use FILL  FILL_3763
timestamp 1713400504
transform 1 0 800 0 -1 970
box -8 -3 16 105
use FILL  FILL_3764
timestamp 1713400504
transform 1 0 696 0 -1 970
box -8 -3 16 105
use FILL  FILL_3765
timestamp 1713400504
transform 1 0 688 0 -1 970
box -8 -3 16 105
use FILL  FILL_3766
timestamp 1713400504
transform 1 0 680 0 -1 970
box -8 -3 16 105
use FILL  FILL_3767
timestamp 1713400504
transform 1 0 672 0 -1 970
box -8 -3 16 105
use FILL  FILL_3768
timestamp 1713400504
transform 1 0 632 0 -1 970
box -8 -3 16 105
use FILL  FILL_3769
timestamp 1713400504
transform 1 0 624 0 -1 970
box -8 -3 16 105
use FILL  FILL_3770
timestamp 1713400504
transform 1 0 616 0 -1 970
box -8 -3 16 105
use FILL  FILL_3771
timestamp 1713400504
transform 1 0 608 0 -1 970
box -8 -3 16 105
use FILL  FILL_3772
timestamp 1713400504
transform 1 0 576 0 -1 970
box -8 -3 16 105
use FILL  FILL_3773
timestamp 1713400504
transform 1 0 568 0 -1 970
box -8 -3 16 105
use FILL  FILL_3774
timestamp 1713400504
transform 1 0 560 0 -1 970
box -8 -3 16 105
use FILL  FILL_3775
timestamp 1713400504
transform 1 0 552 0 -1 970
box -8 -3 16 105
use FILL  FILL_3776
timestamp 1713400504
transform 1 0 448 0 -1 970
box -8 -3 16 105
use FILL  FILL_3777
timestamp 1713400504
transform 1 0 440 0 -1 970
box -8 -3 16 105
use FILL  FILL_3778
timestamp 1713400504
transform 1 0 432 0 -1 970
box -8 -3 16 105
use FILL  FILL_3779
timestamp 1713400504
transform 1 0 424 0 -1 970
box -8 -3 16 105
use FILL  FILL_3780
timestamp 1713400504
transform 1 0 416 0 -1 970
box -8 -3 16 105
use FILL  FILL_3781
timestamp 1713400504
transform 1 0 368 0 -1 970
box -8 -3 16 105
use FILL  FILL_3782
timestamp 1713400504
transform 1 0 360 0 -1 970
box -8 -3 16 105
use FILL  FILL_3783
timestamp 1713400504
transform 1 0 352 0 -1 970
box -8 -3 16 105
use FILL  FILL_3784
timestamp 1713400504
transform 1 0 344 0 -1 970
box -8 -3 16 105
use FILL  FILL_3785
timestamp 1713400504
transform 1 0 336 0 -1 970
box -8 -3 16 105
use FILL  FILL_3786
timestamp 1713400504
transform 1 0 232 0 -1 970
box -8 -3 16 105
use FILL  FILL_3787
timestamp 1713400504
transform 1 0 224 0 -1 970
box -8 -3 16 105
use FILL  FILL_3788
timestamp 1713400504
transform 1 0 216 0 -1 970
box -8 -3 16 105
use FILL  FILL_3789
timestamp 1713400504
transform 1 0 208 0 -1 970
box -8 -3 16 105
use FILL  FILL_3790
timestamp 1713400504
transform 1 0 176 0 -1 970
box -8 -3 16 105
use FILL  FILL_3791
timestamp 1713400504
transform 1 0 168 0 -1 970
box -8 -3 16 105
use FILL  FILL_3792
timestamp 1713400504
transform 1 0 160 0 -1 970
box -8 -3 16 105
use FILL  FILL_3793
timestamp 1713400504
transform 1 0 152 0 -1 970
box -8 -3 16 105
use FILL  FILL_3794
timestamp 1713400504
transform 1 0 144 0 -1 970
box -8 -3 16 105
use FILL  FILL_3795
timestamp 1713400504
transform 1 0 104 0 -1 970
box -8 -3 16 105
use FILL  FILL_3796
timestamp 1713400504
transform 1 0 96 0 -1 970
box -8 -3 16 105
use FILL  FILL_3797
timestamp 1713400504
transform 1 0 88 0 -1 970
box -8 -3 16 105
use FILL  FILL_3798
timestamp 1713400504
transform 1 0 80 0 -1 970
box -8 -3 16 105
use FILL  FILL_3799
timestamp 1713400504
transform 1 0 72 0 -1 970
box -8 -3 16 105
use FILL  FILL_3800
timestamp 1713400504
transform 1 0 3008 0 1 770
box -8 -3 16 105
use FILL  FILL_3801
timestamp 1713400504
transform 1 0 2920 0 1 770
box -8 -3 16 105
use FILL  FILL_3802
timestamp 1713400504
transform 1 0 2912 0 1 770
box -8 -3 16 105
use FILL  FILL_3803
timestamp 1713400504
transform 1 0 2904 0 1 770
box -8 -3 16 105
use FILL  FILL_3804
timestamp 1713400504
transform 1 0 2856 0 1 770
box -8 -3 16 105
use FILL  FILL_3805
timestamp 1713400504
transform 1 0 2848 0 1 770
box -8 -3 16 105
use FILL  FILL_3806
timestamp 1713400504
transform 1 0 2840 0 1 770
box -8 -3 16 105
use FILL  FILL_3807
timestamp 1713400504
transform 1 0 2752 0 1 770
box -8 -3 16 105
use FILL  FILL_3808
timestamp 1713400504
transform 1 0 2744 0 1 770
box -8 -3 16 105
use FILL  FILL_3809
timestamp 1713400504
transform 1 0 2736 0 1 770
box -8 -3 16 105
use FILL  FILL_3810
timestamp 1713400504
transform 1 0 2728 0 1 770
box -8 -3 16 105
use FILL  FILL_3811
timestamp 1713400504
transform 1 0 2680 0 1 770
box -8 -3 16 105
use FILL  FILL_3812
timestamp 1713400504
transform 1 0 2672 0 1 770
box -8 -3 16 105
use FILL  FILL_3813
timestamp 1713400504
transform 1 0 2648 0 1 770
box -8 -3 16 105
use FILL  FILL_3814
timestamp 1713400504
transform 1 0 2640 0 1 770
box -8 -3 16 105
use FILL  FILL_3815
timestamp 1713400504
transform 1 0 2536 0 1 770
box -8 -3 16 105
use FILL  FILL_3816
timestamp 1713400504
transform 1 0 2528 0 1 770
box -8 -3 16 105
use FILL  FILL_3817
timestamp 1713400504
transform 1 0 2520 0 1 770
box -8 -3 16 105
use FILL  FILL_3818
timestamp 1713400504
transform 1 0 2496 0 1 770
box -8 -3 16 105
use FILL  FILL_3819
timestamp 1713400504
transform 1 0 2456 0 1 770
box -8 -3 16 105
use FILL  FILL_3820
timestamp 1713400504
transform 1 0 2448 0 1 770
box -8 -3 16 105
use FILL  FILL_3821
timestamp 1713400504
transform 1 0 2440 0 1 770
box -8 -3 16 105
use FILL  FILL_3822
timestamp 1713400504
transform 1 0 2432 0 1 770
box -8 -3 16 105
use FILL  FILL_3823
timestamp 1713400504
transform 1 0 2424 0 1 770
box -8 -3 16 105
use FILL  FILL_3824
timestamp 1713400504
transform 1 0 2416 0 1 770
box -8 -3 16 105
use FILL  FILL_3825
timestamp 1713400504
transform 1 0 2408 0 1 770
box -8 -3 16 105
use FILL  FILL_3826
timestamp 1713400504
transform 1 0 2376 0 1 770
box -8 -3 16 105
use FILL  FILL_3827
timestamp 1713400504
transform 1 0 2368 0 1 770
box -8 -3 16 105
use FILL  FILL_3828
timestamp 1713400504
transform 1 0 2360 0 1 770
box -8 -3 16 105
use FILL  FILL_3829
timestamp 1713400504
transform 1 0 2352 0 1 770
box -8 -3 16 105
use FILL  FILL_3830
timestamp 1713400504
transform 1 0 2312 0 1 770
box -8 -3 16 105
use FILL  FILL_3831
timestamp 1713400504
transform 1 0 2304 0 1 770
box -8 -3 16 105
use FILL  FILL_3832
timestamp 1713400504
transform 1 0 2296 0 1 770
box -8 -3 16 105
use FILL  FILL_3833
timestamp 1713400504
transform 1 0 2288 0 1 770
box -8 -3 16 105
use FILL  FILL_3834
timestamp 1713400504
transform 1 0 2280 0 1 770
box -8 -3 16 105
use FILL  FILL_3835
timestamp 1713400504
transform 1 0 2216 0 1 770
box -8 -3 16 105
use FILL  FILL_3836
timestamp 1713400504
transform 1 0 2208 0 1 770
box -8 -3 16 105
use FILL  FILL_3837
timestamp 1713400504
transform 1 0 2184 0 1 770
box -8 -3 16 105
use FILL  FILL_3838
timestamp 1713400504
transform 1 0 2176 0 1 770
box -8 -3 16 105
use FILL  FILL_3839
timestamp 1713400504
transform 1 0 2168 0 1 770
box -8 -3 16 105
use FILL  FILL_3840
timestamp 1713400504
transform 1 0 2160 0 1 770
box -8 -3 16 105
use FILL  FILL_3841
timestamp 1713400504
transform 1 0 2152 0 1 770
box -8 -3 16 105
use FILL  FILL_3842
timestamp 1713400504
transform 1 0 2144 0 1 770
box -8 -3 16 105
use FILL  FILL_3843
timestamp 1713400504
transform 1 0 2136 0 1 770
box -8 -3 16 105
use FILL  FILL_3844
timestamp 1713400504
transform 1 0 2104 0 1 770
box -8 -3 16 105
use FILL  FILL_3845
timestamp 1713400504
transform 1 0 2096 0 1 770
box -8 -3 16 105
use FILL  FILL_3846
timestamp 1713400504
transform 1 0 2088 0 1 770
box -8 -3 16 105
use FILL  FILL_3847
timestamp 1713400504
transform 1 0 2080 0 1 770
box -8 -3 16 105
use FILL  FILL_3848
timestamp 1713400504
transform 1 0 2072 0 1 770
box -8 -3 16 105
use FILL  FILL_3849
timestamp 1713400504
transform 1 0 2064 0 1 770
box -8 -3 16 105
use FILL  FILL_3850
timestamp 1713400504
transform 1 0 2032 0 1 770
box -8 -3 16 105
use FILL  FILL_3851
timestamp 1713400504
transform 1 0 2024 0 1 770
box -8 -3 16 105
use FILL  FILL_3852
timestamp 1713400504
transform 1 0 2016 0 1 770
box -8 -3 16 105
use FILL  FILL_3853
timestamp 1713400504
transform 1 0 2008 0 1 770
box -8 -3 16 105
use FILL  FILL_3854
timestamp 1713400504
transform 1 0 2000 0 1 770
box -8 -3 16 105
use FILL  FILL_3855
timestamp 1713400504
transform 1 0 1992 0 1 770
box -8 -3 16 105
use FILL  FILL_3856
timestamp 1713400504
transform 1 0 1984 0 1 770
box -8 -3 16 105
use FILL  FILL_3857
timestamp 1713400504
transform 1 0 1976 0 1 770
box -8 -3 16 105
use FILL  FILL_3858
timestamp 1713400504
transform 1 0 1968 0 1 770
box -8 -3 16 105
use FILL  FILL_3859
timestamp 1713400504
transform 1 0 1928 0 1 770
box -8 -3 16 105
use FILL  FILL_3860
timestamp 1713400504
transform 1 0 1920 0 1 770
box -8 -3 16 105
use FILL  FILL_3861
timestamp 1713400504
transform 1 0 1912 0 1 770
box -8 -3 16 105
use FILL  FILL_3862
timestamp 1713400504
transform 1 0 1904 0 1 770
box -8 -3 16 105
use FILL  FILL_3863
timestamp 1713400504
transform 1 0 1896 0 1 770
box -8 -3 16 105
use FILL  FILL_3864
timestamp 1713400504
transform 1 0 1888 0 1 770
box -8 -3 16 105
use FILL  FILL_3865
timestamp 1713400504
transform 1 0 1880 0 1 770
box -8 -3 16 105
use FILL  FILL_3866
timestamp 1713400504
transform 1 0 1856 0 1 770
box -8 -3 16 105
use FILL  FILL_3867
timestamp 1713400504
transform 1 0 1848 0 1 770
box -8 -3 16 105
use FILL  FILL_3868
timestamp 1713400504
transform 1 0 1840 0 1 770
box -8 -3 16 105
use FILL  FILL_3869
timestamp 1713400504
transform 1 0 1832 0 1 770
box -8 -3 16 105
use FILL  FILL_3870
timestamp 1713400504
transform 1 0 1824 0 1 770
box -8 -3 16 105
use FILL  FILL_3871
timestamp 1713400504
transform 1 0 1816 0 1 770
box -8 -3 16 105
use FILL  FILL_3872
timestamp 1713400504
transform 1 0 1808 0 1 770
box -8 -3 16 105
use FILL  FILL_3873
timestamp 1713400504
transform 1 0 1800 0 1 770
box -8 -3 16 105
use FILL  FILL_3874
timestamp 1713400504
transform 1 0 1768 0 1 770
box -8 -3 16 105
use FILL  FILL_3875
timestamp 1713400504
transform 1 0 1760 0 1 770
box -8 -3 16 105
use FILL  FILL_3876
timestamp 1713400504
transform 1 0 1752 0 1 770
box -8 -3 16 105
use FILL  FILL_3877
timestamp 1713400504
transform 1 0 1744 0 1 770
box -8 -3 16 105
use FILL  FILL_3878
timestamp 1713400504
transform 1 0 1736 0 1 770
box -8 -3 16 105
use FILL  FILL_3879
timestamp 1713400504
transform 1 0 1728 0 1 770
box -8 -3 16 105
use FILL  FILL_3880
timestamp 1713400504
transform 1 0 1720 0 1 770
box -8 -3 16 105
use FILL  FILL_3881
timestamp 1713400504
transform 1 0 1712 0 1 770
box -8 -3 16 105
use FILL  FILL_3882
timestamp 1713400504
transform 1 0 1680 0 1 770
box -8 -3 16 105
use FILL  FILL_3883
timestamp 1713400504
transform 1 0 1672 0 1 770
box -8 -3 16 105
use FILL  FILL_3884
timestamp 1713400504
transform 1 0 1664 0 1 770
box -8 -3 16 105
use FILL  FILL_3885
timestamp 1713400504
transform 1 0 1656 0 1 770
box -8 -3 16 105
use FILL  FILL_3886
timestamp 1713400504
transform 1 0 1648 0 1 770
box -8 -3 16 105
use FILL  FILL_3887
timestamp 1713400504
transform 1 0 1640 0 1 770
box -8 -3 16 105
use FILL  FILL_3888
timestamp 1713400504
transform 1 0 1632 0 1 770
box -8 -3 16 105
use FILL  FILL_3889
timestamp 1713400504
transform 1 0 1624 0 1 770
box -8 -3 16 105
use FILL  FILL_3890
timestamp 1713400504
transform 1 0 1592 0 1 770
box -8 -3 16 105
use FILL  FILL_3891
timestamp 1713400504
transform 1 0 1584 0 1 770
box -8 -3 16 105
use FILL  FILL_3892
timestamp 1713400504
transform 1 0 1576 0 1 770
box -8 -3 16 105
use FILL  FILL_3893
timestamp 1713400504
transform 1 0 1568 0 1 770
box -8 -3 16 105
use FILL  FILL_3894
timestamp 1713400504
transform 1 0 1560 0 1 770
box -8 -3 16 105
use FILL  FILL_3895
timestamp 1713400504
transform 1 0 1552 0 1 770
box -8 -3 16 105
use FILL  FILL_3896
timestamp 1713400504
transform 1 0 1544 0 1 770
box -8 -3 16 105
use FILL  FILL_3897
timestamp 1713400504
transform 1 0 1536 0 1 770
box -8 -3 16 105
use FILL  FILL_3898
timestamp 1713400504
transform 1 0 1528 0 1 770
box -8 -3 16 105
use FILL  FILL_3899
timestamp 1713400504
transform 1 0 1480 0 1 770
box -8 -3 16 105
use FILL  FILL_3900
timestamp 1713400504
transform 1 0 1472 0 1 770
box -8 -3 16 105
use FILL  FILL_3901
timestamp 1713400504
transform 1 0 1464 0 1 770
box -8 -3 16 105
use FILL  FILL_3902
timestamp 1713400504
transform 1 0 1456 0 1 770
box -8 -3 16 105
use FILL  FILL_3903
timestamp 1713400504
transform 1 0 1448 0 1 770
box -8 -3 16 105
use FILL  FILL_3904
timestamp 1713400504
transform 1 0 1440 0 1 770
box -8 -3 16 105
use FILL  FILL_3905
timestamp 1713400504
transform 1 0 1432 0 1 770
box -8 -3 16 105
use FILL  FILL_3906
timestamp 1713400504
transform 1 0 1424 0 1 770
box -8 -3 16 105
use FILL  FILL_3907
timestamp 1713400504
transform 1 0 1376 0 1 770
box -8 -3 16 105
use FILL  FILL_3908
timestamp 1713400504
transform 1 0 1368 0 1 770
box -8 -3 16 105
use FILL  FILL_3909
timestamp 1713400504
transform 1 0 1360 0 1 770
box -8 -3 16 105
use FILL  FILL_3910
timestamp 1713400504
transform 1 0 1352 0 1 770
box -8 -3 16 105
use FILL  FILL_3911
timestamp 1713400504
transform 1 0 1344 0 1 770
box -8 -3 16 105
use FILL  FILL_3912
timestamp 1713400504
transform 1 0 1336 0 1 770
box -8 -3 16 105
use FILL  FILL_3913
timestamp 1713400504
transform 1 0 1328 0 1 770
box -8 -3 16 105
use FILL  FILL_3914
timestamp 1713400504
transform 1 0 1320 0 1 770
box -8 -3 16 105
use FILL  FILL_3915
timestamp 1713400504
transform 1 0 1312 0 1 770
box -8 -3 16 105
use FILL  FILL_3916
timestamp 1713400504
transform 1 0 1264 0 1 770
box -8 -3 16 105
use FILL  FILL_3917
timestamp 1713400504
transform 1 0 1256 0 1 770
box -8 -3 16 105
use FILL  FILL_3918
timestamp 1713400504
transform 1 0 1248 0 1 770
box -8 -3 16 105
use FILL  FILL_3919
timestamp 1713400504
transform 1 0 1240 0 1 770
box -8 -3 16 105
use FILL  FILL_3920
timestamp 1713400504
transform 1 0 1232 0 1 770
box -8 -3 16 105
use FILL  FILL_3921
timestamp 1713400504
transform 1 0 1224 0 1 770
box -8 -3 16 105
use FILL  FILL_3922
timestamp 1713400504
transform 1 0 1216 0 1 770
box -8 -3 16 105
use FILL  FILL_3923
timestamp 1713400504
transform 1 0 1184 0 1 770
box -8 -3 16 105
use FILL  FILL_3924
timestamp 1713400504
transform 1 0 1176 0 1 770
box -8 -3 16 105
use FILL  FILL_3925
timestamp 1713400504
transform 1 0 1168 0 1 770
box -8 -3 16 105
use FILL  FILL_3926
timestamp 1713400504
transform 1 0 1160 0 1 770
box -8 -3 16 105
use FILL  FILL_3927
timestamp 1713400504
transform 1 0 1152 0 1 770
box -8 -3 16 105
use FILL  FILL_3928
timestamp 1713400504
transform 1 0 1144 0 1 770
box -8 -3 16 105
use FILL  FILL_3929
timestamp 1713400504
transform 1 0 1136 0 1 770
box -8 -3 16 105
use FILL  FILL_3930
timestamp 1713400504
transform 1 0 1104 0 1 770
box -8 -3 16 105
use FILL  FILL_3931
timestamp 1713400504
transform 1 0 1096 0 1 770
box -8 -3 16 105
use FILL  FILL_3932
timestamp 1713400504
transform 1 0 1088 0 1 770
box -8 -3 16 105
use FILL  FILL_3933
timestamp 1713400504
transform 1 0 1080 0 1 770
box -8 -3 16 105
use FILL  FILL_3934
timestamp 1713400504
transform 1 0 1072 0 1 770
box -8 -3 16 105
use FILL  FILL_3935
timestamp 1713400504
transform 1 0 1064 0 1 770
box -8 -3 16 105
use FILL  FILL_3936
timestamp 1713400504
transform 1 0 1056 0 1 770
box -8 -3 16 105
use FILL  FILL_3937
timestamp 1713400504
transform 1 0 1024 0 1 770
box -8 -3 16 105
use FILL  FILL_3938
timestamp 1713400504
transform 1 0 1016 0 1 770
box -8 -3 16 105
use FILL  FILL_3939
timestamp 1713400504
transform 1 0 1008 0 1 770
box -8 -3 16 105
use FILL  FILL_3940
timestamp 1713400504
transform 1 0 1000 0 1 770
box -8 -3 16 105
use FILL  FILL_3941
timestamp 1713400504
transform 1 0 992 0 1 770
box -8 -3 16 105
use FILL  FILL_3942
timestamp 1713400504
transform 1 0 984 0 1 770
box -8 -3 16 105
use FILL  FILL_3943
timestamp 1713400504
transform 1 0 976 0 1 770
box -8 -3 16 105
use FILL  FILL_3944
timestamp 1713400504
transform 1 0 872 0 1 770
box -8 -3 16 105
use FILL  FILL_3945
timestamp 1713400504
transform 1 0 864 0 1 770
box -8 -3 16 105
use FILL  FILL_3946
timestamp 1713400504
transform 1 0 856 0 1 770
box -8 -3 16 105
use FILL  FILL_3947
timestamp 1713400504
transform 1 0 848 0 1 770
box -8 -3 16 105
use FILL  FILL_3948
timestamp 1713400504
transform 1 0 808 0 1 770
box -8 -3 16 105
use FILL  FILL_3949
timestamp 1713400504
transform 1 0 800 0 1 770
box -8 -3 16 105
use FILL  FILL_3950
timestamp 1713400504
transform 1 0 792 0 1 770
box -8 -3 16 105
use FILL  FILL_3951
timestamp 1713400504
transform 1 0 784 0 1 770
box -8 -3 16 105
use FILL  FILL_3952
timestamp 1713400504
transform 1 0 776 0 1 770
box -8 -3 16 105
use FILL  FILL_3953
timestamp 1713400504
transform 1 0 768 0 1 770
box -8 -3 16 105
use FILL  FILL_3954
timestamp 1713400504
transform 1 0 760 0 1 770
box -8 -3 16 105
use FILL  FILL_3955
timestamp 1713400504
transform 1 0 728 0 1 770
box -8 -3 16 105
use FILL  FILL_3956
timestamp 1713400504
transform 1 0 720 0 1 770
box -8 -3 16 105
use FILL  FILL_3957
timestamp 1713400504
transform 1 0 712 0 1 770
box -8 -3 16 105
use FILL  FILL_3958
timestamp 1713400504
transform 1 0 704 0 1 770
box -8 -3 16 105
use FILL  FILL_3959
timestamp 1713400504
transform 1 0 680 0 1 770
box -8 -3 16 105
use FILL  FILL_3960
timestamp 1713400504
transform 1 0 672 0 1 770
box -8 -3 16 105
use FILL  FILL_3961
timestamp 1713400504
transform 1 0 664 0 1 770
box -8 -3 16 105
use FILL  FILL_3962
timestamp 1713400504
transform 1 0 656 0 1 770
box -8 -3 16 105
use FILL  FILL_3963
timestamp 1713400504
transform 1 0 632 0 1 770
box -8 -3 16 105
use FILL  FILL_3964
timestamp 1713400504
transform 1 0 624 0 1 770
box -8 -3 16 105
use FILL  FILL_3965
timestamp 1713400504
transform 1 0 592 0 1 770
box -8 -3 16 105
use FILL  FILL_3966
timestamp 1713400504
transform 1 0 584 0 1 770
box -8 -3 16 105
use FILL  FILL_3967
timestamp 1713400504
transform 1 0 576 0 1 770
box -8 -3 16 105
use FILL  FILL_3968
timestamp 1713400504
transform 1 0 568 0 1 770
box -8 -3 16 105
use FILL  FILL_3969
timestamp 1713400504
transform 1 0 536 0 1 770
box -8 -3 16 105
use FILL  FILL_3970
timestamp 1713400504
transform 1 0 528 0 1 770
box -8 -3 16 105
use FILL  FILL_3971
timestamp 1713400504
transform 1 0 520 0 1 770
box -8 -3 16 105
use FILL  FILL_3972
timestamp 1713400504
transform 1 0 488 0 1 770
box -8 -3 16 105
use FILL  FILL_3973
timestamp 1713400504
transform 1 0 480 0 1 770
box -8 -3 16 105
use FILL  FILL_3974
timestamp 1713400504
transform 1 0 472 0 1 770
box -8 -3 16 105
use FILL  FILL_3975
timestamp 1713400504
transform 1 0 440 0 1 770
box -8 -3 16 105
use FILL  FILL_3976
timestamp 1713400504
transform 1 0 432 0 1 770
box -8 -3 16 105
use FILL  FILL_3977
timestamp 1713400504
transform 1 0 424 0 1 770
box -8 -3 16 105
use FILL  FILL_3978
timestamp 1713400504
transform 1 0 392 0 1 770
box -8 -3 16 105
use FILL  FILL_3979
timestamp 1713400504
transform 1 0 384 0 1 770
box -8 -3 16 105
use FILL  FILL_3980
timestamp 1713400504
transform 1 0 376 0 1 770
box -8 -3 16 105
use FILL  FILL_3981
timestamp 1713400504
transform 1 0 368 0 1 770
box -8 -3 16 105
use FILL  FILL_3982
timestamp 1713400504
transform 1 0 336 0 1 770
box -8 -3 16 105
use FILL  FILL_3983
timestamp 1713400504
transform 1 0 328 0 1 770
box -8 -3 16 105
use FILL  FILL_3984
timestamp 1713400504
transform 1 0 304 0 1 770
box -8 -3 16 105
use FILL  FILL_3985
timestamp 1713400504
transform 1 0 296 0 1 770
box -8 -3 16 105
use FILL  FILL_3986
timestamp 1713400504
transform 1 0 288 0 1 770
box -8 -3 16 105
use FILL  FILL_3987
timestamp 1713400504
transform 1 0 280 0 1 770
box -8 -3 16 105
use FILL  FILL_3988
timestamp 1713400504
transform 1 0 248 0 1 770
box -8 -3 16 105
use FILL  FILL_3989
timestamp 1713400504
transform 1 0 240 0 1 770
box -8 -3 16 105
use FILL  FILL_3990
timestamp 1713400504
transform 1 0 232 0 1 770
box -8 -3 16 105
use FILL  FILL_3991
timestamp 1713400504
transform 1 0 224 0 1 770
box -8 -3 16 105
use FILL  FILL_3992
timestamp 1713400504
transform 1 0 184 0 1 770
box -8 -3 16 105
use FILL  FILL_3993
timestamp 1713400504
transform 1 0 176 0 1 770
box -8 -3 16 105
use FILL  FILL_3994
timestamp 1713400504
transform 1 0 168 0 1 770
box -8 -3 16 105
use FILL  FILL_3995
timestamp 1713400504
transform 1 0 3008 0 -1 770
box -8 -3 16 105
use FILL  FILL_3996
timestamp 1713400504
transform 1 0 2976 0 -1 770
box -8 -3 16 105
use FILL  FILL_3997
timestamp 1713400504
transform 1 0 2968 0 -1 770
box -8 -3 16 105
use FILL  FILL_3998
timestamp 1713400504
transform 1 0 2960 0 -1 770
box -8 -3 16 105
use FILL  FILL_3999
timestamp 1713400504
transform 1 0 2952 0 -1 770
box -8 -3 16 105
use FILL  FILL_4000
timestamp 1713400504
transform 1 0 2848 0 -1 770
box -8 -3 16 105
use FILL  FILL_4001
timestamp 1713400504
transform 1 0 2840 0 -1 770
box -8 -3 16 105
use FILL  FILL_4002
timestamp 1713400504
transform 1 0 2832 0 -1 770
box -8 -3 16 105
use FILL  FILL_4003
timestamp 1713400504
transform 1 0 2808 0 -1 770
box -8 -3 16 105
use FILL  FILL_4004
timestamp 1713400504
transform 1 0 2800 0 -1 770
box -8 -3 16 105
use FILL  FILL_4005
timestamp 1713400504
transform 1 0 2792 0 -1 770
box -8 -3 16 105
use FILL  FILL_4006
timestamp 1713400504
transform 1 0 2784 0 -1 770
box -8 -3 16 105
use FILL  FILL_4007
timestamp 1713400504
transform 1 0 2776 0 -1 770
box -8 -3 16 105
use FILL  FILL_4008
timestamp 1713400504
transform 1 0 2768 0 -1 770
box -8 -3 16 105
use FILL  FILL_4009
timestamp 1713400504
transform 1 0 2760 0 -1 770
box -8 -3 16 105
use FILL  FILL_4010
timestamp 1713400504
transform 1 0 2720 0 -1 770
box -8 -3 16 105
use FILL  FILL_4011
timestamp 1713400504
transform 1 0 2712 0 -1 770
box -8 -3 16 105
use FILL  FILL_4012
timestamp 1713400504
transform 1 0 2704 0 -1 770
box -8 -3 16 105
use FILL  FILL_4013
timestamp 1713400504
transform 1 0 2696 0 -1 770
box -8 -3 16 105
use FILL  FILL_4014
timestamp 1713400504
transform 1 0 2688 0 -1 770
box -8 -3 16 105
use FILL  FILL_4015
timestamp 1713400504
transform 1 0 2680 0 -1 770
box -8 -3 16 105
use FILL  FILL_4016
timestamp 1713400504
transform 1 0 2648 0 -1 770
box -8 -3 16 105
use FILL  FILL_4017
timestamp 1713400504
transform 1 0 2640 0 -1 770
box -8 -3 16 105
use FILL  FILL_4018
timestamp 1713400504
transform 1 0 2632 0 -1 770
box -8 -3 16 105
use FILL  FILL_4019
timestamp 1713400504
transform 1 0 2624 0 -1 770
box -8 -3 16 105
use FILL  FILL_4020
timestamp 1713400504
transform 1 0 2600 0 -1 770
box -8 -3 16 105
use FILL  FILL_4021
timestamp 1713400504
transform 1 0 2592 0 -1 770
box -8 -3 16 105
use FILL  FILL_4022
timestamp 1713400504
transform 1 0 2584 0 -1 770
box -8 -3 16 105
use FILL  FILL_4023
timestamp 1713400504
transform 1 0 2576 0 -1 770
box -8 -3 16 105
use FILL  FILL_4024
timestamp 1713400504
transform 1 0 2568 0 -1 770
box -8 -3 16 105
use FILL  FILL_4025
timestamp 1713400504
transform 1 0 2560 0 -1 770
box -8 -3 16 105
use FILL  FILL_4026
timestamp 1713400504
transform 1 0 2520 0 -1 770
box -8 -3 16 105
use FILL  FILL_4027
timestamp 1713400504
transform 1 0 2512 0 -1 770
box -8 -3 16 105
use FILL  FILL_4028
timestamp 1713400504
transform 1 0 2504 0 -1 770
box -8 -3 16 105
use FILL  FILL_4029
timestamp 1713400504
transform 1 0 2496 0 -1 770
box -8 -3 16 105
use FILL  FILL_4030
timestamp 1713400504
transform 1 0 2488 0 -1 770
box -8 -3 16 105
use FILL  FILL_4031
timestamp 1713400504
transform 1 0 2464 0 -1 770
box -8 -3 16 105
use FILL  FILL_4032
timestamp 1713400504
transform 1 0 2456 0 -1 770
box -8 -3 16 105
use FILL  FILL_4033
timestamp 1713400504
transform 1 0 2424 0 -1 770
box -8 -3 16 105
use FILL  FILL_4034
timestamp 1713400504
transform 1 0 2416 0 -1 770
box -8 -3 16 105
use FILL  FILL_4035
timestamp 1713400504
transform 1 0 2408 0 -1 770
box -8 -3 16 105
use FILL  FILL_4036
timestamp 1713400504
transform 1 0 2400 0 -1 770
box -8 -3 16 105
use FILL  FILL_4037
timestamp 1713400504
transform 1 0 2392 0 -1 770
box -8 -3 16 105
use FILL  FILL_4038
timestamp 1713400504
transform 1 0 2384 0 -1 770
box -8 -3 16 105
use FILL  FILL_4039
timestamp 1713400504
transform 1 0 2376 0 -1 770
box -8 -3 16 105
use FILL  FILL_4040
timestamp 1713400504
transform 1 0 2336 0 -1 770
box -8 -3 16 105
use FILL  FILL_4041
timestamp 1713400504
transform 1 0 2328 0 -1 770
box -8 -3 16 105
use FILL  FILL_4042
timestamp 1713400504
transform 1 0 2320 0 -1 770
box -8 -3 16 105
use FILL  FILL_4043
timestamp 1713400504
transform 1 0 2312 0 -1 770
box -8 -3 16 105
use FILL  FILL_4044
timestamp 1713400504
transform 1 0 2304 0 -1 770
box -8 -3 16 105
use FILL  FILL_4045
timestamp 1713400504
transform 1 0 2272 0 -1 770
box -8 -3 16 105
use FILL  FILL_4046
timestamp 1713400504
transform 1 0 2264 0 -1 770
box -8 -3 16 105
use FILL  FILL_4047
timestamp 1713400504
transform 1 0 2256 0 -1 770
box -8 -3 16 105
use FILL  FILL_4048
timestamp 1713400504
transform 1 0 2248 0 -1 770
box -8 -3 16 105
use FILL  FILL_4049
timestamp 1713400504
transform 1 0 2240 0 -1 770
box -8 -3 16 105
use FILL  FILL_4050
timestamp 1713400504
transform 1 0 2232 0 -1 770
box -8 -3 16 105
use FILL  FILL_4051
timestamp 1713400504
transform 1 0 2200 0 -1 770
box -8 -3 16 105
use FILL  FILL_4052
timestamp 1713400504
transform 1 0 2192 0 -1 770
box -8 -3 16 105
use FILL  FILL_4053
timestamp 1713400504
transform 1 0 2184 0 -1 770
box -8 -3 16 105
use FILL  FILL_4054
timestamp 1713400504
transform 1 0 2176 0 -1 770
box -8 -3 16 105
use FILL  FILL_4055
timestamp 1713400504
transform 1 0 2168 0 -1 770
box -8 -3 16 105
use FILL  FILL_4056
timestamp 1713400504
transform 1 0 2128 0 -1 770
box -8 -3 16 105
use FILL  FILL_4057
timestamp 1713400504
transform 1 0 2120 0 -1 770
box -8 -3 16 105
use FILL  FILL_4058
timestamp 1713400504
transform 1 0 2112 0 -1 770
box -8 -3 16 105
use FILL  FILL_4059
timestamp 1713400504
transform 1 0 2104 0 -1 770
box -8 -3 16 105
use FILL  FILL_4060
timestamp 1713400504
transform 1 0 2096 0 -1 770
box -8 -3 16 105
use FILL  FILL_4061
timestamp 1713400504
transform 1 0 2088 0 -1 770
box -8 -3 16 105
use FILL  FILL_4062
timestamp 1713400504
transform 1 0 2080 0 -1 770
box -8 -3 16 105
use FILL  FILL_4063
timestamp 1713400504
transform 1 0 2048 0 -1 770
box -8 -3 16 105
use FILL  FILL_4064
timestamp 1713400504
transform 1 0 2040 0 -1 770
box -8 -3 16 105
use FILL  FILL_4065
timestamp 1713400504
transform 1 0 2032 0 -1 770
box -8 -3 16 105
use FILL  FILL_4066
timestamp 1713400504
transform 1 0 2024 0 -1 770
box -8 -3 16 105
use FILL  FILL_4067
timestamp 1713400504
transform 1 0 2016 0 -1 770
box -8 -3 16 105
use FILL  FILL_4068
timestamp 1713400504
transform 1 0 1992 0 -1 770
box -8 -3 16 105
use FILL  FILL_4069
timestamp 1713400504
transform 1 0 1984 0 -1 770
box -8 -3 16 105
use FILL  FILL_4070
timestamp 1713400504
transform 1 0 1976 0 -1 770
box -8 -3 16 105
use FILL  FILL_4071
timestamp 1713400504
transform 1 0 1968 0 -1 770
box -8 -3 16 105
use FILL  FILL_4072
timestamp 1713400504
transform 1 0 1960 0 -1 770
box -8 -3 16 105
use FILL  FILL_4073
timestamp 1713400504
transform 1 0 1952 0 -1 770
box -8 -3 16 105
use FILL  FILL_4074
timestamp 1713400504
transform 1 0 1912 0 -1 770
box -8 -3 16 105
use FILL  FILL_4075
timestamp 1713400504
transform 1 0 1904 0 -1 770
box -8 -3 16 105
use FILL  FILL_4076
timestamp 1713400504
transform 1 0 1896 0 -1 770
box -8 -3 16 105
use FILL  FILL_4077
timestamp 1713400504
transform 1 0 1888 0 -1 770
box -8 -3 16 105
use FILL  FILL_4078
timestamp 1713400504
transform 1 0 1880 0 -1 770
box -8 -3 16 105
use FILL  FILL_4079
timestamp 1713400504
transform 1 0 1872 0 -1 770
box -8 -3 16 105
use FILL  FILL_4080
timestamp 1713400504
transform 1 0 1864 0 -1 770
box -8 -3 16 105
use FILL  FILL_4081
timestamp 1713400504
transform 1 0 1824 0 -1 770
box -8 -3 16 105
use FILL  FILL_4082
timestamp 1713400504
transform 1 0 1816 0 -1 770
box -8 -3 16 105
use FILL  FILL_4083
timestamp 1713400504
transform 1 0 1808 0 -1 770
box -8 -3 16 105
use FILL  FILL_4084
timestamp 1713400504
transform 1 0 1800 0 -1 770
box -8 -3 16 105
use FILL  FILL_4085
timestamp 1713400504
transform 1 0 1792 0 -1 770
box -8 -3 16 105
use FILL  FILL_4086
timestamp 1713400504
transform 1 0 1688 0 -1 770
box -8 -3 16 105
use FILL  FILL_4087
timestamp 1713400504
transform 1 0 1680 0 -1 770
box -8 -3 16 105
use FILL  FILL_4088
timestamp 1713400504
transform 1 0 1672 0 -1 770
box -8 -3 16 105
use FILL  FILL_4089
timestamp 1713400504
transform 1 0 1664 0 -1 770
box -8 -3 16 105
use FILL  FILL_4090
timestamp 1713400504
transform 1 0 1656 0 -1 770
box -8 -3 16 105
use FILL  FILL_4091
timestamp 1713400504
transform 1 0 1648 0 -1 770
box -8 -3 16 105
use FILL  FILL_4092
timestamp 1713400504
transform 1 0 1624 0 -1 770
box -8 -3 16 105
use FILL  FILL_4093
timestamp 1713400504
transform 1 0 1616 0 -1 770
box -8 -3 16 105
use FILL  FILL_4094
timestamp 1713400504
transform 1 0 1608 0 -1 770
box -8 -3 16 105
use FILL  FILL_4095
timestamp 1713400504
transform 1 0 1600 0 -1 770
box -8 -3 16 105
use FILL  FILL_4096
timestamp 1713400504
transform 1 0 1592 0 -1 770
box -8 -3 16 105
use FILL  FILL_4097
timestamp 1713400504
transform 1 0 1584 0 -1 770
box -8 -3 16 105
use FILL  FILL_4098
timestamp 1713400504
transform 1 0 1576 0 -1 770
box -8 -3 16 105
use FILL  FILL_4099
timestamp 1713400504
transform 1 0 1544 0 -1 770
box -8 -3 16 105
use FILL  FILL_4100
timestamp 1713400504
transform 1 0 1536 0 -1 770
box -8 -3 16 105
use FILL  FILL_4101
timestamp 1713400504
transform 1 0 1528 0 -1 770
box -8 -3 16 105
use FILL  FILL_4102
timestamp 1713400504
transform 1 0 1520 0 -1 770
box -8 -3 16 105
use FILL  FILL_4103
timestamp 1713400504
transform 1 0 1512 0 -1 770
box -8 -3 16 105
use FILL  FILL_4104
timestamp 1713400504
transform 1 0 1504 0 -1 770
box -8 -3 16 105
use FILL  FILL_4105
timestamp 1713400504
transform 1 0 1496 0 -1 770
box -8 -3 16 105
use FILL  FILL_4106
timestamp 1713400504
transform 1 0 1488 0 -1 770
box -8 -3 16 105
use FILL  FILL_4107
timestamp 1713400504
transform 1 0 1480 0 -1 770
box -8 -3 16 105
use FILL  FILL_4108
timestamp 1713400504
transform 1 0 1472 0 -1 770
box -8 -3 16 105
use FILL  FILL_4109
timestamp 1713400504
transform 1 0 1464 0 -1 770
box -8 -3 16 105
use FILL  FILL_4110
timestamp 1713400504
transform 1 0 1456 0 -1 770
box -8 -3 16 105
use FILL  FILL_4111
timestamp 1713400504
transform 1 0 1448 0 -1 770
box -8 -3 16 105
use FILL  FILL_4112
timestamp 1713400504
transform 1 0 1440 0 -1 770
box -8 -3 16 105
use FILL  FILL_4113
timestamp 1713400504
transform 1 0 1432 0 -1 770
box -8 -3 16 105
use FILL  FILL_4114
timestamp 1713400504
transform 1 0 1424 0 -1 770
box -8 -3 16 105
use FILL  FILL_4115
timestamp 1713400504
transform 1 0 1416 0 -1 770
box -8 -3 16 105
use FILL  FILL_4116
timestamp 1713400504
transform 1 0 1408 0 -1 770
box -8 -3 16 105
use FILL  FILL_4117
timestamp 1713400504
transform 1 0 1400 0 -1 770
box -8 -3 16 105
use FILL  FILL_4118
timestamp 1713400504
transform 1 0 1392 0 -1 770
box -8 -3 16 105
use FILL  FILL_4119
timestamp 1713400504
transform 1 0 1384 0 -1 770
box -8 -3 16 105
use FILL  FILL_4120
timestamp 1713400504
transform 1 0 1376 0 -1 770
box -8 -3 16 105
use FILL  FILL_4121
timestamp 1713400504
transform 1 0 1368 0 -1 770
box -8 -3 16 105
use FILL  FILL_4122
timestamp 1713400504
transform 1 0 1360 0 -1 770
box -8 -3 16 105
use FILL  FILL_4123
timestamp 1713400504
transform 1 0 1352 0 -1 770
box -8 -3 16 105
use FILL  FILL_4124
timestamp 1713400504
transform 1 0 1344 0 -1 770
box -8 -3 16 105
use FILL  FILL_4125
timestamp 1713400504
transform 1 0 1336 0 -1 770
box -8 -3 16 105
use FILL  FILL_4126
timestamp 1713400504
transform 1 0 1328 0 -1 770
box -8 -3 16 105
use FILL  FILL_4127
timestamp 1713400504
transform 1 0 1320 0 -1 770
box -8 -3 16 105
use FILL  FILL_4128
timestamp 1713400504
transform 1 0 1312 0 -1 770
box -8 -3 16 105
use FILL  FILL_4129
timestamp 1713400504
transform 1 0 1304 0 -1 770
box -8 -3 16 105
use FILL  FILL_4130
timestamp 1713400504
transform 1 0 1296 0 -1 770
box -8 -3 16 105
use FILL  FILL_4131
timestamp 1713400504
transform 1 0 1288 0 -1 770
box -8 -3 16 105
use FILL  FILL_4132
timestamp 1713400504
transform 1 0 1248 0 -1 770
box -8 -3 16 105
use FILL  FILL_4133
timestamp 1713400504
transform 1 0 1240 0 -1 770
box -8 -3 16 105
use FILL  FILL_4134
timestamp 1713400504
transform 1 0 1232 0 -1 770
box -8 -3 16 105
use FILL  FILL_4135
timestamp 1713400504
transform 1 0 1224 0 -1 770
box -8 -3 16 105
use FILL  FILL_4136
timestamp 1713400504
transform 1 0 1216 0 -1 770
box -8 -3 16 105
use FILL  FILL_4137
timestamp 1713400504
transform 1 0 1208 0 -1 770
box -8 -3 16 105
use FILL  FILL_4138
timestamp 1713400504
transform 1 0 1200 0 -1 770
box -8 -3 16 105
use FILL  FILL_4139
timestamp 1713400504
transform 1 0 1192 0 -1 770
box -8 -3 16 105
use FILL  FILL_4140
timestamp 1713400504
transform 1 0 1184 0 -1 770
box -8 -3 16 105
use FILL  FILL_4141
timestamp 1713400504
transform 1 0 1152 0 -1 770
box -8 -3 16 105
use FILL  FILL_4142
timestamp 1713400504
transform 1 0 1144 0 -1 770
box -8 -3 16 105
use FILL  FILL_4143
timestamp 1713400504
transform 1 0 1136 0 -1 770
box -8 -3 16 105
use FILL  FILL_4144
timestamp 1713400504
transform 1 0 1128 0 -1 770
box -8 -3 16 105
use FILL  FILL_4145
timestamp 1713400504
transform 1 0 1120 0 -1 770
box -8 -3 16 105
use FILL  FILL_4146
timestamp 1713400504
transform 1 0 1112 0 -1 770
box -8 -3 16 105
use FILL  FILL_4147
timestamp 1713400504
transform 1 0 1104 0 -1 770
box -8 -3 16 105
use FILL  FILL_4148
timestamp 1713400504
transform 1 0 1072 0 -1 770
box -8 -3 16 105
use FILL  FILL_4149
timestamp 1713400504
transform 1 0 1064 0 -1 770
box -8 -3 16 105
use FILL  FILL_4150
timestamp 1713400504
transform 1 0 1056 0 -1 770
box -8 -3 16 105
use FILL  FILL_4151
timestamp 1713400504
transform 1 0 1048 0 -1 770
box -8 -3 16 105
use FILL  FILL_4152
timestamp 1713400504
transform 1 0 944 0 -1 770
box -8 -3 16 105
use FILL  FILL_4153
timestamp 1713400504
transform 1 0 936 0 -1 770
box -8 -3 16 105
use FILL  FILL_4154
timestamp 1713400504
transform 1 0 928 0 -1 770
box -8 -3 16 105
use FILL  FILL_4155
timestamp 1713400504
transform 1 0 920 0 -1 770
box -8 -3 16 105
use FILL  FILL_4156
timestamp 1713400504
transform 1 0 912 0 -1 770
box -8 -3 16 105
use FILL  FILL_4157
timestamp 1713400504
transform 1 0 904 0 -1 770
box -8 -3 16 105
use FILL  FILL_4158
timestamp 1713400504
transform 1 0 864 0 -1 770
box -8 -3 16 105
use FILL  FILL_4159
timestamp 1713400504
transform 1 0 856 0 -1 770
box -8 -3 16 105
use FILL  FILL_4160
timestamp 1713400504
transform 1 0 848 0 -1 770
box -8 -3 16 105
use FILL  FILL_4161
timestamp 1713400504
transform 1 0 840 0 -1 770
box -8 -3 16 105
use FILL  FILL_4162
timestamp 1713400504
transform 1 0 832 0 -1 770
box -8 -3 16 105
use FILL  FILL_4163
timestamp 1713400504
transform 1 0 824 0 -1 770
box -8 -3 16 105
use FILL  FILL_4164
timestamp 1713400504
transform 1 0 792 0 -1 770
box -8 -3 16 105
use FILL  FILL_4165
timestamp 1713400504
transform 1 0 784 0 -1 770
box -8 -3 16 105
use FILL  FILL_4166
timestamp 1713400504
transform 1 0 776 0 -1 770
box -8 -3 16 105
use FILL  FILL_4167
timestamp 1713400504
transform 1 0 768 0 -1 770
box -8 -3 16 105
use FILL  FILL_4168
timestamp 1713400504
transform 1 0 760 0 -1 770
box -8 -3 16 105
use FILL  FILL_4169
timestamp 1713400504
transform 1 0 736 0 -1 770
box -8 -3 16 105
use FILL  FILL_4170
timestamp 1713400504
transform 1 0 728 0 -1 770
box -8 -3 16 105
use FILL  FILL_4171
timestamp 1713400504
transform 1 0 720 0 -1 770
box -8 -3 16 105
use FILL  FILL_4172
timestamp 1713400504
transform 1 0 712 0 -1 770
box -8 -3 16 105
use FILL  FILL_4173
timestamp 1713400504
transform 1 0 672 0 -1 770
box -8 -3 16 105
use FILL  FILL_4174
timestamp 1713400504
transform 1 0 664 0 -1 770
box -8 -3 16 105
use FILL  FILL_4175
timestamp 1713400504
transform 1 0 656 0 -1 770
box -8 -3 16 105
use FILL  FILL_4176
timestamp 1713400504
transform 1 0 648 0 -1 770
box -8 -3 16 105
use FILL  FILL_4177
timestamp 1713400504
transform 1 0 640 0 -1 770
box -8 -3 16 105
use FILL  FILL_4178
timestamp 1713400504
transform 1 0 632 0 -1 770
box -8 -3 16 105
use FILL  FILL_4179
timestamp 1713400504
transform 1 0 624 0 -1 770
box -8 -3 16 105
use FILL  FILL_4180
timestamp 1713400504
transform 1 0 584 0 -1 770
box -8 -3 16 105
use FILL  FILL_4181
timestamp 1713400504
transform 1 0 576 0 -1 770
box -8 -3 16 105
use FILL  FILL_4182
timestamp 1713400504
transform 1 0 568 0 -1 770
box -8 -3 16 105
use FILL  FILL_4183
timestamp 1713400504
transform 1 0 560 0 -1 770
box -8 -3 16 105
use FILL  FILL_4184
timestamp 1713400504
transform 1 0 552 0 -1 770
box -8 -3 16 105
use FILL  FILL_4185
timestamp 1713400504
transform 1 0 544 0 -1 770
box -8 -3 16 105
use FILL  FILL_4186
timestamp 1713400504
transform 1 0 504 0 -1 770
box -8 -3 16 105
use FILL  FILL_4187
timestamp 1713400504
transform 1 0 496 0 -1 770
box -8 -3 16 105
use FILL  FILL_4188
timestamp 1713400504
transform 1 0 488 0 -1 770
box -8 -3 16 105
use FILL  FILL_4189
timestamp 1713400504
transform 1 0 480 0 -1 770
box -8 -3 16 105
use FILL  FILL_4190
timestamp 1713400504
transform 1 0 472 0 -1 770
box -8 -3 16 105
use FILL  FILL_4191
timestamp 1713400504
transform 1 0 464 0 -1 770
box -8 -3 16 105
use FILL  FILL_4192
timestamp 1713400504
transform 1 0 456 0 -1 770
box -8 -3 16 105
use FILL  FILL_4193
timestamp 1713400504
transform 1 0 448 0 -1 770
box -8 -3 16 105
use FILL  FILL_4194
timestamp 1713400504
transform 1 0 408 0 -1 770
box -8 -3 16 105
use FILL  FILL_4195
timestamp 1713400504
transform 1 0 400 0 -1 770
box -8 -3 16 105
use FILL  FILL_4196
timestamp 1713400504
transform 1 0 392 0 -1 770
box -8 -3 16 105
use FILL  FILL_4197
timestamp 1713400504
transform 1 0 384 0 -1 770
box -8 -3 16 105
use FILL  FILL_4198
timestamp 1713400504
transform 1 0 376 0 -1 770
box -8 -3 16 105
use FILL  FILL_4199
timestamp 1713400504
transform 1 0 368 0 -1 770
box -8 -3 16 105
use FILL  FILL_4200
timestamp 1713400504
transform 1 0 328 0 -1 770
box -8 -3 16 105
use FILL  FILL_4201
timestamp 1713400504
transform 1 0 320 0 -1 770
box -8 -3 16 105
use FILL  FILL_4202
timestamp 1713400504
transform 1 0 312 0 -1 770
box -8 -3 16 105
use FILL  FILL_4203
timestamp 1713400504
transform 1 0 304 0 -1 770
box -8 -3 16 105
use FILL  FILL_4204
timestamp 1713400504
transform 1 0 296 0 -1 770
box -8 -3 16 105
use FILL  FILL_4205
timestamp 1713400504
transform 1 0 288 0 -1 770
box -8 -3 16 105
use FILL  FILL_4206
timestamp 1713400504
transform 1 0 256 0 -1 770
box -8 -3 16 105
use FILL  FILL_4207
timestamp 1713400504
transform 1 0 248 0 -1 770
box -8 -3 16 105
use FILL  FILL_4208
timestamp 1713400504
transform 1 0 240 0 -1 770
box -8 -3 16 105
use FILL  FILL_4209
timestamp 1713400504
transform 1 0 232 0 -1 770
box -8 -3 16 105
use FILL  FILL_4210
timestamp 1713400504
transform 1 0 208 0 -1 770
box -8 -3 16 105
use FILL  FILL_4211
timestamp 1713400504
transform 1 0 200 0 -1 770
box -8 -3 16 105
use FILL  FILL_4212
timestamp 1713400504
transform 1 0 192 0 -1 770
box -8 -3 16 105
use FILL  FILL_4213
timestamp 1713400504
transform 1 0 184 0 -1 770
box -8 -3 16 105
use FILL  FILL_4214
timestamp 1713400504
transform 1 0 176 0 -1 770
box -8 -3 16 105
use FILL  FILL_4215
timestamp 1713400504
transform 1 0 168 0 -1 770
box -8 -3 16 105
use FILL  FILL_4216
timestamp 1713400504
transform 1 0 160 0 -1 770
box -8 -3 16 105
use FILL  FILL_4217
timestamp 1713400504
transform 1 0 152 0 -1 770
box -8 -3 16 105
use FILL  FILL_4218
timestamp 1713400504
transform 1 0 144 0 -1 770
box -8 -3 16 105
use FILL  FILL_4219
timestamp 1713400504
transform 1 0 136 0 -1 770
box -8 -3 16 105
use FILL  FILL_4220
timestamp 1713400504
transform 1 0 128 0 -1 770
box -8 -3 16 105
use FILL  FILL_4221
timestamp 1713400504
transform 1 0 120 0 -1 770
box -8 -3 16 105
use FILL  FILL_4222
timestamp 1713400504
transform 1 0 112 0 -1 770
box -8 -3 16 105
use FILL  FILL_4223
timestamp 1713400504
transform 1 0 104 0 -1 770
box -8 -3 16 105
use FILL  FILL_4224
timestamp 1713400504
transform 1 0 96 0 -1 770
box -8 -3 16 105
use FILL  FILL_4225
timestamp 1713400504
transform 1 0 88 0 -1 770
box -8 -3 16 105
use FILL  FILL_4226
timestamp 1713400504
transform 1 0 80 0 -1 770
box -8 -3 16 105
use FILL  FILL_4227
timestamp 1713400504
transform 1 0 72 0 -1 770
box -8 -3 16 105
use FILL  FILL_4228
timestamp 1713400504
transform 1 0 3008 0 1 570
box -8 -3 16 105
use FILL  FILL_4229
timestamp 1713400504
transform 1 0 3000 0 1 570
box -8 -3 16 105
use FILL  FILL_4230
timestamp 1713400504
transform 1 0 2992 0 1 570
box -8 -3 16 105
use FILL  FILL_4231
timestamp 1713400504
transform 1 0 2984 0 1 570
box -8 -3 16 105
use FILL  FILL_4232
timestamp 1713400504
transform 1 0 2944 0 1 570
box -8 -3 16 105
use FILL  FILL_4233
timestamp 1713400504
transform 1 0 2936 0 1 570
box -8 -3 16 105
use FILL  FILL_4234
timestamp 1713400504
transform 1 0 2928 0 1 570
box -8 -3 16 105
use FILL  FILL_4235
timestamp 1713400504
transform 1 0 2904 0 1 570
box -8 -3 16 105
use FILL  FILL_4236
timestamp 1713400504
transform 1 0 2896 0 1 570
box -8 -3 16 105
use FILL  FILL_4237
timestamp 1713400504
transform 1 0 2888 0 1 570
box -8 -3 16 105
use FILL  FILL_4238
timestamp 1713400504
transform 1 0 2880 0 1 570
box -8 -3 16 105
use FILL  FILL_4239
timestamp 1713400504
transform 1 0 2872 0 1 570
box -8 -3 16 105
use FILL  FILL_4240
timestamp 1713400504
transform 1 0 2832 0 1 570
box -8 -3 16 105
use FILL  FILL_4241
timestamp 1713400504
transform 1 0 2824 0 1 570
box -8 -3 16 105
use FILL  FILL_4242
timestamp 1713400504
transform 1 0 2816 0 1 570
box -8 -3 16 105
use FILL  FILL_4243
timestamp 1713400504
transform 1 0 2808 0 1 570
box -8 -3 16 105
use FILL  FILL_4244
timestamp 1713400504
transform 1 0 2768 0 1 570
box -8 -3 16 105
use FILL  FILL_4245
timestamp 1713400504
transform 1 0 2760 0 1 570
box -8 -3 16 105
use FILL  FILL_4246
timestamp 1713400504
transform 1 0 2752 0 1 570
box -8 -3 16 105
use FILL  FILL_4247
timestamp 1713400504
transform 1 0 2744 0 1 570
box -8 -3 16 105
use FILL  FILL_4248
timestamp 1713400504
transform 1 0 2704 0 1 570
box -8 -3 16 105
use FILL  FILL_4249
timestamp 1713400504
transform 1 0 2696 0 1 570
box -8 -3 16 105
use FILL  FILL_4250
timestamp 1713400504
transform 1 0 2688 0 1 570
box -8 -3 16 105
use FILL  FILL_4251
timestamp 1713400504
transform 1 0 2680 0 1 570
box -8 -3 16 105
use FILL  FILL_4252
timestamp 1713400504
transform 1 0 2672 0 1 570
box -8 -3 16 105
use FILL  FILL_4253
timestamp 1713400504
transform 1 0 2632 0 1 570
box -8 -3 16 105
use FILL  FILL_4254
timestamp 1713400504
transform 1 0 2624 0 1 570
box -8 -3 16 105
use FILL  FILL_4255
timestamp 1713400504
transform 1 0 2616 0 1 570
box -8 -3 16 105
use FILL  FILL_4256
timestamp 1713400504
transform 1 0 2608 0 1 570
box -8 -3 16 105
use FILL  FILL_4257
timestamp 1713400504
transform 1 0 2600 0 1 570
box -8 -3 16 105
use FILL  FILL_4258
timestamp 1713400504
transform 1 0 2560 0 1 570
box -8 -3 16 105
use FILL  FILL_4259
timestamp 1713400504
transform 1 0 2552 0 1 570
box -8 -3 16 105
use FILL  FILL_4260
timestamp 1713400504
transform 1 0 2544 0 1 570
box -8 -3 16 105
use FILL  FILL_4261
timestamp 1713400504
transform 1 0 2440 0 1 570
box -8 -3 16 105
use FILL  FILL_4262
timestamp 1713400504
transform 1 0 2336 0 1 570
box -8 -3 16 105
use FILL  FILL_4263
timestamp 1713400504
transform 1 0 2328 0 1 570
box -8 -3 16 105
use FILL  FILL_4264
timestamp 1713400504
transform 1 0 2320 0 1 570
box -8 -3 16 105
use FILL  FILL_4265
timestamp 1713400504
transform 1 0 2288 0 1 570
box -8 -3 16 105
use FILL  FILL_4266
timestamp 1713400504
transform 1 0 2280 0 1 570
box -8 -3 16 105
use FILL  FILL_4267
timestamp 1713400504
transform 1 0 2272 0 1 570
box -8 -3 16 105
use FILL  FILL_4268
timestamp 1713400504
transform 1 0 2264 0 1 570
box -8 -3 16 105
use FILL  FILL_4269
timestamp 1713400504
transform 1 0 2224 0 1 570
box -8 -3 16 105
use FILL  FILL_4270
timestamp 1713400504
transform 1 0 2216 0 1 570
box -8 -3 16 105
use FILL  FILL_4271
timestamp 1713400504
transform 1 0 2208 0 1 570
box -8 -3 16 105
use FILL  FILL_4272
timestamp 1713400504
transform 1 0 2200 0 1 570
box -8 -3 16 105
use FILL  FILL_4273
timestamp 1713400504
transform 1 0 2192 0 1 570
box -8 -3 16 105
use FILL  FILL_4274
timestamp 1713400504
transform 1 0 2168 0 1 570
box -8 -3 16 105
use FILL  FILL_4275
timestamp 1713400504
transform 1 0 2160 0 1 570
box -8 -3 16 105
use FILL  FILL_4276
timestamp 1713400504
transform 1 0 2152 0 1 570
box -8 -3 16 105
use FILL  FILL_4277
timestamp 1713400504
transform 1 0 2128 0 1 570
box -8 -3 16 105
use FILL  FILL_4278
timestamp 1713400504
transform 1 0 2120 0 1 570
box -8 -3 16 105
use FILL  FILL_4279
timestamp 1713400504
transform 1 0 2112 0 1 570
box -8 -3 16 105
use FILL  FILL_4280
timestamp 1713400504
transform 1 0 2088 0 1 570
box -8 -3 16 105
use FILL  FILL_4281
timestamp 1713400504
transform 1 0 2080 0 1 570
box -8 -3 16 105
use FILL  FILL_4282
timestamp 1713400504
transform 1 0 2072 0 1 570
box -8 -3 16 105
use FILL  FILL_4283
timestamp 1713400504
transform 1 0 1968 0 1 570
box -8 -3 16 105
use FILL  FILL_4284
timestamp 1713400504
transform 1 0 1960 0 1 570
box -8 -3 16 105
use FILL  FILL_4285
timestamp 1713400504
transform 1 0 1856 0 1 570
box -8 -3 16 105
use FILL  FILL_4286
timestamp 1713400504
transform 1 0 1848 0 1 570
box -8 -3 16 105
use FILL  FILL_4287
timestamp 1713400504
transform 1 0 1840 0 1 570
box -8 -3 16 105
use FILL  FILL_4288
timestamp 1713400504
transform 1 0 1800 0 1 570
box -8 -3 16 105
use FILL  FILL_4289
timestamp 1713400504
transform 1 0 1792 0 1 570
box -8 -3 16 105
use FILL  FILL_4290
timestamp 1713400504
transform 1 0 1784 0 1 570
box -8 -3 16 105
use FILL  FILL_4291
timestamp 1713400504
transform 1 0 1776 0 1 570
box -8 -3 16 105
use FILL  FILL_4292
timestamp 1713400504
transform 1 0 1768 0 1 570
box -8 -3 16 105
use FILL  FILL_4293
timestamp 1713400504
transform 1 0 1760 0 1 570
box -8 -3 16 105
use FILL  FILL_4294
timestamp 1713400504
transform 1 0 1720 0 1 570
box -8 -3 16 105
use FILL  FILL_4295
timestamp 1713400504
transform 1 0 1712 0 1 570
box -8 -3 16 105
use FILL  FILL_4296
timestamp 1713400504
transform 1 0 1704 0 1 570
box -8 -3 16 105
use FILL  FILL_4297
timestamp 1713400504
transform 1 0 1640 0 1 570
box -8 -3 16 105
use FILL  FILL_4298
timestamp 1713400504
transform 1 0 1632 0 1 570
box -8 -3 16 105
use FILL  FILL_4299
timestamp 1713400504
transform 1 0 1624 0 1 570
box -8 -3 16 105
use FILL  FILL_4300
timestamp 1713400504
transform 1 0 1616 0 1 570
box -8 -3 16 105
use FILL  FILL_4301
timestamp 1713400504
transform 1 0 1576 0 1 570
box -8 -3 16 105
use FILL  FILL_4302
timestamp 1713400504
transform 1 0 1568 0 1 570
box -8 -3 16 105
use FILL  FILL_4303
timestamp 1713400504
transform 1 0 1560 0 1 570
box -8 -3 16 105
use FILL  FILL_4304
timestamp 1713400504
transform 1 0 1552 0 1 570
box -8 -3 16 105
use FILL  FILL_4305
timestamp 1713400504
transform 1 0 1544 0 1 570
box -8 -3 16 105
use FILL  FILL_4306
timestamp 1713400504
transform 1 0 1536 0 1 570
box -8 -3 16 105
use FILL  FILL_4307
timestamp 1713400504
transform 1 0 1496 0 1 570
box -8 -3 16 105
use FILL  FILL_4308
timestamp 1713400504
transform 1 0 1488 0 1 570
box -8 -3 16 105
use FILL  FILL_4309
timestamp 1713400504
transform 1 0 1480 0 1 570
box -8 -3 16 105
use FILL  FILL_4310
timestamp 1713400504
transform 1 0 1472 0 1 570
box -8 -3 16 105
use FILL  FILL_4311
timestamp 1713400504
transform 1 0 1408 0 1 570
box -8 -3 16 105
use FILL  FILL_4312
timestamp 1713400504
transform 1 0 1400 0 1 570
box -8 -3 16 105
use FILL  FILL_4313
timestamp 1713400504
transform 1 0 1392 0 1 570
box -8 -3 16 105
use FILL  FILL_4314
timestamp 1713400504
transform 1 0 1352 0 1 570
box -8 -3 16 105
use FILL  FILL_4315
timestamp 1713400504
transform 1 0 1344 0 1 570
box -8 -3 16 105
use FILL  FILL_4316
timestamp 1713400504
transform 1 0 1336 0 1 570
box -8 -3 16 105
use FILL  FILL_4317
timestamp 1713400504
transform 1 0 1328 0 1 570
box -8 -3 16 105
use FILL  FILL_4318
timestamp 1713400504
transform 1 0 1320 0 1 570
box -8 -3 16 105
use FILL  FILL_4319
timestamp 1713400504
transform 1 0 1312 0 1 570
box -8 -3 16 105
use FILL  FILL_4320
timestamp 1713400504
transform 1 0 1304 0 1 570
box -8 -3 16 105
use FILL  FILL_4321
timestamp 1713400504
transform 1 0 1296 0 1 570
box -8 -3 16 105
use FILL  FILL_4322
timestamp 1713400504
transform 1 0 1256 0 1 570
box -8 -3 16 105
use FILL  FILL_4323
timestamp 1713400504
transform 1 0 1248 0 1 570
box -8 -3 16 105
use FILL  FILL_4324
timestamp 1713400504
transform 1 0 1240 0 1 570
box -8 -3 16 105
use FILL  FILL_4325
timestamp 1713400504
transform 1 0 1232 0 1 570
box -8 -3 16 105
use FILL  FILL_4326
timestamp 1713400504
transform 1 0 1224 0 1 570
box -8 -3 16 105
use FILL  FILL_4327
timestamp 1713400504
transform 1 0 1216 0 1 570
box -8 -3 16 105
use FILL  FILL_4328
timestamp 1713400504
transform 1 0 1208 0 1 570
box -8 -3 16 105
use FILL  FILL_4329
timestamp 1713400504
transform 1 0 1200 0 1 570
box -8 -3 16 105
use FILL  FILL_4330
timestamp 1713400504
transform 1 0 1152 0 1 570
box -8 -3 16 105
use FILL  FILL_4331
timestamp 1713400504
transform 1 0 1144 0 1 570
box -8 -3 16 105
use FILL  FILL_4332
timestamp 1713400504
transform 1 0 1136 0 1 570
box -8 -3 16 105
use FILL  FILL_4333
timestamp 1713400504
transform 1 0 1128 0 1 570
box -8 -3 16 105
use FILL  FILL_4334
timestamp 1713400504
transform 1 0 1120 0 1 570
box -8 -3 16 105
use FILL  FILL_4335
timestamp 1713400504
transform 1 0 1112 0 1 570
box -8 -3 16 105
use FILL  FILL_4336
timestamp 1713400504
transform 1 0 1104 0 1 570
box -8 -3 16 105
use FILL  FILL_4337
timestamp 1713400504
transform 1 0 1096 0 1 570
box -8 -3 16 105
use FILL  FILL_4338
timestamp 1713400504
transform 1 0 1064 0 1 570
box -8 -3 16 105
use FILL  FILL_4339
timestamp 1713400504
transform 1 0 1056 0 1 570
box -8 -3 16 105
use FILL  FILL_4340
timestamp 1713400504
transform 1 0 1048 0 1 570
box -8 -3 16 105
use FILL  FILL_4341
timestamp 1713400504
transform 1 0 1040 0 1 570
box -8 -3 16 105
use FILL  FILL_4342
timestamp 1713400504
transform 1 0 1032 0 1 570
box -8 -3 16 105
use FILL  FILL_4343
timestamp 1713400504
transform 1 0 1024 0 1 570
box -8 -3 16 105
use FILL  FILL_4344
timestamp 1713400504
transform 1 0 1016 0 1 570
box -8 -3 16 105
use FILL  FILL_4345
timestamp 1713400504
transform 1 0 1008 0 1 570
box -8 -3 16 105
use FILL  FILL_4346
timestamp 1713400504
transform 1 0 1000 0 1 570
box -8 -3 16 105
use FILL  FILL_4347
timestamp 1713400504
transform 1 0 960 0 1 570
box -8 -3 16 105
use FILL  FILL_4348
timestamp 1713400504
transform 1 0 952 0 1 570
box -8 -3 16 105
use FILL  FILL_4349
timestamp 1713400504
transform 1 0 944 0 1 570
box -8 -3 16 105
use FILL  FILL_4350
timestamp 1713400504
transform 1 0 936 0 1 570
box -8 -3 16 105
use FILL  FILL_4351
timestamp 1713400504
transform 1 0 928 0 1 570
box -8 -3 16 105
use FILL  FILL_4352
timestamp 1713400504
transform 1 0 920 0 1 570
box -8 -3 16 105
use FILL  FILL_4353
timestamp 1713400504
transform 1 0 912 0 1 570
box -8 -3 16 105
use FILL  FILL_4354
timestamp 1713400504
transform 1 0 904 0 1 570
box -8 -3 16 105
use FILL  FILL_4355
timestamp 1713400504
transform 1 0 896 0 1 570
box -8 -3 16 105
use FILL  FILL_4356
timestamp 1713400504
transform 1 0 872 0 1 570
box -8 -3 16 105
use FILL  FILL_4357
timestamp 1713400504
transform 1 0 864 0 1 570
box -8 -3 16 105
use FILL  FILL_4358
timestamp 1713400504
transform 1 0 856 0 1 570
box -8 -3 16 105
use FILL  FILL_4359
timestamp 1713400504
transform 1 0 848 0 1 570
box -8 -3 16 105
use FILL  FILL_4360
timestamp 1713400504
transform 1 0 840 0 1 570
box -8 -3 16 105
use FILL  FILL_4361
timestamp 1713400504
transform 1 0 832 0 1 570
box -8 -3 16 105
use FILL  FILL_4362
timestamp 1713400504
transform 1 0 824 0 1 570
box -8 -3 16 105
use FILL  FILL_4363
timestamp 1713400504
transform 1 0 784 0 1 570
box -8 -3 16 105
use FILL  FILL_4364
timestamp 1713400504
transform 1 0 776 0 1 570
box -8 -3 16 105
use FILL  FILL_4365
timestamp 1713400504
transform 1 0 768 0 1 570
box -8 -3 16 105
use FILL  FILL_4366
timestamp 1713400504
transform 1 0 760 0 1 570
box -8 -3 16 105
use FILL  FILL_4367
timestamp 1713400504
transform 1 0 752 0 1 570
box -8 -3 16 105
use FILL  FILL_4368
timestamp 1713400504
transform 1 0 744 0 1 570
box -8 -3 16 105
use FILL  FILL_4369
timestamp 1713400504
transform 1 0 736 0 1 570
box -8 -3 16 105
use FILL  FILL_4370
timestamp 1713400504
transform 1 0 696 0 1 570
box -8 -3 16 105
use FILL  FILL_4371
timestamp 1713400504
transform 1 0 688 0 1 570
box -8 -3 16 105
use FILL  FILL_4372
timestamp 1713400504
transform 1 0 680 0 1 570
box -8 -3 16 105
use FILL  FILL_4373
timestamp 1713400504
transform 1 0 672 0 1 570
box -8 -3 16 105
use FILL  FILL_4374
timestamp 1713400504
transform 1 0 648 0 1 570
box -8 -3 16 105
use FILL  FILL_4375
timestamp 1713400504
transform 1 0 640 0 1 570
box -8 -3 16 105
use FILL  FILL_4376
timestamp 1713400504
transform 1 0 632 0 1 570
box -8 -3 16 105
use FILL  FILL_4377
timestamp 1713400504
transform 1 0 624 0 1 570
box -8 -3 16 105
use FILL  FILL_4378
timestamp 1713400504
transform 1 0 592 0 1 570
box -8 -3 16 105
use FILL  FILL_4379
timestamp 1713400504
transform 1 0 584 0 1 570
box -8 -3 16 105
use FILL  FILL_4380
timestamp 1713400504
transform 1 0 576 0 1 570
box -8 -3 16 105
use FILL  FILL_4381
timestamp 1713400504
transform 1 0 568 0 1 570
box -8 -3 16 105
use FILL  FILL_4382
timestamp 1713400504
transform 1 0 560 0 1 570
box -8 -3 16 105
use FILL  FILL_4383
timestamp 1713400504
transform 1 0 520 0 1 570
box -8 -3 16 105
use FILL  FILL_4384
timestamp 1713400504
transform 1 0 512 0 1 570
box -8 -3 16 105
use FILL  FILL_4385
timestamp 1713400504
transform 1 0 504 0 1 570
box -8 -3 16 105
use FILL  FILL_4386
timestamp 1713400504
transform 1 0 400 0 1 570
box -8 -3 16 105
use FILL  FILL_4387
timestamp 1713400504
transform 1 0 392 0 1 570
box -8 -3 16 105
use FILL  FILL_4388
timestamp 1713400504
transform 1 0 384 0 1 570
box -8 -3 16 105
use FILL  FILL_4389
timestamp 1713400504
transform 1 0 376 0 1 570
box -8 -3 16 105
use FILL  FILL_4390
timestamp 1713400504
transform 1 0 368 0 1 570
box -8 -3 16 105
use FILL  FILL_4391
timestamp 1713400504
transform 1 0 320 0 1 570
box -8 -3 16 105
use FILL  FILL_4392
timestamp 1713400504
transform 1 0 312 0 1 570
box -8 -3 16 105
use FILL  FILL_4393
timestamp 1713400504
transform 1 0 304 0 1 570
box -8 -3 16 105
use FILL  FILL_4394
timestamp 1713400504
transform 1 0 296 0 1 570
box -8 -3 16 105
use FILL  FILL_4395
timestamp 1713400504
transform 1 0 288 0 1 570
box -8 -3 16 105
use FILL  FILL_4396
timestamp 1713400504
transform 1 0 280 0 1 570
box -8 -3 16 105
use FILL  FILL_4397
timestamp 1713400504
transform 1 0 248 0 1 570
box -8 -3 16 105
use FILL  FILL_4398
timestamp 1713400504
transform 1 0 240 0 1 570
box -8 -3 16 105
use FILL  FILL_4399
timestamp 1713400504
transform 1 0 232 0 1 570
box -8 -3 16 105
use FILL  FILL_4400
timestamp 1713400504
transform 1 0 192 0 1 570
box -8 -3 16 105
use FILL  FILL_4401
timestamp 1713400504
transform 1 0 184 0 1 570
box -8 -3 16 105
use FILL  FILL_4402
timestamp 1713400504
transform 1 0 176 0 1 570
box -8 -3 16 105
use FILL  FILL_4403
timestamp 1713400504
transform 1 0 72 0 1 570
box -8 -3 16 105
use FILL  FILL_4404
timestamp 1713400504
transform 1 0 3008 0 -1 570
box -8 -3 16 105
use FILL  FILL_4405
timestamp 1713400504
transform 1 0 3000 0 -1 570
box -8 -3 16 105
use FILL  FILL_4406
timestamp 1713400504
transform 1 0 2976 0 -1 570
box -8 -3 16 105
use FILL  FILL_4407
timestamp 1713400504
transform 1 0 2968 0 -1 570
box -8 -3 16 105
use FILL  FILL_4408
timestamp 1713400504
transform 1 0 2960 0 -1 570
box -8 -3 16 105
use FILL  FILL_4409
timestamp 1713400504
transform 1 0 2952 0 -1 570
box -8 -3 16 105
use FILL  FILL_4410
timestamp 1713400504
transform 1 0 2912 0 -1 570
box -8 -3 16 105
use FILL  FILL_4411
timestamp 1713400504
transform 1 0 2904 0 -1 570
box -8 -3 16 105
use FILL  FILL_4412
timestamp 1713400504
transform 1 0 2896 0 -1 570
box -8 -3 16 105
use FILL  FILL_4413
timestamp 1713400504
transform 1 0 2888 0 -1 570
box -8 -3 16 105
use FILL  FILL_4414
timestamp 1713400504
transform 1 0 2864 0 -1 570
box -8 -3 16 105
use FILL  FILL_4415
timestamp 1713400504
transform 1 0 2856 0 -1 570
box -8 -3 16 105
use FILL  FILL_4416
timestamp 1713400504
transform 1 0 2752 0 -1 570
box -8 -3 16 105
use FILL  FILL_4417
timestamp 1713400504
transform 1 0 2744 0 -1 570
box -8 -3 16 105
use FILL  FILL_4418
timestamp 1713400504
transform 1 0 2736 0 -1 570
box -8 -3 16 105
use FILL  FILL_4419
timestamp 1713400504
transform 1 0 2696 0 -1 570
box -8 -3 16 105
use FILL  FILL_4420
timestamp 1713400504
transform 1 0 2688 0 -1 570
box -8 -3 16 105
use FILL  FILL_4421
timestamp 1713400504
transform 1 0 2680 0 -1 570
box -8 -3 16 105
use FILL  FILL_4422
timestamp 1713400504
transform 1 0 2672 0 -1 570
box -8 -3 16 105
use FILL  FILL_4423
timestamp 1713400504
transform 1 0 2664 0 -1 570
box -8 -3 16 105
use FILL  FILL_4424
timestamp 1713400504
transform 1 0 2632 0 -1 570
box -8 -3 16 105
use FILL  FILL_4425
timestamp 1713400504
transform 1 0 2624 0 -1 570
box -8 -3 16 105
use FILL  FILL_4426
timestamp 1713400504
transform 1 0 2616 0 -1 570
box -8 -3 16 105
use FILL  FILL_4427
timestamp 1713400504
transform 1 0 2416 0 -1 570
box -8 -3 16 105
use FILL  FILL_4428
timestamp 1713400504
transform 1 0 2408 0 -1 570
box -8 -3 16 105
use FILL  FILL_4429
timestamp 1713400504
transform 1 0 2304 0 -1 570
box -8 -3 16 105
use FILL  FILL_4430
timestamp 1713400504
transform 1 0 2296 0 -1 570
box -8 -3 16 105
use FILL  FILL_4431
timestamp 1713400504
transform 1 0 2288 0 -1 570
box -8 -3 16 105
use FILL  FILL_4432
timestamp 1713400504
transform 1 0 2280 0 -1 570
box -8 -3 16 105
use FILL  FILL_4433
timestamp 1713400504
transform 1 0 2240 0 -1 570
box -8 -3 16 105
use FILL  FILL_4434
timestamp 1713400504
transform 1 0 2232 0 -1 570
box -8 -3 16 105
use FILL  FILL_4435
timestamp 1713400504
transform 1 0 2224 0 -1 570
box -8 -3 16 105
use FILL  FILL_4436
timestamp 1713400504
transform 1 0 2216 0 -1 570
box -8 -3 16 105
use FILL  FILL_4437
timestamp 1713400504
transform 1 0 2208 0 -1 570
box -8 -3 16 105
use FILL  FILL_4438
timestamp 1713400504
transform 1 0 2200 0 -1 570
box -8 -3 16 105
use FILL  FILL_4439
timestamp 1713400504
transform 1 0 2192 0 -1 570
box -8 -3 16 105
use FILL  FILL_4440
timestamp 1713400504
transform 1 0 2152 0 -1 570
box -8 -3 16 105
use FILL  FILL_4441
timestamp 1713400504
transform 1 0 2144 0 -1 570
box -8 -3 16 105
use FILL  FILL_4442
timestamp 1713400504
transform 1 0 2136 0 -1 570
box -8 -3 16 105
use FILL  FILL_4443
timestamp 1713400504
transform 1 0 2128 0 -1 570
box -8 -3 16 105
use FILL  FILL_4444
timestamp 1713400504
transform 1 0 2120 0 -1 570
box -8 -3 16 105
use FILL  FILL_4445
timestamp 1713400504
transform 1 0 2112 0 -1 570
box -8 -3 16 105
use FILL  FILL_4446
timestamp 1713400504
transform 1 0 2072 0 -1 570
box -8 -3 16 105
use FILL  FILL_4447
timestamp 1713400504
transform 1 0 2064 0 -1 570
box -8 -3 16 105
use FILL  FILL_4448
timestamp 1713400504
transform 1 0 2056 0 -1 570
box -8 -3 16 105
use FILL  FILL_4449
timestamp 1713400504
transform 1 0 2048 0 -1 570
box -8 -3 16 105
use FILL  FILL_4450
timestamp 1713400504
transform 1 0 2040 0 -1 570
box -8 -3 16 105
use FILL  FILL_4451
timestamp 1713400504
transform 1 0 2008 0 -1 570
box -8 -3 16 105
use FILL  FILL_4452
timestamp 1713400504
transform 1 0 2000 0 -1 570
box -8 -3 16 105
use FILL  FILL_4453
timestamp 1713400504
transform 1 0 1992 0 -1 570
box -8 -3 16 105
use FILL  FILL_4454
timestamp 1713400504
transform 1 0 1984 0 -1 570
box -8 -3 16 105
use FILL  FILL_4455
timestamp 1713400504
transform 1 0 1976 0 -1 570
box -8 -3 16 105
use FILL  FILL_4456
timestamp 1713400504
transform 1 0 1968 0 -1 570
box -8 -3 16 105
use FILL  FILL_4457
timestamp 1713400504
transform 1 0 1960 0 -1 570
box -8 -3 16 105
use FILL  FILL_4458
timestamp 1713400504
transform 1 0 1920 0 -1 570
box -8 -3 16 105
use FILL  FILL_4459
timestamp 1713400504
transform 1 0 1912 0 -1 570
box -8 -3 16 105
use FILL  FILL_4460
timestamp 1713400504
transform 1 0 1904 0 -1 570
box -8 -3 16 105
use FILL  FILL_4461
timestamp 1713400504
transform 1 0 1896 0 -1 570
box -8 -3 16 105
use FILL  FILL_4462
timestamp 1713400504
transform 1 0 1888 0 -1 570
box -8 -3 16 105
use FILL  FILL_4463
timestamp 1713400504
transform 1 0 1880 0 -1 570
box -8 -3 16 105
use FILL  FILL_4464
timestamp 1713400504
transform 1 0 1872 0 -1 570
box -8 -3 16 105
use FILL  FILL_4465
timestamp 1713400504
transform 1 0 1864 0 -1 570
box -8 -3 16 105
use FILL  FILL_4466
timestamp 1713400504
transform 1 0 1856 0 -1 570
box -8 -3 16 105
use FILL  FILL_4467
timestamp 1713400504
transform 1 0 1848 0 -1 570
box -8 -3 16 105
use FILL  FILL_4468
timestamp 1713400504
transform 1 0 1840 0 -1 570
box -8 -3 16 105
use FILL  FILL_4469
timestamp 1713400504
transform 1 0 1832 0 -1 570
box -8 -3 16 105
use FILL  FILL_4470
timestamp 1713400504
transform 1 0 1824 0 -1 570
box -8 -3 16 105
use FILL  FILL_4471
timestamp 1713400504
transform 1 0 1816 0 -1 570
box -8 -3 16 105
use FILL  FILL_4472
timestamp 1713400504
transform 1 0 1808 0 -1 570
box -8 -3 16 105
use FILL  FILL_4473
timestamp 1713400504
transform 1 0 1800 0 -1 570
box -8 -3 16 105
use FILL  FILL_4474
timestamp 1713400504
transform 1 0 1792 0 -1 570
box -8 -3 16 105
use FILL  FILL_4475
timestamp 1713400504
transform 1 0 1784 0 -1 570
box -8 -3 16 105
use FILL  FILL_4476
timestamp 1713400504
transform 1 0 1776 0 -1 570
box -8 -3 16 105
use FILL  FILL_4477
timestamp 1713400504
transform 1 0 1736 0 -1 570
box -8 -3 16 105
use FILL  FILL_4478
timestamp 1713400504
transform 1 0 1728 0 -1 570
box -8 -3 16 105
use FILL  FILL_4479
timestamp 1713400504
transform 1 0 1720 0 -1 570
box -8 -3 16 105
use FILL  FILL_4480
timestamp 1713400504
transform 1 0 1712 0 -1 570
box -8 -3 16 105
use FILL  FILL_4481
timestamp 1713400504
transform 1 0 1704 0 -1 570
box -8 -3 16 105
use FILL  FILL_4482
timestamp 1713400504
transform 1 0 1696 0 -1 570
box -8 -3 16 105
use FILL  FILL_4483
timestamp 1713400504
transform 1 0 1688 0 -1 570
box -8 -3 16 105
use FILL  FILL_4484
timestamp 1713400504
transform 1 0 1680 0 -1 570
box -8 -3 16 105
use FILL  FILL_4485
timestamp 1713400504
transform 1 0 1672 0 -1 570
box -8 -3 16 105
use FILL  FILL_4486
timestamp 1713400504
transform 1 0 1632 0 -1 570
box -8 -3 16 105
use FILL  FILL_4487
timestamp 1713400504
transform 1 0 1624 0 -1 570
box -8 -3 16 105
use FILL  FILL_4488
timestamp 1713400504
transform 1 0 1616 0 -1 570
box -8 -3 16 105
use FILL  FILL_4489
timestamp 1713400504
transform 1 0 1608 0 -1 570
box -8 -3 16 105
use FILL  FILL_4490
timestamp 1713400504
transform 1 0 1600 0 -1 570
box -8 -3 16 105
use FILL  FILL_4491
timestamp 1713400504
transform 1 0 1592 0 -1 570
box -8 -3 16 105
use FILL  FILL_4492
timestamp 1713400504
transform 1 0 1584 0 -1 570
box -8 -3 16 105
use FILL  FILL_4493
timestamp 1713400504
transform 1 0 1576 0 -1 570
box -8 -3 16 105
use FILL  FILL_4494
timestamp 1713400504
transform 1 0 1568 0 -1 570
box -8 -3 16 105
use FILL  FILL_4495
timestamp 1713400504
transform 1 0 1560 0 -1 570
box -8 -3 16 105
use FILL  FILL_4496
timestamp 1713400504
transform 1 0 1512 0 -1 570
box -8 -3 16 105
use FILL  FILL_4497
timestamp 1713400504
transform 1 0 1504 0 -1 570
box -8 -3 16 105
use FILL  FILL_4498
timestamp 1713400504
transform 1 0 1496 0 -1 570
box -8 -3 16 105
use FILL  FILL_4499
timestamp 1713400504
transform 1 0 1488 0 -1 570
box -8 -3 16 105
use FILL  FILL_4500
timestamp 1713400504
transform 1 0 1480 0 -1 570
box -8 -3 16 105
use FILL  FILL_4501
timestamp 1713400504
transform 1 0 1472 0 -1 570
box -8 -3 16 105
use FILL  FILL_4502
timestamp 1713400504
transform 1 0 1464 0 -1 570
box -8 -3 16 105
use FILL  FILL_4503
timestamp 1713400504
transform 1 0 1440 0 -1 570
box -8 -3 16 105
use FILL  FILL_4504
timestamp 1713400504
transform 1 0 1432 0 -1 570
box -8 -3 16 105
use FILL  FILL_4505
timestamp 1713400504
transform 1 0 1424 0 -1 570
box -8 -3 16 105
use FILL  FILL_4506
timestamp 1713400504
transform 1 0 1416 0 -1 570
box -8 -3 16 105
use FILL  FILL_4507
timestamp 1713400504
transform 1 0 1376 0 -1 570
box -8 -3 16 105
use FILL  FILL_4508
timestamp 1713400504
transform 1 0 1368 0 -1 570
box -8 -3 16 105
use FILL  FILL_4509
timestamp 1713400504
transform 1 0 1360 0 -1 570
box -8 -3 16 105
use FILL  FILL_4510
timestamp 1713400504
transform 1 0 1352 0 -1 570
box -8 -3 16 105
use FILL  FILL_4511
timestamp 1713400504
transform 1 0 1344 0 -1 570
box -8 -3 16 105
use FILL  FILL_4512
timestamp 1713400504
transform 1 0 1336 0 -1 570
box -8 -3 16 105
use FILL  FILL_4513
timestamp 1713400504
transform 1 0 1328 0 -1 570
box -8 -3 16 105
use FILL  FILL_4514
timestamp 1713400504
transform 1 0 1320 0 -1 570
box -8 -3 16 105
use FILL  FILL_4515
timestamp 1713400504
transform 1 0 1272 0 -1 570
box -8 -3 16 105
use FILL  FILL_4516
timestamp 1713400504
transform 1 0 1264 0 -1 570
box -8 -3 16 105
use FILL  FILL_4517
timestamp 1713400504
transform 1 0 1256 0 -1 570
box -8 -3 16 105
use FILL  FILL_4518
timestamp 1713400504
transform 1 0 1248 0 -1 570
box -8 -3 16 105
use FILL  FILL_4519
timestamp 1713400504
transform 1 0 1240 0 -1 570
box -8 -3 16 105
use FILL  FILL_4520
timestamp 1713400504
transform 1 0 1232 0 -1 570
box -8 -3 16 105
use FILL  FILL_4521
timestamp 1713400504
transform 1 0 1224 0 -1 570
box -8 -3 16 105
use FILL  FILL_4522
timestamp 1713400504
transform 1 0 1176 0 -1 570
box -8 -3 16 105
use FILL  FILL_4523
timestamp 1713400504
transform 1 0 1168 0 -1 570
box -8 -3 16 105
use FILL  FILL_4524
timestamp 1713400504
transform 1 0 1160 0 -1 570
box -8 -3 16 105
use FILL  FILL_4525
timestamp 1713400504
transform 1 0 1152 0 -1 570
box -8 -3 16 105
use FILL  FILL_4526
timestamp 1713400504
transform 1 0 1048 0 -1 570
box -8 -3 16 105
use FILL  FILL_4527
timestamp 1713400504
transform 1 0 1040 0 -1 570
box -8 -3 16 105
use FILL  FILL_4528
timestamp 1713400504
transform 1 0 1032 0 -1 570
box -8 -3 16 105
use FILL  FILL_4529
timestamp 1713400504
transform 1 0 1000 0 -1 570
box -8 -3 16 105
use FILL  FILL_4530
timestamp 1713400504
transform 1 0 992 0 -1 570
box -8 -3 16 105
use FILL  FILL_4531
timestamp 1713400504
transform 1 0 984 0 -1 570
box -8 -3 16 105
use FILL  FILL_4532
timestamp 1713400504
transform 1 0 944 0 -1 570
box -8 -3 16 105
use FILL  FILL_4533
timestamp 1713400504
transform 1 0 936 0 -1 570
box -8 -3 16 105
use FILL  FILL_4534
timestamp 1713400504
transform 1 0 928 0 -1 570
box -8 -3 16 105
use FILL  FILL_4535
timestamp 1713400504
transform 1 0 824 0 -1 570
box -8 -3 16 105
use FILL  FILL_4536
timestamp 1713400504
transform 1 0 816 0 -1 570
box -8 -3 16 105
use FILL  FILL_4537
timestamp 1713400504
transform 1 0 808 0 -1 570
box -8 -3 16 105
use FILL  FILL_4538
timestamp 1713400504
transform 1 0 776 0 -1 570
box -8 -3 16 105
use FILL  FILL_4539
timestamp 1713400504
transform 1 0 768 0 -1 570
box -8 -3 16 105
use FILL  FILL_4540
timestamp 1713400504
transform 1 0 760 0 -1 570
box -8 -3 16 105
use FILL  FILL_4541
timestamp 1713400504
transform 1 0 752 0 -1 570
box -8 -3 16 105
use FILL  FILL_4542
timestamp 1713400504
transform 1 0 712 0 -1 570
box -8 -3 16 105
use FILL  FILL_4543
timestamp 1713400504
transform 1 0 704 0 -1 570
box -8 -3 16 105
use FILL  FILL_4544
timestamp 1713400504
transform 1 0 696 0 -1 570
box -8 -3 16 105
use FILL  FILL_4545
timestamp 1713400504
transform 1 0 688 0 -1 570
box -8 -3 16 105
use FILL  FILL_4546
timestamp 1713400504
transform 1 0 680 0 -1 570
box -8 -3 16 105
use FILL  FILL_4547
timestamp 1713400504
transform 1 0 672 0 -1 570
box -8 -3 16 105
use FILL  FILL_4548
timestamp 1713400504
transform 1 0 664 0 -1 570
box -8 -3 16 105
use FILL  FILL_4549
timestamp 1713400504
transform 1 0 624 0 -1 570
box -8 -3 16 105
use FILL  FILL_4550
timestamp 1713400504
transform 1 0 616 0 -1 570
box -8 -3 16 105
use FILL  FILL_4551
timestamp 1713400504
transform 1 0 608 0 -1 570
box -8 -3 16 105
use FILL  FILL_4552
timestamp 1713400504
transform 1 0 600 0 -1 570
box -8 -3 16 105
use FILL  FILL_4553
timestamp 1713400504
transform 1 0 560 0 -1 570
box -8 -3 16 105
use FILL  FILL_4554
timestamp 1713400504
transform 1 0 552 0 -1 570
box -8 -3 16 105
use FILL  FILL_4555
timestamp 1713400504
transform 1 0 544 0 -1 570
box -8 -3 16 105
use FILL  FILL_4556
timestamp 1713400504
transform 1 0 536 0 -1 570
box -8 -3 16 105
use FILL  FILL_4557
timestamp 1713400504
transform 1 0 528 0 -1 570
box -8 -3 16 105
use FILL  FILL_4558
timestamp 1713400504
transform 1 0 504 0 -1 570
box -8 -3 16 105
use FILL  FILL_4559
timestamp 1713400504
transform 1 0 496 0 -1 570
box -8 -3 16 105
use FILL  FILL_4560
timestamp 1713400504
transform 1 0 488 0 -1 570
box -8 -3 16 105
use FILL  FILL_4561
timestamp 1713400504
transform 1 0 448 0 -1 570
box -8 -3 16 105
use FILL  FILL_4562
timestamp 1713400504
transform 1 0 440 0 -1 570
box -8 -3 16 105
use FILL  FILL_4563
timestamp 1713400504
transform 1 0 432 0 -1 570
box -8 -3 16 105
use FILL  FILL_4564
timestamp 1713400504
transform 1 0 424 0 -1 570
box -8 -3 16 105
use FILL  FILL_4565
timestamp 1713400504
transform 1 0 416 0 -1 570
box -8 -3 16 105
use FILL  FILL_4566
timestamp 1713400504
transform 1 0 408 0 -1 570
box -8 -3 16 105
use FILL  FILL_4567
timestamp 1713400504
transform 1 0 400 0 -1 570
box -8 -3 16 105
use FILL  FILL_4568
timestamp 1713400504
transform 1 0 360 0 -1 570
box -8 -3 16 105
use FILL  FILL_4569
timestamp 1713400504
transform 1 0 352 0 -1 570
box -8 -3 16 105
use FILL  FILL_4570
timestamp 1713400504
transform 1 0 344 0 -1 570
box -8 -3 16 105
use FILL  FILL_4571
timestamp 1713400504
transform 1 0 336 0 -1 570
box -8 -3 16 105
use FILL  FILL_4572
timestamp 1713400504
transform 1 0 328 0 -1 570
box -8 -3 16 105
use FILL  FILL_4573
timestamp 1713400504
transform 1 0 288 0 -1 570
box -8 -3 16 105
use FILL  FILL_4574
timestamp 1713400504
transform 1 0 280 0 -1 570
box -8 -3 16 105
use FILL  FILL_4575
timestamp 1713400504
transform 1 0 272 0 -1 570
box -8 -3 16 105
use FILL  FILL_4576
timestamp 1713400504
transform 1 0 264 0 -1 570
box -8 -3 16 105
use FILL  FILL_4577
timestamp 1713400504
transform 1 0 256 0 -1 570
box -8 -3 16 105
use FILL  FILL_4578
timestamp 1713400504
transform 1 0 216 0 -1 570
box -8 -3 16 105
use FILL  FILL_4579
timestamp 1713400504
transform 1 0 208 0 -1 570
box -8 -3 16 105
use FILL  FILL_4580
timestamp 1713400504
transform 1 0 200 0 -1 570
box -8 -3 16 105
use FILL  FILL_4581
timestamp 1713400504
transform 1 0 192 0 -1 570
box -8 -3 16 105
use FILL  FILL_4582
timestamp 1713400504
transform 1 0 184 0 -1 570
box -8 -3 16 105
use FILL  FILL_4583
timestamp 1713400504
transform 1 0 176 0 -1 570
box -8 -3 16 105
use FILL  FILL_4584
timestamp 1713400504
transform 1 0 72 0 -1 570
box -8 -3 16 105
use FILL  FILL_4585
timestamp 1713400504
transform 1 0 3008 0 1 370
box -8 -3 16 105
use FILL  FILL_4586
timestamp 1713400504
transform 1 0 3000 0 1 370
box -8 -3 16 105
use FILL  FILL_4587
timestamp 1713400504
transform 1 0 2992 0 1 370
box -8 -3 16 105
use FILL  FILL_4588
timestamp 1713400504
transform 1 0 2984 0 1 370
box -8 -3 16 105
use FILL  FILL_4589
timestamp 1713400504
transform 1 0 2976 0 1 370
box -8 -3 16 105
use FILL  FILL_4590
timestamp 1713400504
transform 1 0 2968 0 1 370
box -8 -3 16 105
use FILL  FILL_4591
timestamp 1713400504
transform 1 0 2960 0 1 370
box -8 -3 16 105
use FILL  FILL_4592
timestamp 1713400504
transform 1 0 2952 0 1 370
box -8 -3 16 105
use FILL  FILL_4593
timestamp 1713400504
transform 1 0 2944 0 1 370
box -8 -3 16 105
use FILL  FILL_4594
timestamp 1713400504
transform 1 0 2936 0 1 370
box -8 -3 16 105
use FILL  FILL_4595
timestamp 1713400504
transform 1 0 2896 0 1 370
box -8 -3 16 105
use FILL  FILL_4596
timestamp 1713400504
transform 1 0 2888 0 1 370
box -8 -3 16 105
use FILL  FILL_4597
timestamp 1713400504
transform 1 0 2880 0 1 370
box -8 -3 16 105
use FILL  FILL_4598
timestamp 1713400504
transform 1 0 2872 0 1 370
box -8 -3 16 105
use FILL  FILL_4599
timestamp 1713400504
transform 1 0 2864 0 1 370
box -8 -3 16 105
use FILL  FILL_4600
timestamp 1713400504
transform 1 0 2856 0 1 370
box -8 -3 16 105
use FILL  FILL_4601
timestamp 1713400504
transform 1 0 2848 0 1 370
box -8 -3 16 105
use FILL  FILL_4602
timestamp 1713400504
transform 1 0 2840 0 1 370
box -8 -3 16 105
use FILL  FILL_4603
timestamp 1713400504
transform 1 0 2832 0 1 370
box -8 -3 16 105
use FILL  FILL_4604
timestamp 1713400504
transform 1 0 2824 0 1 370
box -8 -3 16 105
use FILL  FILL_4605
timestamp 1713400504
transform 1 0 2784 0 1 370
box -8 -3 16 105
use FILL  FILL_4606
timestamp 1713400504
transform 1 0 2776 0 1 370
box -8 -3 16 105
use FILL  FILL_4607
timestamp 1713400504
transform 1 0 2768 0 1 370
box -8 -3 16 105
use FILL  FILL_4608
timestamp 1713400504
transform 1 0 2760 0 1 370
box -8 -3 16 105
use FILL  FILL_4609
timestamp 1713400504
transform 1 0 2752 0 1 370
box -8 -3 16 105
use FILL  FILL_4610
timestamp 1713400504
transform 1 0 2744 0 1 370
box -8 -3 16 105
use FILL  FILL_4611
timestamp 1713400504
transform 1 0 2736 0 1 370
box -8 -3 16 105
use FILL  FILL_4612
timestamp 1713400504
transform 1 0 2728 0 1 370
box -8 -3 16 105
use FILL  FILL_4613
timestamp 1713400504
transform 1 0 2680 0 1 370
box -8 -3 16 105
use FILL  FILL_4614
timestamp 1713400504
transform 1 0 2672 0 1 370
box -8 -3 16 105
use FILL  FILL_4615
timestamp 1713400504
transform 1 0 2664 0 1 370
box -8 -3 16 105
use FILL  FILL_4616
timestamp 1713400504
transform 1 0 2656 0 1 370
box -8 -3 16 105
use FILL  FILL_4617
timestamp 1713400504
transform 1 0 2648 0 1 370
box -8 -3 16 105
use FILL  FILL_4618
timestamp 1713400504
transform 1 0 2640 0 1 370
box -8 -3 16 105
use FILL  FILL_4619
timestamp 1713400504
transform 1 0 2632 0 1 370
box -8 -3 16 105
use FILL  FILL_4620
timestamp 1713400504
transform 1 0 2624 0 1 370
box -8 -3 16 105
use FILL  FILL_4621
timestamp 1713400504
transform 1 0 2592 0 1 370
box -8 -3 16 105
use FILL  FILL_4622
timestamp 1713400504
transform 1 0 2584 0 1 370
box -8 -3 16 105
use FILL  FILL_4623
timestamp 1713400504
transform 1 0 2576 0 1 370
box -8 -3 16 105
use FILL  FILL_4624
timestamp 1713400504
transform 1 0 2568 0 1 370
box -8 -3 16 105
use FILL  FILL_4625
timestamp 1713400504
transform 1 0 2464 0 1 370
box -8 -3 16 105
use FILL  FILL_4626
timestamp 1713400504
transform 1 0 2456 0 1 370
box -8 -3 16 105
use FILL  FILL_4627
timestamp 1713400504
transform 1 0 2448 0 1 370
box -8 -3 16 105
use FILL  FILL_4628
timestamp 1713400504
transform 1 0 2440 0 1 370
box -8 -3 16 105
use FILL  FILL_4629
timestamp 1713400504
transform 1 0 2432 0 1 370
box -8 -3 16 105
use FILL  FILL_4630
timestamp 1713400504
transform 1 0 2408 0 1 370
box -8 -3 16 105
use FILL  FILL_4631
timestamp 1713400504
transform 1 0 2384 0 1 370
box -8 -3 16 105
use FILL  FILL_4632
timestamp 1713400504
transform 1 0 2376 0 1 370
box -8 -3 16 105
use FILL  FILL_4633
timestamp 1713400504
transform 1 0 2368 0 1 370
box -8 -3 16 105
use FILL  FILL_4634
timestamp 1713400504
transform 1 0 2360 0 1 370
box -8 -3 16 105
use FILL  FILL_4635
timestamp 1713400504
transform 1 0 2352 0 1 370
box -8 -3 16 105
use FILL  FILL_4636
timestamp 1713400504
transform 1 0 2344 0 1 370
box -8 -3 16 105
use FILL  FILL_4637
timestamp 1713400504
transform 1 0 2336 0 1 370
box -8 -3 16 105
use FILL  FILL_4638
timestamp 1713400504
transform 1 0 2328 0 1 370
box -8 -3 16 105
use FILL  FILL_4639
timestamp 1713400504
transform 1 0 2320 0 1 370
box -8 -3 16 105
use FILL  FILL_4640
timestamp 1713400504
transform 1 0 2280 0 1 370
box -8 -3 16 105
use FILL  FILL_4641
timestamp 1713400504
transform 1 0 2272 0 1 370
box -8 -3 16 105
use FILL  FILL_4642
timestamp 1713400504
transform 1 0 2264 0 1 370
box -8 -3 16 105
use FILL  FILL_4643
timestamp 1713400504
transform 1 0 2256 0 1 370
box -8 -3 16 105
use FILL  FILL_4644
timestamp 1713400504
transform 1 0 2248 0 1 370
box -8 -3 16 105
use FILL  FILL_4645
timestamp 1713400504
transform 1 0 2240 0 1 370
box -8 -3 16 105
use FILL  FILL_4646
timestamp 1713400504
transform 1 0 2232 0 1 370
box -8 -3 16 105
use FILL  FILL_4647
timestamp 1713400504
transform 1 0 2208 0 1 370
box -8 -3 16 105
use FILL  FILL_4648
timestamp 1713400504
transform 1 0 2200 0 1 370
box -8 -3 16 105
use FILL  FILL_4649
timestamp 1713400504
transform 1 0 2192 0 1 370
box -8 -3 16 105
use FILL  FILL_4650
timestamp 1713400504
transform 1 0 2184 0 1 370
box -8 -3 16 105
use FILL  FILL_4651
timestamp 1713400504
transform 1 0 2144 0 1 370
box -8 -3 16 105
use FILL  FILL_4652
timestamp 1713400504
transform 1 0 2136 0 1 370
box -8 -3 16 105
use FILL  FILL_4653
timestamp 1713400504
transform 1 0 2128 0 1 370
box -8 -3 16 105
use FILL  FILL_4654
timestamp 1713400504
transform 1 0 2120 0 1 370
box -8 -3 16 105
use FILL  FILL_4655
timestamp 1713400504
transform 1 0 2112 0 1 370
box -8 -3 16 105
use FILL  FILL_4656
timestamp 1713400504
transform 1 0 2104 0 1 370
box -8 -3 16 105
use FILL  FILL_4657
timestamp 1713400504
transform 1 0 2072 0 1 370
box -8 -3 16 105
use FILL  FILL_4658
timestamp 1713400504
transform 1 0 2064 0 1 370
box -8 -3 16 105
use FILL  FILL_4659
timestamp 1713400504
transform 1 0 2056 0 1 370
box -8 -3 16 105
use FILL  FILL_4660
timestamp 1713400504
transform 1 0 2048 0 1 370
box -8 -3 16 105
use FILL  FILL_4661
timestamp 1713400504
transform 1 0 2040 0 1 370
box -8 -3 16 105
use FILL  FILL_4662
timestamp 1713400504
transform 1 0 2032 0 1 370
box -8 -3 16 105
use FILL  FILL_4663
timestamp 1713400504
transform 1 0 1960 0 1 370
box -8 -3 16 105
use FILL  FILL_4664
timestamp 1713400504
transform 1 0 1952 0 1 370
box -8 -3 16 105
use FILL  FILL_4665
timestamp 1713400504
transform 1 0 1944 0 1 370
box -8 -3 16 105
use FILL  FILL_4666
timestamp 1713400504
transform 1 0 1936 0 1 370
box -8 -3 16 105
use FILL  FILL_4667
timestamp 1713400504
transform 1 0 1832 0 1 370
box -8 -3 16 105
use FILL  FILL_4668
timestamp 1713400504
transform 1 0 1824 0 1 370
box -8 -3 16 105
use FILL  FILL_4669
timestamp 1713400504
transform 1 0 1816 0 1 370
box -8 -3 16 105
use FILL  FILL_4670
timestamp 1713400504
transform 1 0 1808 0 1 370
box -8 -3 16 105
use FILL  FILL_4671
timestamp 1713400504
transform 1 0 1768 0 1 370
box -8 -3 16 105
use FILL  FILL_4672
timestamp 1713400504
transform 1 0 1760 0 1 370
box -8 -3 16 105
use FILL  FILL_4673
timestamp 1713400504
transform 1 0 1752 0 1 370
box -8 -3 16 105
use FILL  FILL_4674
timestamp 1713400504
transform 1 0 1744 0 1 370
box -8 -3 16 105
use FILL  FILL_4675
timestamp 1713400504
transform 1 0 1736 0 1 370
box -8 -3 16 105
use FILL  FILL_4676
timestamp 1713400504
transform 1 0 1632 0 1 370
box -8 -3 16 105
use FILL  FILL_4677
timestamp 1713400504
transform 1 0 1624 0 1 370
box -8 -3 16 105
use FILL  FILL_4678
timestamp 1713400504
transform 1 0 1616 0 1 370
box -8 -3 16 105
use FILL  FILL_4679
timestamp 1713400504
transform 1 0 1608 0 1 370
box -8 -3 16 105
use FILL  FILL_4680
timestamp 1713400504
transform 1 0 1600 0 1 370
box -8 -3 16 105
use FILL  FILL_4681
timestamp 1713400504
transform 1 0 1592 0 1 370
box -8 -3 16 105
use FILL  FILL_4682
timestamp 1713400504
transform 1 0 1584 0 1 370
box -8 -3 16 105
use FILL  FILL_4683
timestamp 1713400504
transform 1 0 1560 0 1 370
box -8 -3 16 105
use FILL  FILL_4684
timestamp 1713400504
transform 1 0 1552 0 1 370
box -8 -3 16 105
use FILL  FILL_4685
timestamp 1713400504
transform 1 0 1544 0 1 370
box -8 -3 16 105
use FILL  FILL_4686
timestamp 1713400504
transform 1 0 1536 0 1 370
box -8 -3 16 105
use FILL  FILL_4687
timestamp 1713400504
transform 1 0 1528 0 1 370
box -8 -3 16 105
use FILL  FILL_4688
timestamp 1713400504
transform 1 0 1520 0 1 370
box -8 -3 16 105
use FILL  FILL_4689
timestamp 1713400504
transform 1 0 1512 0 1 370
box -8 -3 16 105
use FILL  FILL_4690
timestamp 1713400504
transform 1 0 1504 0 1 370
box -8 -3 16 105
use FILL  FILL_4691
timestamp 1713400504
transform 1 0 1496 0 1 370
box -8 -3 16 105
use FILL  FILL_4692
timestamp 1713400504
transform 1 0 1488 0 1 370
box -8 -3 16 105
use FILL  FILL_4693
timestamp 1713400504
transform 1 0 1480 0 1 370
box -8 -3 16 105
use FILL  FILL_4694
timestamp 1713400504
transform 1 0 1472 0 1 370
box -8 -3 16 105
use FILL  FILL_4695
timestamp 1713400504
transform 1 0 1432 0 1 370
box -8 -3 16 105
use FILL  FILL_4696
timestamp 1713400504
transform 1 0 1424 0 1 370
box -8 -3 16 105
use FILL  FILL_4697
timestamp 1713400504
transform 1 0 1416 0 1 370
box -8 -3 16 105
use FILL  FILL_4698
timestamp 1713400504
transform 1 0 1408 0 1 370
box -8 -3 16 105
use FILL  FILL_4699
timestamp 1713400504
transform 1 0 1400 0 1 370
box -8 -3 16 105
use FILL  FILL_4700
timestamp 1713400504
transform 1 0 1392 0 1 370
box -8 -3 16 105
use FILL  FILL_4701
timestamp 1713400504
transform 1 0 1384 0 1 370
box -8 -3 16 105
use FILL  FILL_4702
timestamp 1713400504
transform 1 0 1376 0 1 370
box -8 -3 16 105
use FILL  FILL_4703
timestamp 1713400504
transform 1 0 1368 0 1 370
box -8 -3 16 105
use FILL  FILL_4704
timestamp 1713400504
transform 1 0 1328 0 1 370
box -8 -3 16 105
use FILL  FILL_4705
timestamp 1713400504
transform 1 0 1320 0 1 370
box -8 -3 16 105
use FILL  FILL_4706
timestamp 1713400504
transform 1 0 1312 0 1 370
box -8 -3 16 105
use FILL  FILL_4707
timestamp 1713400504
transform 1 0 1304 0 1 370
box -8 -3 16 105
use FILL  FILL_4708
timestamp 1713400504
transform 1 0 1296 0 1 370
box -8 -3 16 105
use FILL  FILL_4709
timestamp 1713400504
transform 1 0 1288 0 1 370
box -8 -3 16 105
use FILL  FILL_4710
timestamp 1713400504
transform 1 0 1280 0 1 370
box -8 -3 16 105
use FILL  FILL_4711
timestamp 1713400504
transform 1 0 1272 0 1 370
box -8 -3 16 105
use FILL  FILL_4712
timestamp 1713400504
transform 1 0 1264 0 1 370
box -8 -3 16 105
use FILL  FILL_4713
timestamp 1713400504
transform 1 0 1216 0 1 370
box -8 -3 16 105
use FILL  FILL_4714
timestamp 1713400504
transform 1 0 1208 0 1 370
box -8 -3 16 105
use FILL  FILL_4715
timestamp 1713400504
transform 1 0 1200 0 1 370
box -8 -3 16 105
use FILL  FILL_4716
timestamp 1713400504
transform 1 0 1192 0 1 370
box -8 -3 16 105
use FILL  FILL_4717
timestamp 1713400504
transform 1 0 1184 0 1 370
box -8 -3 16 105
use FILL  FILL_4718
timestamp 1713400504
transform 1 0 1176 0 1 370
box -8 -3 16 105
use FILL  FILL_4719
timestamp 1713400504
transform 1 0 1168 0 1 370
box -8 -3 16 105
use FILL  FILL_4720
timestamp 1713400504
transform 1 0 1160 0 1 370
box -8 -3 16 105
use FILL  FILL_4721
timestamp 1713400504
transform 1 0 1152 0 1 370
box -8 -3 16 105
use FILL  FILL_4722
timestamp 1713400504
transform 1 0 1144 0 1 370
box -8 -3 16 105
use FILL  FILL_4723
timestamp 1713400504
transform 1 0 1112 0 1 370
box -8 -3 16 105
use FILL  FILL_4724
timestamp 1713400504
transform 1 0 1104 0 1 370
box -8 -3 16 105
use FILL  FILL_4725
timestamp 1713400504
transform 1 0 1096 0 1 370
box -8 -3 16 105
use FILL  FILL_4726
timestamp 1713400504
transform 1 0 1088 0 1 370
box -8 -3 16 105
use FILL  FILL_4727
timestamp 1713400504
transform 1 0 1080 0 1 370
box -8 -3 16 105
use FILL  FILL_4728
timestamp 1713400504
transform 1 0 1072 0 1 370
box -8 -3 16 105
use FILL  FILL_4729
timestamp 1713400504
transform 1 0 1064 0 1 370
box -8 -3 16 105
use FILL  FILL_4730
timestamp 1713400504
transform 1 0 1024 0 1 370
box -8 -3 16 105
use FILL  FILL_4731
timestamp 1713400504
transform 1 0 1016 0 1 370
box -8 -3 16 105
use FILL  FILL_4732
timestamp 1713400504
transform 1 0 1008 0 1 370
box -8 -3 16 105
use FILL  FILL_4733
timestamp 1713400504
transform 1 0 1000 0 1 370
box -8 -3 16 105
use FILL  FILL_4734
timestamp 1713400504
transform 1 0 992 0 1 370
box -8 -3 16 105
use FILL  FILL_4735
timestamp 1713400504
transform 1 0 984 0 1 370
box -8 -3 16 105
use FILL  FILL_4736
timestamp 1713400504
transform 1 0 976 0 1 370
box -8 -3 16 105
use FILL  FILL_4737
timestamp 1713400504
transform 1 0 952 0 1 370
box -8 -3 16 105
use FILL  FILL_4738
timestamp 1713400504
transform 1 0 944 0 1 370
box -8 -3 16 105
use FILL  FILL_4739
timestamp 1713400504
transform 1 0 936 0 1 370
box -8 -3 16 105
use FILL  FILL_4740
timestamp 1713400504
transform 1 0 928 0 1 370
box -8 -3 16 105
use FILL  FILL_4741
timestamp 1713400504
transform 1 0 920 0 1 370
box -8 -3 16 105
use FILL  FILL_4742
timestamp 1713400504
transform 1 0 912 0 1 370
box -8 -3 16 105
use FILL  FILL_4743
timestamp 1713400504
transform 1 0 880 0 1 370
box -8 -3 16 105
use FILL  FILL_4744
timestamp 1713400504
transform 1 0 872 0 1 370
box -8 -3 16 105
use FILL  FILL_4745
timestamp 1713400504
transform 1 0 864 0 1 370
box -8 -3 16 105
use FILL  FILL_4746
timestamp 1713400504
transform 1 0 856 0 1 370
box -8 -3 16 105
use FILL  FILL_4747
timestamp 1713400504
transform 1 0 832 0 1 370
box -8 -3 16 105
use FILL  FILL_4748
timestamp 1713400504
transform 1 0 824 0 1 370
box -8 -3 16 105
use FILL  FILL_4749
timestamp 1713400504
transform 1 0 816 0 1 370
box -8 -3 16 105
use FILL  FILL_4750
timestamp 1713400504
transform 1 0 808 0 1 370
box -8 -3 16 105
use FILL  FILL_4751
timestamp 1713400504
transform 1 0 800 0 1 370
box -8 -3 16 105
use FILL  FILL_4752
timestamp 1713400504
transform 1 0 760 0 1 370
box -8 -3 16 105
use FILL  FILL_4753
timestamp 1713400504
transform 1 0 752 0 1 370
box -8 -3 16 105
use FILL  FILL_4754
timestamp 1713400504
transform 1 0 744 0 1 370
box -8 -3 16 105
use FILL  FILL_4755
timestamp 1713400504
transform 1 0 736 0 1 370
box -8 -3 16 105
use FILL  FILL_4756
timestamp 1713400504
transform 1 0 728 0 1 370
box -8 -3 16 105
use FILL  FILL_4757
timestamp 1713400504
transform 1 0 720 0 1 370
box -8 -3 16 105
use FILL  FILL_4758
timestamp 1713400504
transform 1 0 712 0 1 370
box -8 -3 16 105
use FILL  FILL_4759
timestamp 1713400504
transform 1 0 704 0 1 370
box -8 -3 16 105
use FILL  FILL_4760
timestamp 1713400504
transform 1 0 664 0 1 370
box -8 -3 16 105
use FILL  FILL_4761
timestamp 1713400504
transform 1 0 656 0 1 370
box -8 -3 16 105
use FILL  FILL_4762
timestamp 1713400504
transform 1 0 648 0 1 370
box -8 -3 16 105
use FILL  FILL_4763
timestamp 1713400504
transform 1 0 640 0 1 370
box -8 -3 16 105
use FILL  FILL_4764
timestamp 1713400504
transform 1 0 632 0 1 370
box -8 -3 16 105
use FILL  FILL_4765
timestamp 1713400504
transform 1 0 624 0 1 370
box -8 -3 16 105
use FILL  FILL_4766
timestamp 1713400504
transform 1 0 592 0 1 370
box -8 -3 16 105
use FILL  FILL_4767
timestamp 1713400504
transform 1 0 584 0 1 370
box -8 -3 16 105
use FILL  FILL_4768
timestamp 1713400504
transform 1 0 576 0 1 370
box -8 -3 16 105
use FILL  FILL_4769
timestamp 1713400504
transform 1 0 568 0 1 370
box -8 -3 16 105
use FILL  FILL_4770
timestamp 1713400504
transform 1 0 560 0 1 370
box -8 -3 16 105
use FILL  FILL_4771
timestamp 1713400504
transform 1 0 520 0 1 370
box -8 -3 16 105
use FILL  FILL_4772
timestamp 1713400504
transform 1 0 512 0 1 370
box -8 -3 16 105
use FILL  FILL_4773
timestamp 1713400504
transform 1 0 504 0 1 370
box -8 -3 16 105
use FILL  FILL_4774
timestamp 1713400504
transform 1 0 496 0 1 370
box -8 -3 16 105
use FILL  FILL_4775
timestamp 1713400504
transform 1 0 392 0 1 370
box -8 -3 16 105
use FILL  FILL_4776
timestamp 1713400504
transform 1 0 384 0 1 370
box -8 -3 16 105
use FILL  FILL_4777
timestamp 1713400504
transform 1 0 376 0 1 370
box -8 -3 16 105
use FILL  FILL_4778
timestamp 1713400504
transform 1 0 368 0 1 370
box -8 -3 16 105
use FILL  FILL_4779
timestamp 1713400504
transform 1 0 360 0 1 370
box -8 -3 16 105
use FILL  FILL_4780
timestamp 1713400504
transform 1 0 352 0 1 370
box -8 -3 16 105
use FILL  FILL_4781
timestamp 1713400504
transform 1 0 312 0 1 370
box -8 -3 16 105
use FILL  FILL_4782
timestamp 1713400504
transform 1 0 304 0 1 370
box -8 -3 16 105
use FILL  FILL_4783
timestamp 1713400504
transform 1 0 296 0 1 370
box -8 -3 16 105
use FILL  FILL_4784
timestamp 1713400504
transform 1 0 288 0 1 370
box -8 -3 16 105
use FILL  FILL_4785
timestamp 1713400504
transform 1 0 280 0 1 370
box -8 -3 16 105
use FILL  FILL_4786
timestamp 1713400504
transform 1 0 272 0 1 370
box -8 -3 16 105
use FILL  FILL_4787
timestamp 1713400504
transform 1 0 240 0 1 370
box -8 -3 16 105
use FILL  FILL_4788
timestamp 1713400504
transform 1 0 232 0 1 370
box -8 -3 16 105
use FILL  FILL_4789
timestamp 1713400504
transform 1 0 224 0 1 370
box -8 -3 16 105
use FILL  FILL_4790
timestamp 1713400504
transform 1 0 216 0 1 370
box -8 -3 16 105
use FILL  FILL_4791
timestamp 1713400504
transform 1 0 208 0 1 370
box -8 -3 16 105
use FILL  FILL_4792
timestamp 1713400504
transform 1 0 200 0 1 370
box -8 -3 16 105
use FILL  FILL_4793
timestamp 1713400504
transform 1 0 192 0 1 370
box -8 -3 16 105
use FILL  FILL_4794
timestamp 1713400504
transform 1 0 144 0 1 370
box -8 -3 16 105
use FILL  FILL_4795
timestamp 1713400504
transform 1 0 136 0 1 370
box -8 -3 16 105
use FILL  FILL_4796
timestamp 1713400504
transform 1 0 128 0 1 370
box -8 -3 16 105
use FILL  FILL_4797
timestamp 1713400504
transform 1 0 120 0 1 370
box -8 -3 16 105
use FILL  FILL_4798
timestamp 1713400504
transform 1 0 112 0 1 370
box -8 -3 16 105
use FILL  FILL_4799
timestamp 1713400504
transform 1 0 104 0 1 370
box -8 -3 16 105
use FILL  FILL_4800
timestamp 1713400504
transform 1 0 96 0 1 370
box -8 -3 16 105
use FILL  FILL_4801
timestamp 1713400504
transform 1 0 72 0 1 370
box -8 -3 16 105
use FILL  FILL_4802
timestamp 1713400504
transform 1 0 3008 0 -1 370
box -8 -3 16 105
use FILL  FILL_4803
timestamp 1713400504
transform 1 0 3000 0 -1 370
box -8 -3 16 105
use FILL  FILL_4804
timestamp 1713400504
transform 1 0 2992 0 -1 370
box -8 -3 16 105
use FILL  FILL_4805
timestamp 1713400504
transform 1 0 2952 0 -1 370
box -8 -3 16 105
use FILL  FILL_4806
timestamp 1713400504
transform 1 0 2944 0 -1 370
box -8 -3 16 105
use FILL  FILL_4807
timestamp 1713400504
transform 1 0 2936 0 -1 370
box -8 -3 16 105
use FILL  FILL_4808
timestamp 1713400504
transform 1 0 2928 0 -1 370
box -8 -3 16 105
use FILL  FILL_4809
timestamp 1713400504
transform 1 0 2920 0 -1 370
box -8 -3 16 105
use FILL  FILL_4810
timestamp 1713400504
transform 1 0 2912 0 -1 370
box -8 -3 16 105
use FILL  FILL_4811
timestamp 1713400504
transform 1 0 2864 0 -1 370
box -8 -3 16 105
use FILL  FILL_4812
timestamp 1713400504
transform 1 0 2856 0 -1 370
box -8 -3 16 105
use FILL  FILL_4813
timestamp 1713400504
transform 1 0 2848 0 -1 370
box -8 -3 16 105
use FILL  FILL_4814
timestamp 1713400504
transform 1 0 2840 0 -1 370
box -8 -3 16 105
use FILL  FILL_4815
timestamp 1713400504
transform 1 0 2832 0 -1 370
box -8 -3 16 105
use FILL  FILL_4816
timestamp 1713400504
transform 1 0 2824 0 -1 370
box -8 -3 16 105
use FILL  FILL_4817
timestamp 1713400504
transform 1 0 2816 0 -1 370
box -8 -3 16 105
use FILL  FILL_4818
timestamp 1713400504
transform 1 0 2768 0 -1 370
box -8 -3 16 105
use FILL  FILL_4819
timestamp 1713400504
transform 1 0 2760 0 -1 370
box -8 -3 16 105
use FILL  FILL_4820
timestamp 1713400504
transform 1 0 2752 0 -1 370
box -8 -3 16 105
use FILL  FILL_4821
timestamp 1713400504
transform 1 0 2744 0 -1 370
box -8 -3 16 105
use FILL  FILL_4822
timestamp 1713400504
transform 1 0 2736 0 -1 370
box -8 -3 16 105
use FILL  FILL_4823
timestamp 1713400504
transform 1 0 2728 0 -1 370
box -8 -3 16 105
use FILL  FILL_4824
timestamp 1713400504
transform 1 0 2720 0 -1 370
box -8 -3 16 105
use FILL  FILL_4825
timestamp 1713400504
transform 1 0 2672 0 -1 370
box -8 -3 16 105
use FILL  FILL_4826
timestamp 1713400504
transform 1 0 2664 0 -1 370
box -8 -3 16 105
use FILL  FILL_4827
timestamp 1713400504
transform 1 0 2656 0 -1 370
box -8 -3 16 105
use FILL  FILL_4828
timestamp 1713400504
transform 1 0 2456 0 -1 370
box -8 -3 16 105
use FILL  FILL_4829
timestamp 1713400504
transform 1 0 2448 0 -1 370
box -8 -3 16 105
use FILL  FILL_4830
timestamp 1713400504
transform 1 0 2416 0 -1 370
box -8 -3 16 105
use FILL  FILL_4831
timestamp 1713400504
transform 1 0 2408 0 -1 370
box -8 -3 16 105
use FILL  FILL_4832
timestamp 1713400504
transform 1 0 2400 0 -1 370
box -8 -3 16 105
use FILL  FILL_4833
timestamp 1713400504
transform 1 0 2336 0 -1 370
box -8 -3 16 105
use FILL  FILL_4834
timestamp 1713400504
transform 1 0 2328 0 -1 370
box -8 -3 16 105
use FILL  FILL_4835
timestamp 1713400504
transform 1 0 2320 0 -1 370
box -8 -3 16 105
use FILL  FILL_4836
timestamp 1713400504
transform 1 0 2288 0 -1 370
box -8 -3 16 105
use FILL  FILL_4837
timestamp 1713400504
transform 1 0 2280 0 -1 370
box -8 -3 16 105
use FILL  FILL_4838
timestamp 1713400504
transform 1 0 2272 0 -1 370
box -8 -3 16 105
use FILL  FILL_4839
timestamp 1713400504
transform 1 0 2264 0 -1 370
box -8 -3 16 105
use FILL  FILL_4840
timestamp 1713400504
transform 1 0 2256 0 -1 370
box -8 -3 16 105
use FILL  FILL_4841
timestamp 1713400504
transform 1 0 2232 0 -1 370
box -8 -3 16 105
use FILL  FILL_4842
timestamp 1713400504
transform 1 0 2224 0 -1 370
box -8 -3 16 105
use FILL  FILL_4843
timestamp 1713400504
transform 1 0 2216 0 -1 370
box -8 -3 16 105
use FILL  FILL_4844
timestamp 1713400504
transform 1 0 2184 0 -1 370
box -8 -3 16 105
use FILL  FILL_4845
timestamp 1713400504
transform 1 0 2176 0 -1 370
box -8 -3 16 105
use FILL  FILL_4846
timestamp 1713400504
transform 1 0 2168 0 -1 370
box -8 -3 16 105
use FILL  FILL_4847
timestamp 1713400504
transform 1 0 2160 0 -1 370
box -8 -3 16 105
use FILL  FILL_4848
timestamp 1713400504
transform 1 0 2152 0 -1 370
box -8 -3 16 105
use FILL  FILL_4849
timestamp 1713400504
transform 1 0 2144 0 -1 370
box -8 -3 16 105
use FILL  FILL_4850
timestamp 1713400504
transform 1 0 2136 0 -1 370
box -8 -3 16 105
use FILL  FILL_4851
timestamp 1713400504
transform 1 0 2096 0 -1 370
box -8 -3 16 105
use FILL  FILL_4852
timestamp 1713400504
transform 1 0 2088 0 -1 370
box -8 -3 16 105
use FILL  FILL_4853
timestamp 1713400504
transform 1 0 2080 0 -1 370
box -8 -3 16 105
use FILL  FILL_4854
timestamp 1713400504
transform 1 0 2072 0 -1 370
box -8 -3 16 105
use FILL  FILL_4855
timestamp 1713400504
transform 1 0 2040 0 -1 370
box -8 -3 16 105
use FILL  FILL_4856
timestamp 1713400504
transform 1 0 2032 0 -1 370
box -8 -3 16 105
use FILL  FILL_4857
timestamp 1713400504
transform 1 0 2024 0 -1 370
box -8 -3 16 105
use FILL  FILL_4858
timestamp 1713400504
transform 1 0 2016 0 -1 370
box -8 -3 16 105
use FILL  FILL_4859
timestamp 1713400504
transform 1 0 2008 0 -1 370
box -8 -3 16 105
use FILL  FILL_4860
timestamp 1713400504
transform 1 0 1976 0 -1 370
box -8 -3 16 105
use FILL  FILL_4861
timestamp 1713400504
transform 1 0 1968 0 -1 370
box -8 -3 16 105
use FILL  FILL_4862
timestamp 1713400504
transform 1 0 1960 0 -1 370
box -8 -3 16 105
use FILL  FILL_4863
timestamp 1713400504
transform 1 0 1952 0 -1 370
box -8 -3 16 105
use FILL  FILL_4864
timestamp 1713400504
transform 1 0 1944 0 -1 370
box -8 -3 16 105
use FILL  FILL_4865
timestamp 1713400504
transform 1 0 1904 0 -1 370
box -8 -3 16 105
use FILL  FILL_4866
timestamp 1713400504
transform 1 0 1896 0 -1 370
box -8 -3 16 105
use FILL  FILL_4867
timestamp 1713400504
transform 1 0 1888 0 -1 370
box -8 -3 16 105
use FILL  FILL_4868
timestamp 1713400504
transform 1 0 1880 0 -1 370
box -8 -3 16 105
use FILL  FILL_4869
timestamp 1713400504
transform 1 0 1872 0 -1 370
box -8 -3 16 105
use FILL  FILL_4870
timestamp 1713400504
transform 1 0 1864 0 -1 370
box -8 -3 16 105
use FILL  FILL_4871
timestamp 1713400504
transform 1 0 1840 0 -1 370
box -8 -3 16 105
use FILL  FILL_4872
timestamp 1713400504
transform 1 0 1808 0 -1 370
box -8 -3 16 105
use FILL  FILL_4873
timestamp 1713400504
transform 1 0 1800 0 -1 370
box -8 -3 16 105
use FILL  FILL_4874
timestamp 1713400504
transform 1 0 1792 0 -1 370
box -8 -3 16 105
use FILL  FILL_4875
timestamp 1713400504
transform 1 0 1784 0 -1 370
box -8 -3 16 105
use FILL  FILL_4876
timestamp 1713400504
transform 1 0 1776 0 -1 370
box -8 -3 16 105
use FILL  FILL_4877
timestamp 1713400504
transform 1 0 1744 0 -1 370
box -8 -3 16 105
use FILL  FILL_4878
timestamp 1713400504
transform 1 0 1736 0 -1 370
box -8 -3 16 105
use FILL  FILL_4879
timestamp 1713400504
transform 1 0 1728 0 -1 370
box -8 -3 16 105
use FILL  FILL_4880
timestamp 1713400504
transform 1 0 1720 0 -1 370
box -8 -3 16 105
use FILL  FILL_4881
timestamp 1713400504
transform 1 0 1680 0 -1 370
box -8 -3 16 105
use FILL  FILL_4882
timestamp 1713400504
transform 1 0 1672 0 -1 370
box -8 -3 16 105
use FILL  FILL_4883
timestamp 1713400504
transform 1 0 1664 0 -1 370
box -8 -3 16 105
use FILL  FILL_4884
timestamp 1713400504
transform 1 0 1560 0 -1 370
box -8 -3 16 105
use FILL  FILL_4885
timestamp 1713400504
transform 1 0 1552 0 -1 370
box -8 -3 16 105
use FILL  FILL_4886
timestamp 1713400504
transform 1 0 1544 0 -1 370
box -8 -3 16 105
use FILL  FILL_4887
timestamp 1713400504
transform 1 0 1512 0 -1 370
box -8 -3 16 105
use FILL  FILL_4888
timestamp 1713400504
transform 1 0 1504 0 -1 370
box -8 -3 16 105
use FILL  FILL_4889
timestamp 1713400504
transform 1 0 1496 0 -1 370
box -8 -3 16 105
use FILL  FILL_4890
timestamp 1713400504
transform 1 0 1488 0 -1 370
box -8 -3 16 105
use FILL  FILL_4891
timestamp 1713400504
transform 1 0 1480 0 -1 370
box -8 -3 16 105
use FILL  FILL_4892
timestamp 1713400504
transform 1 0 1472 0 -1 370
box -8 -3 16 105
use FILL  FILL_4893
timestamp 1713400504
transform 1 0 1432 0 -1 370
box -8 -3 16 105
use FILL  FILL_4894
timestamp 1713400504
transform 1 0 1424 0 -1 370
box -8 -3 16 105
use FILL  FILL_4895
timestamp 1713400504
transform 1 0 1416 0 -1 370
box -8 -3 16 105
use FILL  FILL_4896
timestamp 1713400504
transform 1 0 1408 0 -1 370
box -8 -3 16 105
use FILL  FILL_4897
timestamp 1713400504
transform 1 0 1400 0 -1 370
box -8 -3 16 105
use FILL  FILL_4898
timestamp 1713400504
transform 1 0 1392 0 -1 370
box -8 -3 16 105
use FILL  FILL_4899
timestamp 1713400504
transform 1 0 1352 0 -1 370
box -8 -3 16 105
use FILL  FILL_4900
timestamp 1713400504
transform 1 0 1344 0 -1 370
box -8 -3 16 105
use FILL  FILL_4901
timestamp 1713400504
transform 1 0 1336 0 -1 370
box -8 -3 16 105
use FILL  FILL_4902
timestamp 1713400504
transform 1 0 1328 0 -1 370
box -8 -3 16 105
use FILL  FILL_4903
timestamp 1713400504
transform 1 0 1320 0 -1 370
box -8 -3 16 105
use FILL  FILL_4904
timestamp 1713400504
transform 1 0 1312 0 -1 370
box -8 -3 16 105
use FILL  FILL_4905
timestamp 1713400504
transform 1 0 1304 0 -1 370
box -8 -3 16 105
use FILL  FILL_4906
timestamp 1713400504
transform 1 0 1256 0 -1 370
box -8 -3 16 105
use FILL  FILL_4907
timestamp 1713400504
transform 1 0 1248 0 -1 370
box -8 -3 16 105
use FILL  FILL_4908
timestamp 1713400504
transform 1 0 1240 0 -1 370
box -8 -3 16 105
use FILL  FILL_4909
timestamp 1713400504
transform 1 0 1232 0 -1 370
box -8 -3 16 105
use FILL  FILL_4910
timestamp 1713400504
transform 1 0 1224 0 -1 370
box -8 -3 16 105
use FILL  FILL_4911
timestamp 1713400504
transform 1 0 1216 0 -1 370
box -8 -3 16 105
use FILL  FILL_4912
timestamp 1713400504
transform 1 0 1208 0 -1 370
box -8 -3 16 105
use FILL  FILL_4913
timestamp 1713400504
transform 1 0 1200 0 -1 370
box -8 -3 16 105
use FILL  FILL_4914
timestamp 1713400504
transform 1 0 1152 0 -1 370
box -8 -3 16 105
use FILL  FILL_4915
timestamp 1713400504
transform 1 0 1144 0 -1 370
box -8 -3 16 105
use FILL  FILL_4916
timestamp 1713400504
transform 1 0 1136 0 -1 370
box -8 -3 16 105
use FILL  FILL_4917
timestamp 1713400504
transform 1 0 1128 0 -1 370
box -8 -3 16 105
use FILL  FILL_4918
timestamp 1713400504
transform 1 0 1024 0 -1 370
box -8 -3 16 105
use FILL  FILL_4919
timestamp 1713400504
transform 1 0 920 0 -1 370
box -8 -3 16 105
use FILL  FILL_4920
timestamp 1713400504
transform 1 0 912 0 -1 370
box -8 -3 16 105
use FILL  FILL_4921
timestamp 1713400504
transform 1 0 904 0 -1 370
box -8 -3 16 105
use FILL  FILL_4922
timestamp 1713400504
transform 1 0 864 0 -1 370
box -8 -3 16 105
use FILL  FILL_4923
timestamp 1713400504
transform 1 0 856 0 -1 370
box -8 -3 16 105
use FILL  FILL_4924
timestamp 1713400504
transform 1 0 848 0 -1 370
box -8 -3 16 105
use FILL  FILL_4925
timestamp 1713400504
transform 1 0 840 0 -1 370
box -8 -3 16 105
use FILL  FILL_4926
timestamp 1713400504
transform 1 0 816 0 -1 370
box -8 -3 16 105
use FILL  FILL_4927
timestamp 1713400504
transform 1 0 808 0 -1 370
box -8 -3 16 105
use FILL  FILL_4928
timestamp 1713400504
transform 1 0 800 0 -1 370
box -8 -3 16 105
use FILL  FILL_4929
timestamp 1713400504
transform 1 0 792 0 -1 370
box -8 -3 16 105
use FILL  FILL_4930
timestamp 1713400504
transform 1 0 752 0 -1 370
box -8 -3 16 105
use FILL  FILL_4931
timestamp 1713400504
transform 1 0 744 0 -1 370
box -8 -3 16 105
use FILL  FILL_4932
timestamp 1713400504
transform 1 0 736 0 -1 370
box -8 -3 16 105
use FILL  FILL_4933
timestamp 1713400504
transform 1 0 728 0 -1 370
box -8 -3 16 105
use FILL  FILL_4934
timestamp 1713400504
transform 1 0 720 0 -1 370
box -8 -3 16 105
use FILL  FILL_4935
timestamp 1713400504
transform 1 0 680 0 -1 370
box -8 -3 16 105
use FILL  FILL_4936
timestamp 1713400504
transform 1 0 672 0 -1 370
box -8 -3 16 105
use FILL  FILL_4937
timestamp 1713400504
transform 1 0 664 0 -1 370
box -8 -3 16 105
use FILL  FILL_4938
timestamp 1713400504
transform 1 0 656 0 -1 370
box -8 -3 16 105
use FILL  FILL_4939
timestamp 1713400504
transform 1 0 616 0 -1 370
box -8 -3 16 105
use FILL  FILL_4940
timestamp 1713400504
transform 1 0 608 0 -1 370
box -8 -3 16 105
use FILL  FILL_4941
timestamp 1713400504
transform 1 0 600 0 -1 370
box -8 -3 16 105
use FILL  FILL_4942
timestamp 1713400504
transform 1 0 592 0 -1 370
box -8 -3 16 105
use FILL  FILL_4943
timestamp 1713400504
transform 1 0 584 0 -1 370
box -8 -3 16 105
use FILL  FILL_4944
timestamp 1713400504
transform 1 0 576 0 -1 370
box -8 -3 16 105
use FILL  FILL_4945
timestamp 1713400504
transform 1 0 536 0 -1 370
box -8 -3 16 105
use FILL  FILL_4946
timestamp 1713400504
transform 1 0 528 0 -1 370
box -8 -3 16 105
use FILL  FILL_4947
timestamp 1713400504
transform 1 0 520 0 -1 370
box -8 -3 16 105
use FILL  FILL_4948
timestamp 1713400504
transform 1 0 496 0 -1 370
box -8 -3 16 105
use FILL  FILL_4949
timestamp 1713400504
transform 1 0 488 0 -1 370
box -8 -3 16 105
use FILL  FILL_4950
timestamp 1713400504
transform 1 0 480 0 -1 370
box -8 -3 16 105
use FILL  FILL_4951
timestamp 1713400504
transform 1 0 472 0 -1 370
box -8 -3 16 105
use FILL  FILL_4952
timestamp 1713400504
transform 1 0 464 0 -1 370
box -8 -3 16 105
use FILL  FILL_4953
timestamp 1713400504
transform 1 0 424 0 -1 370
box -8 -3 16 105
use FILL  FILL_4954
timestamp 1713400504
transform 1 0 416 0 -1 370
box -8 -3 16 105
use FILL  FILL_4955
timestamp 1713400504
transform 1 0 408 0 -1 370
box -8 -3 16 105
use FILL  FILL_4956
timestamp 1713400504
transform 1 0 400 0 -1 370
box -8 -3 16 105
use FILL  FILL_4957
timestamp 1713400504
transform 1 0 392 0 -1 370
box -8 -3 16 105
use FILL  FILL_4958
timestamp 1713400504
transform 1 0 384 0 -1 370
box -8 -3 16 105
use FILL  FILL_4959
timestamp 1713400504
transform 1 0 376 0 -1 370
box -8 -3 16 105
use FILL  FILL_4960
timestamp 1713400504
transform 1 0 328 0 -1 370
box -8 -3 16 105
use FILL  FILL_4961
timestamp 1713400504
transform 1 0 320 0 -1 370
box -8 -3 16 105
use FILL  FILL_4962
timestamp 1713400504
transform 1 0 312 0 -1 370
box -8 -3 16 105
use FILL  FILL_4963
timestamp 1713400504
transform 1 0 304 0 -1 370
box -8 -3 16 105
use FILL  FILL_4964
timestamp 1713400504
transform 1 0 280 0 -1 370
box -8 -3 16 105
use FILL  FILL_4965
timestamp 1713400504
transform 1 0 272 0 -1 370
box -8 -3 16 105
use FILL  FILL_4966
timestamp 1713400504
transform 1 0 264 0 -1 370
box -8 -3 16 105
use FILL  FILL_4967
timestamp 1713400504
transform 1 0 256 0 -1 370
box -8 -3 16 105
use FILL  FILL_4968
timestamp 1713400504
transform 1 0 216 0 -1 370
box -8 -3 16 105
use FILL  FILL_4969
timestamp 1713400504
transform 1 0 208 0 -1 370
box -8 -3 16 105
use FILL  FILL_4970
timestamp 1713400504
transform 1 0 200 0 -1 370
box -8 -3 16 105
use FILL  FILL_4971
timestamp 1713400504
transform 1 0 192 0 -1 370
box -8 -3 16 105
use FILL  FILL_4972
timestamp 1713400504
transform 1 0 184 0 -1 370
box -8 -3 16 105
use FILL  FILL_4973
timestamp 1713400504
transform 1 0 176 0 -1 370
box -8 -3 16 105
use FILL  FILL_4974
timestamp 1713400504
transform 1 0 136 0 -1 370
box -8 -3 16 105
use FILL  FILL_4975
timestamp 1713400504
transform 1 0 128 0 -1 370
box -8 -3 16 105
use FILL  FILL_4976
timestamp 1713400504
transform 1 0 120 0 -1 370
box -8 -3 16 105
use FILL  FILL_4977
timestamp 1713400504
transform 1 0 112 0 -1 370
box -8 -3 16 105
use FILL  FILL_4978
timestamp 1713400504
transform 1 0 104 0 -1 370
box -8 -3 16 105
use FILL  FILL_4979
timestamp 1713400504
transform 1 0 80 0 -1 370
box -8 -3 16 105
use FILL  FILL_4980
timestamp 1713400504
transform 1 0 72 0 -1 370
box -8 -3 16 105
use FILL  FILL_4981
timestamp 1713400504
transform 1 0 3008 0 1 170
box -8 -3 16 105
use FILL  FILL_4982
timestamp 1713400504
transform 1 0 3000 0 1 170
box -8 -3 16 105
use FILL  FILL_4983
timestamp 1713400504
transform 1 0 2992 0 1 170
box -8 -3 16 105
use FILL  FILL_4984
timestamp 1713400504
transform 1 0 2984 0 1 170
box -8 -3 16 105
use FILL  FILL_4985
timestamp 1713400504
transform 1 0 2976 0 1 170
box -8 -3 16 105
use FILL  FILL_4986
timestamp 1713400504
transform 1 0 2936 0 1 170
box -8 -3 16 105
use FILL  FILL_4987
timestamp 1713400504
transform 1 0 2928 0 1 170
box -8 -3 16 105
use FILL  FILL_4988
timestamp 1713400504
transform 1 0 2920 0 1 170
box -8 -3 16 105
use FILL  FILL_4989
timestamp 1713400504
transform 1 0 2912 0 1 170
box -8 -3 16 105
use FILL  FILL_4990
timestamp 1713400504
transform 1 0 2904 0 1 170
box -8 -3 16 105
use FILL  FILL_4991
timestamp 1713400504
transform 1 0 2872 0 1 170
box -8 -3 16 105
use FILL  FILL_4992
timestamp 1713400504
transform 1 0 2864 0 1 170
box -8 -3 16 105
use FILL  FILL_4993
timestamp 1713400504
transform 1 0 2856 0 1 170
box -8 -3 16 105
use FILL  FILL_4994
timestamp 1713400504
transform 1 0 2848 0 1 170
box -8 -3 16 105
use FILL  FILL_4995
timestamp 1713400504
transform 1 0 2840 0 1 170
box -8 -3 16 105
use FILL  FILL_4996
timestamp 1713400504
transform 1 0 2832 0 1 170
box -8 -3 16 105
use FILL  FILL_4997
timestamp 1713400504
transform 1 0 2824 0 1 170
box -8 -3 16 105
use FILL  FILL_4998
timestamp 1713400504
transform 1 0 2816 0 1 170
box -8 -3 16 105
use FILL  FILL_4999
timestamp 1713400504
transform 1 0 2776 0 1 170
box -8 -3 16 105
use FILL  FILL_5000
timestamp 1713400504
transform 1 0 2768 0 1 170
box -8 -3 16 105
use FILL  FILL_5001
timestamp 1713400504
transform 1 0 2760 0 1 170
box -8 -3 16 105
use FILL  FILL_5002
timestamp 1713400504
transform 1 0 2752 0 1 170
box -8 -3 16 105
use FILL  FILL_5003
timestamp 1713400504
transform 1 0 2744 0 1 170
box -8 -3 16 105
use FILL  FILL_5004
timestamp 1713400504
transform 1 0 2736 0 1 170
box -8 -3 16 105
use FILL  FILL_5005
timestamp 1713400504
transform 1 0 2728 0 1 170
box -8 -3 16 105
use FILL  FILL_5006
timestamp 1713400504
transform 1 0 2688 0 1 170
box -8 -3 16 105
use FILL  FILL_5007
timestamp 1713400504
transform 1 0 2680 0 1 170
box -8 -3 16 105
use FILL  FILL_5008
timestamp 1713400504
transform 1 0 2672 0 1 170
box -8 -3 16 105
use FILL  FILL_5009
timestamp 1713400504
transform 1 0 2664 0 1 170
box -8 -3 16 105
use FILL  FILL_5010
timestamp 1713400504
transform 1 0 2656 0 1 170
box -8 -3 16 105
use FILL  FILL_5011
timestamp 1713400504
transform 1 0 2632 0 1 170
box -8 -3 16 105
use FILL  FILL_5012
timestamp 1713400504
transform 1 0 2624 0 1 170
box -8 -3 16 105
use FILL  FILL_5013
timestamp 1713400504
transform 1 0 2520 0 1 170
box -8 -3 16 105
use FILL  FILL_5014
timestamp 1713400504
transform 1 0 2512 0 1 170
box -8 -3 16 105
use FILL  FILL_5015
timestamp 1713400504
transform 1 0 2504 0 1 170
box -8 -3 16 105
use FILL  FILL_5016
timestamp 1713400504
transform 1 0 2496 0 1 170
box -8 -3 16 105
use FILL  FILL_5017
timestamp 1713400504
transform 1 0 2456 0 1 170
box -8 -3 16 105
use FILL  FILL_5018
timestamp 1713400504
transform 1 0 2448 0 1 170
box -8 -3 16 105
use FILL  FILL_5019
timestamp 1713400504
transform 1 0 2440 0 1 170
box -8 -3 16 105
use FILL  FILL_5020
timestamp 1713400504
transform 1 0 2432 0 1 170
box -8 -3 16 105
use FILL  FILL_5021
timestamp 1713400504
transform 1 0 2424 0 1 170
box -8 -3 16 105
use FILL  FILL_5022
timestamp 1713400504
transform 1 0 2400 0 1 170
box -8 -3 16 105
use FILL  FILL_5023
timestamp 1713400504
transform 1 0 2392 0 1 170
box -8 -3 16 105
use FILL  FILL_5024
timestamp 1713400504
transform 1 0 2384 0 1 170
box -8 -3 16 105
use FILL  FILL_5025
timestamp 1713400504
transform 1 0 2376 0 1 170
box -8 -3 16 105
use FILL  FILL_5026
timestamp 1713400504
transform 1 0 2368 0 1 170
box -8 -3 16 105
use FILL  FILL_5027
timestamp 1713400504
transform 1 0 2360 0 1 170
box -8 -3 16 105
use FILL  FILL_5028
timestamp 1713400504
transform 1 0 2320 0 1 170
box -8 -3 16 105
use FILL  FILL_5029
timestamp 1713400504
transform 1 0 2312 0 1 170
box -8 -3 16 105
use FILL  FILL_5030
timestamp 1713400504
transform 1 0 2304 0 1 170
box -8 -3 16 105
use FILL  FILL_5031
timestamp 1713400504
transform 1 0 2296 0 1 170
box -8 -3 16 105
use FILL  FILL_5032
timestamp 1713400504
transform 1 0 2288 0 1 170
box -8 -3 16 105
use FILL  FILL_5033
timestamp 1713400504
transform 1 0 2280 0 1 170
box -8 -3 16 105
use FILL  FILL_5034
timestamp 1713400504
transform 1 0 2272 0 1 170
box -8 -3 16 105
use FILL  FILL_5035
timestamp 1713400504
transform 1 0 2232 0 1 170
box -8 -3 16 105
use FILL  FILL_5036
timestamp 1713400504
transform 1 0 2224 0 1 170
box -8 -3 16 105
use FILL  FILL_5037
timestamp 1713400504
transform 1 0 2216 0 1 170
box -8 -3 16 105
use FILL  FILL_5038
timestamp 1713400504
transform 1 0 2208 0 1 170
box -8 -3 16 105
use FILL  FILL_5039
timestamp 1713400504
transform 1 0 2200 0 1 170
box -8 -3 16 105
use FILL  FILL_5040
timestamp 1713400504
transform 1 0 2192 0 1 170
box -8 -3 16 105
use FILL  FILL_5041
timestamp 1713400504
transform 1 0 2184 0 1 170
box -8 -3 16 105
use FILL  FILL_5042
timestamp 1713400504
transform 1 0 2176 0 1 170
box -8 -3 16 105
use FILL  FILL_5043
timestamp 1713400504
transform 1 0 2168 0 1 170
box -8 -3 16 105
use FILL  FILL_5044
timestamp 1713400504
transform 1 0 2128 0 1 170
box -8 -3 16 105
use FILL  FILL_5045
timestamp 1713400504
transform 1 0 2120 0 1 170
box -8 -3 16 105
use FILL  FILL_5046
timestamp 1713400504
transform 1 0 2112 0 1 170
box -8 -3 16 105
use FILL  FILL_5047
timestamp 1713400504
transform 1 0 2104 0 1 170
box -8 -3 16 105
use FILL  FILL_5048
timestamp 1713400504
transform 1 0 2096 0 1 170
box -8 -3 16 105
use FILL  FILL_5049
timestamp 1713400504
transform 1 0 2088 0 1 170
box -8 -3 16 105
use FILL  FILL_5050
timestamp 1713400504
transform 1 0 2064 0 1 170
box -8 -3 16 105
use FILL  FILL_5051
timestamp 1713400504
transform 1 0 2056 0 1 170
box -8 -3 16 105
use FILL  FILL_5052
timestamp 1713400504
transform 1 0 2048 0 1 170
box -8 -3 16 105
use FILL  FILL_5053
timestamp 1713400504
transform 1 0 2040 0 1 170
box -8 -3 16 105
use FILL  FILL_5054
timestamp 1713400504
transform 1 0 2032 0 1 170
box -8 -3 16 105
use FILL  FILL_5055
timestamp 1713400504
transform 1 0 2024 0 1 170
box -8 -3 16 105
use FILL  FILL_5056
timestamp 1713400504
transform 1 0 1920 0 1 170
box -8 -3 16 105
use FILL  FILL_5057
timestamp 1713400504
transform 1 0 1912 0 1 170
box -8 -3 16 105
use FILL  FILL_5058
timestamp 1713400504
transform 1 0 1904 0 1 170
box -8 -3 16 105
use FILL  FILL_5059
timestamp 1713400504
transform 1 0 1896 0 1 170
box -8 -3 16 105
use FILL  FILL_5060
timestamp 1713400504
transform 1 0 1888 0 1 170
box -8 -3 16 105
use FILL  FILL_5061
timestamp 1713400504
transform 1 0 1864 0 1 170
box -8 -3 16 105
use FILL  FILL_5062
timestamp 1713400504
transform 1 0 1856 0 1 170
box -8 -3 16 105
use FILL  FILL_5063
timestamp 1713400504
transform 1 0 1848 0 1 170
box -8 -3 16 105
use FILL  FILL_5064
timestamp 1713400504
transform 1 0 1840 0 1 170
box -8 -3 16 105
use FILL  FILL_5065
timestamp 1713400504
transform 1 0 1832 0 1 170
box -8 -3 16 105
use FILL  FILL_5066
timestamp 1713400504
transform 1 0 1824 0 1 170
box -8 -3 16 105
use FILL  FILL_5067
timestamp 1713400504
transform 1 0 1816 0 1 170
box -8 -3 16 105
use FILL  FILL_5068
timestamp 1713400504
transform 1 0 1784 0 1 170
box -8 -3 16 105
use FILL  FILL_5069
timestamp 1713400504
transform 1 0 1776 0 1 170
box -8 -3 16 105
use FILL  FILL_5070
timestamp 1713400504
transform 1 0 1768 0 1 170
box -8 -3 16 105
use FILL  FILL_5071
timestamp 1713400504
transform 1 0 1760 0 1 170
box -8 -3 16 105
use FILL  FILL_5072
timestamp 1713400504
transform 1 0 1752 0 1 170
box -8 -3 16 105
use FILL  FILL_5073
timestamp 1713400504
transform 1 0 1744 0 1 170
box -8 -3 16 105
use FILL  FILL_5074
timestamp 1713400504
transform 1 0 1712 0 1 170
box -8 -3 16 105
use FILL  FILL_5075
timestamp 1713400504
transform 1 0 1704 0 1 170
box -8 -3 16 105
use FILL  FILL_5076
timestamp 1713400504
transform 1 0 1696 0 1 170
box -8 -3 16 105
use FILL  FILL_5077
timestamp 1713400504
transform 1 0 1688 0 1 170
box -8 -3 16 105
use FILL  FILL_5078
timestamp 1713400504
transform 1 0 1680 0 1 170
box -8 -3 16 105
use FILL  FILL_5079
timestamp 1713400504
transform 1 0 1672 0 1 170
box -8 -3 16 105
use FILL  FILL_5080
timestamp 1713400504
transform 1 0 1664 0 1 170
box -8 -3 16 105
use FILL  FILL_5081
timestamp 1713400504
transform 1 0 1624 0 1 170
box -8 -3 16 105
use FILL  FILL_5082
timestamp 1713400504
transform 1 0 1616 0 1 170
box -8 -3 16 105
use FILL  FILL_5083
timestamp 1713400504
transform 1 0 1608 0 1 170
box -8 -3 16 105
use FILL  FILL_5084
timestamp 1713400504
transform 1 0 1600 0 1 170
box -8 -3 16 105
use FILL  FILL_5085
timestamp 1713400504
transform 1 0 1592 0 1 170
box -8 -3 16 105
use FILL  FILL_5086
timestamp 1713400504
transform 1 0 1584 0 1 170
box -8 -3 16 105
use FILL  FILL_5087
timestamp 1713400504
transform 1 0 1576 0 1 170
box -8 -3 16 105
use FILL  FILL_5088
timestamp 1713400504
transform 1 0 1568 0 1 170
box -8 -3 16 105
use FILL  FILL_5089
timestamp 1713400504
transform 1 0 1560 0 1 170
box -8 -3 16 105
use FILL  FILL_5090
timestamp 1713400504
transform 1 0 1528 0 1 170
box -8 -3 16 105
use FILL  FILL_5091
timestamp 1713400504
transform 1 0 1520 0 1 170
box -8 -3 16 105
use FILL  FILL_5092
timestamp 1713400504
transform 1 0 1512 0 1 170
box -8 -3 16 105
use FILL  FILL_5093
timestamp 1713400504
transform 1 0 1504 0 1 170
box -8 -3 16 105
use FILL  FILL_5094
timestamp 1713400504
transform 1 0 1496 0 1 170
box -8 -3 16 105
use FILL  FILL_5095
timestamp 1713400504
transform 1 0 1488 0 1 170
box -8 -3 16 105
use FILL  FILL_5096
timestamp 1713400504
transform 1 0 1480 0 1 170
box -8 -3 16 105
use FILL  FILL_5097
timestamp 1713400504
transform 1 0 1472 0 1 170
box -8 -3 16 105
use FILL  FILL_5098
timestamp 1713400504
transform 1 0 1464 0 1 170
box -8 -3 16 105
use FILL  FILL_5099
timestamp 1713400504
transform 1 0 1424 0 1 170
box -8 -3 16 105
use FILL  FILL_5100
timestamp 1713400504
transform 1 0 1416 0 1 170
box -8 -3 16 105
use FILL  FILL_5101
timestamp 1713400504
transform 1 0 1408 0 1 170
box -8 -3 16 105
use FILL  FILL_5102
timestamp 1713400504
transform 1 0 1400 0 1 170
box -8 -3 16 105
use FILL  FILL_5103
timestamp 1713400504
transform 1 0 1392 0 1 170
box -8 -3 16 105
use FILL  FILL_5104
timestamp 1713400504
transform 1 0 1384 0 1 170
box -8 -3 16 105
use FILL  FILL_5105
timestamp 1713400504
transform 1 0 1376 0 1 170
box -8 -3 16 105
use FILL  FILL_5106
timestamp 1713400504
transform 1 0 1368 0 1 170
box -8 -3 16 105
use FILL  FILL_5107
timestamp 1713400504
transform 1 0 1360 0 1 170
box -8 -3 16 105
use FILL  FILL_5108
timestamp 1713400504
transform 1 0 1352 0 1 170
box -8 -3 16 105
use FILL  FILL_5109
timestamp 1713400504
transform 1 0 1344 0 1 170
box -8 -3 16 105
use FILL  FILL_5110
timestamp 1713400504
transform 1 0 1304 0 1 170
box -8 -3 16 105
use FILL  FILL_5111
timestamp 1713400504
transform 1 0 1296 0 1 170
box -8 -3 16 105
use FILL  FILL_5112
timestamp 1713400504
transform 1 0 1288 0 1 170
box -8 -3 16 105
use FILL  FILL_5113
timestamp 1713400504
transform 1 0 1280 0 1 170
box -8 -3 16 105
use FILL  FILL_5114
timestamp 1713400504
transform 1 0 1272 0 1 170
box -8 -3 16 105
use FILL  FILL_5115
timestamp 1713400504
transform 1 0 1264 0 1 170
box -8 -3 16 105
use FILL  FILL_5116
timestamp 1713400504
transform 1 0 1256 0 1 170
box -8 -3 16 105
use FILL  FILL_5117
timestamp 1713400504
transform 1 0 1248 0 1 170
box -8 -3 16 105
use FILL  FILL_5118
timestamp 1713400504
transform 1 0 1240 0 1 170
box -8 -3 16 105
use FILL  FILL_5119
timestamp 1713400504
transform 1 0 1232 0 1 170
box -8 -3 16 105
use FILL  FILL_5120
timestamp 1713400504
transform 1 0 1224 0 1 170
box -8 -3 16 105
use FILL  FILL_5121
timestamp 1713400504
transform 1 0 1216 0 1 170
box -8 -3 16 105
use FILL  FILL_5122
timestamp 1713400504
transform 1 0 1208 0 1 170
box -8 -3 16 105
use FILL  FILL_5123
timestamp 1713400504
transform 1 0 1200 0 1 170
box -8 -3 16 105
use FILL  FILL_5124
timestamp 1713400504
transform 1 0 1192 0 1 170
box -8 -3 16 105
use FILL  FILL_5125
timestamp 1713400504
transform 1 0 1184 0 1 170
box -8 -3 16 105
use FILL  FILL_5126
timestamp 1713400504
transform 1 0 1176 0 1 170
box -8 -3 16 105
use FILL  FILL_5127
timestamp 1713400504
transform 1 0 1152 0 1 170
box -8 -3 16 105
use FILL  FILL_5128
timestamp 1713400504
transform 1 0 1144 0 1 170
box -8 -3 16 105
use FILL  FILL_5129
timestamp 1713400504
transform 1 0 1136 0 1 170
box -8 -3 16 105
use FILL  FILL_5130
timestamp 1713400504
transform 1 0 1128 0 1 170
box -8 -3 16 105
use FILL  FILL_5131
timestamp 1713400504
transform 1 0 1120 0 1 170
box -8 -3 16 105
use FILL  FILL_5132
timestamp 1713400504
transform 1 0 1016 0 1 170
box -8 -3 16 105
use FILL  FILL_5133
timestamp 1713400504
transform 1 0 1008 0 1 170
box -8 -3 16 105
use FILL  FILL_5134
timestamp 1713400504
transform 1 0 1000 0 1 170
box -8 -3 16 105
use FILL  FILL_5135
timestamp 1713400504
transform 1 0 992 0 1 170
box -8 -3 16 105
use FILL  FILL_5136
timestamp 1713400504
transform 1 0 984 0 1 170
box -8 -3 16 105
use FILL  FILL_5137
timestamp 1713400504
transform 1 0 944 0 1 170
box -8 -3 16 105
use FILL  FILL_5138
timestamp 1713400504
transform 1 0 936 0 1 170
box -8 -3 16 105
use FILL  FILL_5139
timestamp 1713400504
transform 1 0 928 0 1 170
box -8 -3 16 105
use FILL  FILL_5140
timestamp 1713400504
transform 1 0 920 0 1 170
box -8 -3 16 105
use FILL  FILL_5141
timestamp 1713400504
transform 1 0 888 0 1 170
box -8 -3 16 105
use FILL  FILL_5142
timestamp 1713400504
transform 1 0 880 0 1 170
box -8 -3 16 105
use FILL  FILL_5143
timestamp 1713400504
transform 1 0 872 0 1 170
box -8 -3 16 105
use FILL  FILL_5144
timestamp 1713400504
transform 1 0 864 0 1 170
box -8 -3 16 105
use FILL  FILL_5145
timestamp 1713400504
transform 1 0 856 0 1 170
box -8 -3 16 105
use FILL  FILL_5146
timestamp 1713400504
transform 1 0 848 0 1 170
box -8 -3 16 105
use FILL  FILL_5147
timestamp 1713400504
transform 1 0 808 0 1 170
box -8 -3 16 105
use FILL  FILL_5148
timestamp 1713400504
transform 1 0 800 0 1 170
box -8 -3 16 105
use FILL  FILL_5149
timestamp 1713400504
transform 1 0 792 0 1 170
box -8 -3 16 105
use FILL  FILL_5150
timestamp 1713400504
transform 1 0 784 0 1 170
box -8 -3 16 105
use FILL  FILL_5151
timestamp 1713400504
transform 1 0 776 0 1 170
box -8 -3 16 105
use FILL  FILL_5152
timestamp 1713400504
transform 1 0 744 0 1 170
box -8 -3 16 105
use FILL  FILL_5153
timestamp 1713400504
transform 1 0 736 0 1 170
box -8 -3 16 105
use FILL  FILL_5154
timestamp 1713400504
transform 1 0 728 0 1 170
box -8 -3 16 105
use FILL  FILL_5155
timestamp 1713400504
transform 1 0 720 0 1 170
box -8 -3 16 105
use FILL  FILL_5156
timestamp 1713400504
transform 1 0 712 0 1 170
box -8 -3 16 105
use FILL  FILL_5157
timestamp 1713400504
transform 1 0 704 0 1 170
box -8 -3 16 105
use FILL  FILL_5158
timestamp 1713400504
transform 1 0 664 0 1 170
box -8 -3 16 105
use FILL  FILL_5159
timestamp 1713400504
transform 1 0 656 0 1 170
box -8 -3 16 105
use FILL  FILL_5160
timestamp 1713400504
transform 1 0 648 0 1 170
box -8 -3 16 105
use FILL  FILL_5161
timestamp 1713400504
transform 1 0 640 0 1 170
box -8 -3 16 105
use FILL  FILL_5162
timestamp 1713400504
transform 1 0 632 0 1 170
box -8 -3 16 105
use FILL  FILL_5163
timestamp 1713400504
transform 1 0 624 0 1 170
box -8 -3 16 105
use FILL  FILL_5164
timestamp 1713400504
transform 1 0 592 0 1 170
box -8 -3 16 105
use FILL  FILL_5165
timestamp 1713400504
transform 1 0 584 0 1 170
box -8 -3 16 105
use FILL  FILL_5166
timestamp 1713400504
transform 1 0 576 0 1 170
box -8 -3 16 105
use FILL  FILL_5167
timestamp 1713400504
transform 1 0 536 0 1 170
box -8 -3 16 105
use FILL  FILL_5168
timestamp 1713400504
transform 1 0 528 0 1 170
box -8 -3 16 105
use FILL  FILL_5169
timestamp 1713400504
transform 1 0 520 0 1 170
box -8 -3 16 105
use FILL  FILL_5170
timestamp 1713400504
transform 1 0 416 0 1 170
box -8 -3 16 105
use FILL  FILL_5171
timestamp 1713400504
transform 1 0 408 0 1 170
box -8 -3 16 105
use FILL  FILL_5172
timestamp 1713400504
transform 1 0 400 0 1 170
box -8 -3 16 105
use FILL  FILL_5173
timestamp 1713400504
transform 1 0 344 0 1 170
box -8 -3 16 105
use FILL  FILL_5174
timestamp 1713400504
transform 1 0 336 0 1 170
box -8 -3 16 105
use FILL  FILL_5175
timestamp 1713400504
transform 1 0 328 0 1 170
box -8 -3 16 105
use FILL  FILL_5176
timestamp 1713400504
transform 1 0 320 0 1 170
box -8 -3 16 105
use FILL  FILL_5177
timestamp 1713400504
transform 1 0 312 0 1 170
box -8 -3 16 105
use FILL  FILL_5178
timestamp 1713400504
transform 1 0 304 0 1 170
box -8 -3 16 105
use FILL  FILL_5179
timestamp 1713400504
transform 1 0 264 0 1 170
box -8 -3 16 105
use FILL  FILL_5180
timestamp 1713400504
transform 1 0 256 0 1 170
box -8 -3 16 105
use FILL  FILL_5181
timestamp 1713400504
transform 1 0 248 0 1 170
box -8 -3 16 105
use FILL  FILL_5182
timestamp 1713400504
transform 1 0 240 0 1 170
box -8 -3 16 105
use FILL  FILL_5183
timestamp 1713400504
transform 1 0 208 0 1 170
box -8 -3 16 105
use FILL  FILL_5184
timestamp 1713400504
transform 1 0 200 0 1 170
box -8 -3 16 105
use FILL  FILL_5185
timestamp 1713400504
transform 1 0 192 0 1 170
box -8 -3 16 105
use FILL  FILL_5186
timestamp 1713400504
transform 1 0 152 0 1 170
box -8 -3 16 105
use FILL  FILL_5187
timestamp 1713400504
transform 1 0 144 0 1 170
box -8 -3 16 105
use FILL  FILL_5188
timestamp 1713400504
transform 1 0 136 0 1 170
box -8 -3 16 105
use FILL  FILL_5189
timestamp 1713400504
transform 1 0 128 0 1 170
box -8 -3 16 105
use FILL  FILL_5190
timestamp 1713400504
transform 1 0 120 0 1 170
box -8 -3 16 105
use FILL  FILL_5191
timestamp 1713400504
transform 1 0 80 0 1 170
box -8 -3 16 105
use FILL  FILL_5192
timestamp 1713400504
transform 1 0 72 0 1 170
box -8 -3 16 105
use FILL  FILL_5193
timestamp 1713400504
transform 1 0 3008 0 -1 170
box -8 -3 16 105
use FILL  FILL_5194
timestamp 1713400504
transform 1 0 3000 0 -1 170
box -8 -3 16 105
use FILL  FILL_5195
timestamp 1713400504
transform 1 0 2992 0 -1 170
box -8 -3 16 105
use FILL  FILL_5196
timestamp 1713400504
transform 1 0 2960 0 -1 170
box -8 -3 16 105
use FILL  FILL_5197
timestamp 1713400504
transform 1 0 2952 0 -1 170
box -8 -3 16 105
use FILL  FILL_5198
timestamp 1713400504
transform 1 0 2944 0 -1 170
box -8 -3 16 105
use FILL  FILL_5199
timestamp 1713400504
transform 1 0 2936 0 -1 170
box -8 -3 16 105
use FILL  FILL_5200
timestamp 1713400504
transform 1 0 2912 0 -1 170
box -8 -3 16 105
use FILL  FILL_5201
timestamp 1713400504
transform 1 0 2904 0 -1 170
box -8 -3 16 105
use FILL  FILL_5202
timestamp 1713400504
transform 1 0 2896 0 -1 170
box -8 -3 16 105
use FILL  FILL_5203
timestamp 1713400504
transform 1 0 2888 0 -1 170
box -8 -3 16 105
use FILL  FILL_5204
timestamp 1713400504
transform 1 0 2880 0 -1 170
box -8 -3 16 105
use FILL  FILL_5205
timestamp 1713400504
transform 1 0 2840 0 -1 170
box -8 -3 16 105
use FILL  FILL_5206
timestamp 1713400504
transform 1 0 2832 0 -1 170
box -8 -3 16 105
use FILL  FILL_5207
timestamp 1713400504
transform 1 0 2824 0 -1 170
box -8 -3 16 105
use FILL  FILL_5208
timestamp 1713400504
transform 1 0 2816 0 -1 170
box -8 -3 16 105
use FILL  FILL_5209
timestamp 1713400504
transform 1 0 2808 0 -1 170
box -8 -3 16 105
use FILL  FILL_5210
timestamp 1713400504
transform 1 0 2800 0 -1 170
box -8 -3 16 105
use FILL  FILL_5211
timestamp 1713400504
transform 1 0 2792 0 -1 170
box -8 -3 16 105
use FILL  FILL_5212
timestamp 1713400504
transform 1 0 2784 0 -1 170
box -8 -3 16 105
use FILL  FILL_5213
timestamp 1713400504
transform 1 0 2736 0 -1 170
box -8 -3 16 105
use FILL  FILL_5214
timestamp 1713400504
transform 1 0 2728 0 -1 170
box -8 -3 16 105
use FILL  FILL_5215
timestamp 1713400504
transform 1 0 2720 0 -1 170
box -8 -3 16 105
use FILL  FILL_5216
timestamp 1713400504
transform 1 0 2712 0 -1 170
box -8 -3 16 105
use FILL  FILL_5217
timestamp 1713400504
transform 1 0 2704 0 -1 170
box -8 -3 16 105
use FILL  FILL_5218
timestamp 1713400504
transform 1 0 2680 0 -1 170
box -8 -3 16 105
use FILL  FILL_5219
timestamp 1713400504
transform 1 0 2672 0 -1 170
box -8 -3 16 105
use FILL  FILL_5220
timestamp 1713400504
transform 1 0 2664 0 -1 170
box -8 -3 16 105
use FILL  FILL_5221
timestamp 1713400504
transform 1 0 2656 0 -1 170
box -8 -3 16 105
use FILL  FILL_5222
timestamp 1713400504
transform 1 0 2648 0 -1 170
box -8 -3 16 105
use FILL  FILL_5223
timestamp 1713400504
transform 1 0 2608 0 -1 170
box -8 -3 16 105
use FILL  FILL_5224
timestamp 1713400504
transform 1 0 2600 0 -1 170
box -8 -3 16 105
use FILL  FILL_5225
timestamp 1713400504
transform 1 0 2592 0 -1 170
box -8 -3 16 105
use FILL  FILL_5226
timestamp 1713400504
transform 1 0 2584 0 -1 170
box -8 -3 16 105
use FILL  FILL_5227
timestamp 1713400504
transform 1 0 2576 0 -1 170
box -8 -3 16 105
use FILL  FILL_5228
timestamp 1713400504
transform 1 0 2544 0 -1 170
box -8 -3 16 105
use FILL  FILL_5229
timestamp 1713400504
transform 1 0 2536 0 -1 170
box -8 -3 16 105
use FILL  FILL_5230
timestamp 1713400504
transform 1 0 2528 0 -1 170
box -8 -3 16 105
use FILL  FILL_5231
timestamp 1713400504
transform 1 0 2424 0 -1 170
box -8 -3 16 105
use FILL  FILL_5232
timestamp 1713400504
transform 1 0 2416 0 -1 170
box -8 -3 16 105
use FILL  FILL_5233
timestamp 1713400504
transform 1 0 2408 0 -1 170
box -8 -3 16 105
use FILL  FILL_5234
timestamp 1713400504
transform 1 0 2304 0 -1 170
box -8 -3 16 105
use FILL  FILL_5235
timestamp 1713400504
transform 1 0 2296 0 -1 170
box -8 -3 16 105
use FILL  FILL_5236
timestamp 1713400504
transform 1 0 2288 0 -1 170
box -8 -3 16 105
use FILL  FILL_5237
timestamp 1713400504
transform 1 0 2280 0 -1 170
box -8 -3 16 105
use FILL  FILL_5238
timestamp 1713400504
transform 1 0 2240 0 -1 170
box -8 -3 16 105
use FILL  FILL_5239
timestamp 1713400504
transform 1 0 2232 0 -1 170
box -8 -3 16 105
use FILL  FILL_5240
timestamp 1713400504
transform 1 0 2224 0 -1 170
box -8 -3 16 105
use FILL  FILL_5241
timestamp 1713400504
transform 1 0 2216 0 -1 170
box -8 -3 16 105
use FILL  FILL_5242
timestamp 1713400504
transform 1 0 2208 0 -1 170
box -8 -3 16 105
use FILL  FILL_5243
timestamp 1713400504
transform 1 0 2200 0 -1 170
box -8 -3 16 105
use FILL  FILL_5244
timestamp 1713400504
transform 1 0 2192 0 -1 170
box -8 -3 16 105
use FILL  FILL_5245
timestamp 1713400504
transform 1 0 2184 0 -1 170
box -8 -3 16 105
use FILL  FILL_5246
timestamp 1713400504
transform 1 0 2144 0 -1 170
box -8 -3 16 105
use FILL  FILL_5247
timestamp 1713400504
transform 1 0 2136 0 -1 170
box -8 -3 16 105
use FILL  FILL_5248
timestamp 1713400504
transform 1 0 2128 0 -1 170
box -8 -3 16 105
use FILL  FILL_5249
timestamp 1713400504
transform 1 0 2120 0 -1 170
box -8 -3 16 105
use FILL  FILL_5250
timestamp 1713400504
transform 1 0 2112 0 -1 170
box -8 -3 16 105
use FILL  FILL_5251
timestamp 1713400504
transform 1 0 2104 0 -1 170
box -8 -3 16 105
use FILL  FILL_5252
timestamp 1713400504
transform 1 0 2096 0 -1 170
box -8 -3 16 105
use FILL  FILL_5253
timestamp 1713400504
transform 1 0 2056 0 -1 170
box -8 -3 16 105
use FILL  FILL_5254
timestamp 1713400504
transform 1 0 2048 0 -1 170
box -8 -3 16 105
use FILL  FILL_5255
timestamp 1713400504
transform 1 0 2040 0 -1 170
box -8 -3 16 105
use FILL  FILL_5256
timestamp 1713400504
transform 1 0 2032 0 -1 170
box -8 -3 16 105
use FILL  FILL_5257
timestamp 1713400504
transform 1 0 2024 0 -1 170
box -8 -3 16 105
use FILL  FILL_5258
timestamp 1713400504
transform 1 0 1920 0 -1 170
box -8 -3 16 105
use FILL  FILL_5259
timestamp 1713400504
transform 1 0 1912 0 -1 170
box -8 -3 16 105
use FILL  FILL_5260
timestamp 1713400504
transform 1 0 1904 0 -1 170
box -8 -3 16 105
use FILL  FILL_5261
timestamp 1713400504
transform 1 0 1896 0 -1 170
box -8 -3 16 105
use FILL  FILL_5262
timestamp 1713400504
transform 1 0 1864 0 -1 170
box -8 -3 16 105
use FILL  FILL_5263
timestamp 1713400504
transform 1 0 1856 0 -1 170
box -8 -3 16 105
use FILL  FILL_5264
timestamp 1713400504
transform 1 0 1848 0 -1 170
box -8 -3 16 105
use FILL  FILL_5265
timestamp 1713400504
transform 1 0 1816 0 -1 170
box -8 -3 16 105
use FILL  FILL_5266
timestamp 1713400504
transform 1 0 1808 0 -1 170
box -8 -3 16 105
use FILL  FILL_5267
timestamp 1713400504
transform 1 0 1800 0 -1 170
box -8 -3 16 105
use FILL  FILL_5268
timestamp 1713400504
transform 1 0 1696 0 -1 170
box -8 -3 16 105
use FILL  FILL_5269
timestamp 1713400504
transform 1 0 1688 0 -1 170
box -8 -3 16 105
use FILL  FILL_5270
timestamp 1713400504
transform 1 0 1680 0 -1 170
box -8 -3 16 105
use FILL  FILL_5271
timestamp 1713400504
transform 1 0 1648 0 -1 170
box -8 -3 16 105
use FILL  FILL_5272
timestamp 1713400504
transform 1 0 1640 0 -1 170
box -8 -3 16 105
use FILL  FILL_5273
timestamp 1713400504
transform 1 0 1632 0 -1 170
box -8 -3 16 105
use FILL  FILL_5274
timestamp 1713400504
transform 1 0 1624 0 -1 170
box -8 -3 16 105
use FILL  FILL_5275
timestamp 1713400504
transform 1 0 1616 0 -1 170
box -8 -3 16 105
use FILL  FILL_5276
timestamp 1713400504
transform 1 0 1576 0 -1 170
box -8 -3 16 105
use FILL  FILL_5277
timestamp 1713400504
transform 1 0 1568 0 -1 170
box -8 -3 16 105
use FILL  FILL_5278
timestamp 1713400504
transform 1 0 1560 0 -1 170
box -8 -3 16 105
use FILL  FILL_5279
timestamp 1713400504
transform 1 0 1456 0 -1 170
box -8 -3 16 105
use FILL  FILL_5280
timestamp 1713400504
transform 1 0 1448 0 -1 170
box -8 -3 16 105
use FILL  FILL_5281
timestamp 1713400504
transform 1 0 1440 0 -1 170
box -8 -3 16 105
use FILL  FILL_5282
timestamp 1713400504
transform 1 0 1416 0 -1 170
box -8 -3 16 105
use FILL  FILL_5283
timestamp 1713400504
transform 1 0 1408 0 -1 170
box -8 -3 16 105
use FILL  FILL_5284
timestamp 1713400504
transform 1 0 1400 0 -1 170
box -8 -3 16 105
use FILL  FILL_5285
timestamp 1713400504
transform 1 0 1360 0 -1 170
box -8 -3 16 105
use FILL  FILL_5286
timestamp 1713400504
transform 1 0 1352 0 -1 170
box -8 -3 16 105
use FILL  FILL_5287
timestamp 1713400504
transform 1 0 1344 0 -1 170
box -8 -3 16 105
use FILL  FILL_5288
timestamp 1713400504
transform 1 0 1336 0 -1 170
box -8 -3 16 105
use FILL  FILL_5289
timestamp 1713400504
transform 1 0 1328 0 -1 170
box -8 -3 16 105
use FILL  FILL_5290
timestamp 1713400504
transform 1 0 1320 0 -1 170
box -8 -3 16 105
use FILL  FILL_5291
timestamp 1713400504
transform 1 0 1312 0 -1 170
box -8 -3 16 105
use FILL  FILL_5292
timestamp 1713400504
transform 1 0 1304 0 -1 170
box -8 -3 16 105
use FILL  FILL_5293
timestamp 1713400504
transform 1 0 1272 0 -1 170
box -8 -3 16 105
use FILL  FILL_5294
timestamp 1713400504
transform 1 0 1264 0 -1 170
box -8 -3 16 105
use FILL  FILL_5295
timestamp 1713400504
transform 1 0 1256 0 -1 170
box -8 -3 16 105
use FILL  FILL_5296
timestamp 1713400504
transform 1 0 1248 0 -1 170
box -8 -3 16 105
use FILL  FILL_5297
timestamp 1713400504
transform 1 0 1240 0 -1 170
box -8 -3 16 105
use FILL  FILL_5298
timestamp 1713400504
transform 1 0 1232 0 -1 170
box -8 -3 16 105
use FILL  FILL_5299
timestamp 1713400504
transform 1 0 1224 0 -1 170
box -8 -3 16 105
use FILL  FILL_5300
timestamp 1713400504
transform 1 0 1120 0 -1 170
box -8 -3 16 105
use FILL  FILL_5301
timestamp 1713400504
transform 1 0 1112 0 -1 170
box -8 -3 16 105
use FILL  FILL_5302
timestamp 1713400504
transform 1 0 1104 0 -1 170
box -8 -3 16 105
use FILL  FILL_5303
timestamp 1713400504
transform 1 0 1096 0 -1 170
box -8 -3 16 105
use FILL  FILL_5304
timestamp 1713400504
transform 1 0 1064 0 -1 170
box -8 -3 16 105
use FILL  FILL_5305
timestamp 1713400504
transform 1 0 1056 0 -1 170
box -8 -3 16 105
use FILL  FILL_5306
timestamp 1713400504
transform 1 0 1048 0 -1 170
box -8 -3 16 105
use FILL  FILL_5307
timestamp 1713400504
transform 1 0 1040 0 -1 170
box -8 -3 16 105
use FILL  FILL_5308
timestamp 1713400504
transform 1 0 1032 0 -1 170
box -8 -3 16 105
use FILL  FILL_5309
timestamp 1713400504
transform 1 0 1024 0 -1 170
box -8 -3 16 105
use FILL  FILL_5310
timestamp 1713400504
transform 1 0 984 0 -1 170
box -8 -3 16 105
use FILL  FILL_5311
timestamp 1713400504
transform 1 0 976 0 -1 170
box -8 -3 16 105
use FILL  FILL_5312
timestamp 1713400504
transform 1 0 968 0 -1 170
box -8 -3 16 105
use FILL  FILL_5313
timestamp 1713400504
transform 1 0 960 0 -1 170
box -8 -3 16 105
use FILL  FILL_5314
timestamp 1713400504
transform 1 0 952 0 -1 170
box -8 -3 16 105
use FILL  FILL_5315
timestamp 1713400504
transform 1 0 944 0 -1 170
box -8 -3 16 105
use FILL  FILL_5316
timestamp 1713400504
transform 1 0 904 0 -1 170
box -8 -3 16 105
use FILL  FILL_5317
timestamp 1713400504
transform 1 0 896 0 -1 170
box -8 -3 16 105
use FILL  FILL_5318
timestamp 1713400504
transform 1 0 888 0 -1 170
box -8 -3 16 105
use FILL  FILL_5319
timestamp 1713400504
transform 1 0 880 0 -1 170
box -8 -3 16 105
use FILL  FILL_5320
timestamp 1713400504
transform 1 0 776 0 -1 170
box -8 -3 16 105
use FILL  FILL_5321
timestamp 1713400504
transform 1 0 768 0 -1 170
box -8 -3 16 105
use FILL  FILL_5322
timestamp 1713400504
transform 1 0 760 0 -1 170
box -8 -3 16 105
use FILL  FILL_5323
timestamp 1713400504
transform 1 0 752 0 -1 170
box -8 -3 16 105
use FILL  FILL_5324
timestamp 1713400504
transform 1 0 720 0 -1 170
box -8 -3 16 105
use FILL  FILL_5325
timestamp 1713400504
transform 1 0 680 0 -1 170
box -8 -3 16 105
use FILL  FILL_5326
timestamp 1713400504
transform 1 0 672 0 -1 170
box -8 -3 16 105
use FILL  FILL_5327
timestamp 1713400504
transform 1 0 664 0 -1 170
box -8 -3 16 105
use FILL  FILL_5328
timestamp 1713400504
transform 1 0 560 0 -1 170
box -8 -3 16 105
use FILL  FILL_5329
timestamp 1713400504
transform 1 0 456 0 -1 170
box -8 -3 16 105
use FILL  FILL_5330
timestamp 1713400504
transform 1 0 448 0 -1 170
box -8 -3 16 105
use FILL  FILL_5331
timestamp 1713400504
transform 1 0 384 0 -1 170
box -8 -3 16 105
use FILL  FILL_5332
timestamp 1713400504
transform 1 0 344 0 -1 170
box -8 -3 16 105
use FILL  FILL_5333
timestamp 1713400504
transform 1 0 336 0 -1 170
box -8 -3 16 105
use FILL  FILL_5334
timestamp 1713400504
transform 1 0 328 0 -1 170
box -8 -3 16 105
use FILL  FILL_5335
timestamp 1713400504
transform 1 0 264 0 -1 170
box -8 -3 16 105
use FILL  FILL_5336
timestamp 1713400504
transform 1 0 256 0 -1 170
box -8 -3 16 105
use FILL  FILL_5337
timestamp 1713400504
transform 1 0 176 0 -1 170
box -8 -3 16 105
use FILL  FILL_5338
timestamp 1713400504
transform 1 0 72 0 -1 170
box -8 -3 16 105
use HAX1  HAX1_0
timestamp 1713400504
transform 1 0 2928 0 1 770
box -5 -3 84 105
use HAX1  HAX1_1
timestamp 1713400504
transform 1 0 2760 0 1 770
box -5 -3 84 105
use HAX1  HAX1_2
timestamp 1713400504
transform 1 0 2816 0 1 970
box -5 -3 84 105
use HAX1  HAX1_3
timestamp 1713400504
transform 1 0 2808 0 -1 1170
box -5 -3 84 105
use HAX1  HAX1_4
timestamp 1713400504
transform 1 0 2912 0 1 1170
box -5 -3 84 105
use HAX1  HAX1_5
timestamp 1713400504
transform 1 0 2808 0 -1 1370
box -5 -3 84 105
use HAX1  HAX1_6
timestamp 1713400504
transform 1 0 424 0 1 2170
box -5 -3 84 105
use HAX1  HAX1_7
timestamp 1713400504
transform 1 0 720 0 -1 2370
box -5 -3 84 105
use HAX1  HAX1_8
timestamp 1713400504
transform 1 0 384 0 -1 2170
box -5 -3 84 105
use HAX1  HAX1_9
timestamp 1713400504
transform 1 0 680 0 -1 2970
box -5 -3 84 105
use HAX1  HAX1_10
timestamp 1713400504
transform 1 0 840 0 -1 2970
box -5 -3 84 105
use HAX1  HAX1_11
timestamp 1713400504
transform 1 0 344 0 1 2770
box -5 -3 84 105
use HAX1  HAX1_12
timestamp 1713400504
transform 1 0 320 0 -1 2970
box -5 -3 84 105
use HAX1  HAX1_13
timestamp 1713400504
transform 1 0 144 0 -1 2770
box -5 -3 84 105
use HAX1  HAX1_14
timestamp 1713400504
transform 1 0 144 0 1 2770
box -5 -3 84 105
use HAX1  HAX1_15
timestamp 1713400504
transform 1 0 80 0 1 1970
box -5 -3 84 105
use HAX1  HAX1_16
timestamp 1713400504
transform 1 0 80 0 -1 2170
box -5 -3 84 105
use INVX1  INVX1_0
timestamp 1713400504
transform 1 0 1600 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_0
timestamp 1713400504
transform 1 0 1424 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_1
timestamp 1713400504
transform 1 0 80 0 1 370
box -9 -3 26 105
use INVX2  INVX2_2
timestamp 1713400504
transform 1 0 552 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_3
timestamp 1713400504
transform 1 0 384 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_4
timestamp 1713400504
transform 1 0 432 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_5
timestamp 1713400504
transform 1 0 456 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_6
timestamp 1713400504
transform 1 0 488 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_7
timestamp 1713400504
transform 1 0 2848 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_8
timestamp 1713400504
transform 1 0 1440 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_9
timestamp 1713400504
transform 1 0 2792 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_10
timestamp 1713400504
transform 1 0 2112 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_11
timestamp 1713400504
transform 1 0 1376 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_12
timestamp 1713400504
transform 1 0 1776 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_13
timestamp 1713400504
transform 1 0 1112 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_14
timestamp 1713400504
transform 1 0 1688 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_15
timestamp 1713400504
transform 1 0 1840 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_16
timestamp 1713400504
transform 1 0 1656 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_17
timestamp 1713400504
transform 1 0 2192 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_18
timestamp 1713400504
transform 1 0 1528 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_19
timestamp 1713400504
transform 1 0 1640 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_20
timestamp 1713400504
transform 1 0 1584 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_21
timestamp 1713400504
transform 1 0 1624 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_22
timestamp 1713400504
transform 1 0 1480 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_23
timestamp 1713400504
transform 1 0 1312 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_24
timestamp 1713400504
transform 1 0 1400 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_25
timestamp 1713400504
transform 1 0 184 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_26
timestamp 1713400504
transform 1 0 384 0 1 170
box -9 -3 26 105
use INVX2  INVX2_27
timestamp 1713400504
transform 1 0 1464 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_28
timestamp 1713400504
transform 1 0 1168 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_29
timestamp 1713400504
transform 1 0 2160 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_30
timestamp 1713400504
transform 1 0 2552 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_31
timestamp 1713400504
transform 1 0 2488 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_32
timestamp 1713400504
transform 1 0 1864 0 1 770
box -9 -3 26 105
use INVX2  INVX2_33
timestamp 1713400504
transform 1 0 1784 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_34
timestamp 1713400504
transform 1 0 1736 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_35
timestamp 1713400504
transform 1 0 1720 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_36
timestamp 1713400504
transform 1 0 1448 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_37
timestamp 1713400504
transform 1 0 1048 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_38
timestamp 1713400504
transform 1 0 1216 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_39
timestamp 1713400504
transform 1 0 1040 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_40
timestamp 1713400504
transform 1 0 800 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_41
timestamp 1713400504
transform 1 0 1296 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_42
timestamp 1713400504
transform 1 0 2040 0 1 970
box -9 -3 26 105
use INVX2  INVX2_43
timestamp 1713400504
transform 1 0 1616 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_44
timestamp 1713400504
transform 1 0 1848 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_45
timestamp 1713400504
transform 1 0 1856 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_46
timestamp 1713400504
transform 1 0 2176 0 1 970
box -9 -3 26 105
use INVX2  INVX2_47
timestamp 1713400504
transform 1 0 2104 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_48
timestamp 1713400504
transform 1 0 1808 0 1 970
box -9 -3 26 105
use INVX2  INVX2_49
timestamp 1713400504
transform 1 0 1800 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_50
timestamp 1713400504
transform 1 0 2216 0 1 970
box -9 -3 26 105
use INVX2  INVX2_51
timestamp 1713400504
transform 1 0 2192 0 1 770
box -9 -3 26 105
use INVX2  INVX2_52
timestamp 1713400504
transform 1 0 2024 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_53
timestamp 1713400504
transform 1 0 1184 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_54
timestamp 1713400504
transform 1 0 936 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_55
timestamp 1713400504
transform 1 0 1096 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_56
timestamp 1713400504
transform 1 0 1896 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_57
timestamp 1713400504
transform 1 0 2080 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_58
timestamp 1713400504
transform 1 0 2112 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_59
timestamp 1713400504
transform 1 0 1736 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_60
timestamp 1713400504
transform 1 0 2424 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_61
timestamp 1713400504
transform 1 0 1760 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_62
timestamp 1713400504
transform 1 0 1656 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_63
timestamp 1713400504
transform 1 0 1480 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_64
timestamp 1713400504
transform 1 0 2480 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_65
timestamp 1713400504
transform 1 0 1408 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_66
timestamp 1713400504
transform 1 0 1528 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_67
timestamp 1713400504
transform 1 0 1408 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_68
timestamp 1713400504
transform 1 0 1488 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_69
timestamp 1713400504
transform 1 0 1928 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_70
timestamp 1713400504
transform 1 0 1944 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_71
timestamp 1713400504
transform 1 0 2192 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_72
timestamp 1713400504
transform 1 0 2384 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_73
timestamp 1713400504
transform 1 0 2496 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_74
timestamp 1713400504
transform 1 0 2288 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_75
timestamp 1713400504
transform 1 0 2416 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_76
timestamp 1713400504
transform 1 0 2832 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_77
timestamp 1713400504
transform 1 0 2736 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_78
timestamp 1713400504
transform 1 0 2616 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_79
timestamp 1713400504
transform 1 0 2864 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_80
timestamp 1713400504
transform 1 0 2496 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_81
timestamp 1713400504
transform 1 0 2472 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_82
timestamp 1713400504
transform 1 0 2576 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_83
timestamp 1713400504
transform 1 0 2672 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_84
timestamp 1713400504
transform 1 0 2976 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_85
timestamp 1713400504
transform 1 0 2952 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_86
timestamp 1713400504
transform 1 0 2712 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_87
timestamp 1713400504
transform 1 0 2216 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_88
timestamp 1713400504
transform 1 0 2336 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_89
timestamp 1713400504
transform 1 0 2384 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_90
timestamp 1713400504
transform 1 0 2488 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_91
timestamp 1713400504
transform 1 0 2376 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_92
timestamp 1713400504
transform 1 0 1872 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_93
timestamp 1713400504
transform 1 0 2088 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_94
timestamp 1713400504
transform 1 0 1552 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_95
timestamp 1713400504
transform 1 0 1400 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_96
timestamp 1713400504
transform 1 0 1664 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_97
timestamp 1713400504
transform 1 0 1352 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_98
timestamp 1713400504
transform 1 0 1184 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_99
timestamp 1713400504
transform 1 0 1168 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_100
timestamp 1713400504
transform 1 0 1288 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_101
timestamp 1713400504
transform 1 0 1168 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_102
timestamp 1713400504
transform 1 0 1752 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_103
timestamp 1713400504
transform 1 0 1944 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_104
timestamp 1713400504
transform 1 0 2096 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_105
timestamp 1713400504
transform 1 0 2528 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_106
timestamp 1713400504
transform 1 0 2704 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_107
timestamp 1713400504
transform 1 0 2784 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_108
timestamp 1713400504
transform 1 0 2976 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_109
timestamp 1713400504
transform 1 0 2888 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_110
timestamp 1713400504
transform 1 0 2904 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_111
timestamp 1713400504
transform 1 0 2576 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_112
timestamp 1713400504
transform 1 0 2728 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_113
timestamp 1713400504
transform 1 0 2872 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_114
timestamp 1713400504
transform 1 0 2992 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_115
timestamp 1713400504
transform 1 0 2984 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_116
timestamp 1713400504
transform 1 0 2872 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_117
timestamp 1713400504
transform 1 0 2864 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_118
timestamp 1713400504
transform 1 0 2608 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_119
timestamp 1713400504
transform 1 0 2872 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_120
timestamp 1713400504
transform 1 0 2392 0 1 370
box -9 -3 26 105
use INVX2  INVX2_121
timestamp 1713400504
transform 1 0 2680 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_122
timestamp 1713400504
transform 1 0 2240 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_123
timestamp 1713400504
transform 1 0 2416 0 1 370
box -9 -3 26 105
use INVX2  INVX2_124
timestamp 1713400504
transform 1 0 2408 0 1 170
box -9 -3 26 105
use INVX2  INVX2_125
timestamp 1713400504
transform 1 0 2912 0 1 570
box -9 -3 26 105
use INVX2  INVX2_126
timestamp 1713400504
transform 1 0 2640 0 1 170
box -9 -3 26 105
use INVX2  INVX2_127
timestamp 1713400504
transform 1 0 2872 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_128
timestamp 1713400504
transform 1 0 2920 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_129
timestamp 1713400504
transform 1 0 2688 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_130
timestamp 1713400504
transform 1 0 2216 0 1 370
box -9 -3 26 105
use INVX2  INVX2_131
timestamp 1713400504
transform 1 0 2072 0 1 170
box -9 -3 26 105
use INVX2  INVX2_132
timestamp 1713400504
transform 1 0 1872 0 1 170
box -9 -3 26 105
use INVX2  INVX2_133
timestamp 1713400504
transform 1 0 2176 0 1 570
box -9 -3 26 105
use INVX2  INVX2_134
timestamp 1713400504
transform 1 0 2136 0 1 570
box -9 -3 26 105
use INVX2  INVX2_135
timestamp 1713400504
transform 1 0 2984 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_136
timestamp 1713400504
transform 1 0 320 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_137
timestamp 1713400504
transform 1 0 424 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_138
timestamp 1713400504
transform 1 0 272 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_139
timestamp 1713400504
transform 1 0 264 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_140
timestamp 1713400504
transform 1 0 288 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_141
timestamp 1713400504
transform 1 0 376 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_142
timestamp 1713400504
transform 1 0 536 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_143
timestamp 1713400504
transform 1 0 584 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_144
timestamp 1713400504
transform 1 0 816 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_145
timestamp 1713400504
transform 1 0 1000 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_146
timestamp 1713400504
transform 1 0 864 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_147
timestamp 1713400504
transform 1 0 736 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_148
timestamp 1713400504
transform 1 0 560 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_149
timestamp 1713400504
transform 1 0 616 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_150
timestamp 1713400504
transform 1 0 488 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_151
timestamp 1713400504
transform 1 0 504 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_152
timestamp 1713400504
transform 1 0 416 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_153
timestamp 1713400504
transform 1 0 440 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_154
timestamp 1713400504
transform 1 0 320 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_155
timestamp 1713400504
transform 1 0 192 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_156
timestamp 1713400504
transform 1 0 240 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_157
timestamp 1713400504
transform 1 0 80 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_158
timestamp 1713400504
transform 1 0 240 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_159
timestamp 1713400504
transform 1 0 224 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_160
timestamp 1713400504
transform 1 0 104 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_161
timestamp 1713400504
transform 1 0 120 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_162
timestamp 1713400504
transform 1 0 136 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_163
timestamp 1713400504
transform 1 0 80 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_164
timestamp 1713400504
transform 1 0 192 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_165
timestamp 1713400504
transform 1 0 96 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_166
timestamp 1713400504
transform 1 0 176 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_167
timestamp 1713400504
transform 1 0 368 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_168
timestamp 1713400504
transform 1 0 288 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_169
timestamp 1713400504
transform 1 0 552 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_170
timestamp 1713400504
transform 1 0 400 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_171
timestamp 1713400504
transform 1 0 352 0 1 570
box -9 -3 26 105
use INVX2  INVX2_172
timestamp 1713400504
transform 1 0 2472 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_173
timestamp 1713400504
transform 1 0 2656 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_174
timestamp 1713400504
transform 1 0 2896 0 1 970
box -9 -3 26 105
use INVX2  INVX2_175
timestamp 1713400504
transform 1 0 2816 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_176
timestamp 1713400504
transform 1 0 2656 0 1 770
box -9 -3 26 105
use INVX2  INVX2_177
timestamp 1713400504
transform 1 0 2720 0 1 970
box -9 -3 26 105
use INVX2  INVX2_178
timestamp 1713400504
transform 1 0 2888 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_179
timestamp 1713400504
transform 1 0 2784 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_180
timestamp 1713400504
transform 1 0 2888 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_181
timestamp 1713400504
transform 1 0 2880 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_182
timestamp 1713400504
transform 1 0 1848 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_183
timestamp 1713400504
transform 1 0 456 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_184
timestamp 1713400504
transform 1 0 592 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_185
timestamp 1713400504
transform 1 0 416 0 1 970
box -9 -3 26 105
use INVX2  INVX2_186
timestamp 1713400504
transform 1 0 216 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_187
timestamp 1713400504
transform 1 0 512 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_188
timestamp 1713400504
transform 1 0 552 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_189
timestamp 1713400504
transform 1 0 248 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_190
timestamp 1713400504
transform 1 0 672 0 1 170
box -9 -3 26 105
use INVX2  INVX2_191
timestamp 1713400504
transform 1 0 504 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_192
timestamp 1713400504
transform 1 0 512 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_193
timestamp 1713400504
transform 1 0 840 0 1 370
box -9 -3 26 105
use INVX2  INVX2_194
timestamp 1713400504
transform 1 0 656 0 1 570
box -9 -3 26 105
use INVX2  INVX2_195
timestamp 1713400504
transform 1 0 224 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_196
timestamp 1713400504
transform 1 0 688 0 1 770
box -9 -3 26 105
use INVX2  INVX2_197
timestamp 1713400504
transform 1 0 744 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_198
timestamp 1713400504
transform 1 0 640 0 1 770
box -9 -3 26 105
use INVX2  INVX2_199
timestamp 1713400504
transform 1 0 880 0 1 570
box -9 -3 26 105
use INVX2  INVX2_200
timestamp 1713400504
transform 1 0 312 0 1 770
box -9 -3 26 105
use INVX2  INVX2_201
timestamp 1713400504
transform 1 0 216 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_202
timestamp 1713400504
transform 1 0 88 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_203
timestamp 1713400504
transform 1 0 240 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_204
timestamp 1713400504
transform 1 0 200 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_205
timestamp 1713400504
transform 1 0 824 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_206
timestamp 1713400504
transform 1 0 688 0 1 170
box -9 -3 26 105
use INVX2  INVX2_207
timestamp 1713400504
transform 1 0 960 0 1 370
box -9 -3 26 105
use INVX2  INVX2_208
timestamp 1713400504
transform 1 0 1160 0 1 170
box -9 -3 26 105
use INVX2  INVX2_209
timestamp 1713400504
transform 1 0 632 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_210
timestamp 1713400504
transform 1 0 648 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_211
timestamp 1713400504
transform 1 0 976 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_212
timestamp 1713400504
transform 1 0 2000 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_213
timestamp 1713400504
transform 1 0 360 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_214
timestamp 1713400504
transform 1 0 2536 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_215
timestamp 1713400504
transform 1 0 288 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_216
timestamp 1713400504
transform 1 0 1272 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_217
timestamp 1713400504
transform 1 0 2096 0 1 570
box -9 -3 26 105
use INVX2  INVX2_218
timestamp 1713400504
transform 1 0 1632 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_219
timestamp 1713400504
transform 1 0 2472 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_220
timestamp 1713400504
transform 1 0 1568 0 1 370
box -9 -3 26 105
use INVX2  INVX2_221
timestamp 1713400504
transform 1 0 2504 0 1 770
box -9 -3 26 105
use INVX2  INVX2_222
timestamp 1713400504
transform 1 0 1584 0 -1 170
box -9 -3 26 105
use M2_M1  M2_M1_0
timestamp 1713400504
transform 1 0 2876 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1
timestamp 1713400504
transform 1 0 2844 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2
timestamp 1713400504
transform 1 0 2948 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3
timestamp 1713400504
transform 1 0 2820 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4
timestamp 1713400504
transform 1 0 2836 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_5
timestamp 1713400504
transform 1 0 2828 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_6
timestamp 1713400504
transform 1 0 2852 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_7
timestamp 1713400504
transform 1 0 2852 0 1 955
box -2 -2 2 2
use M2_M1  M2_M1_8
timestamp 1713400504
transform 1 0 2772 0 1 955
box -2 -2 2 2
use M2_M1  M2_M1_9
timestamp 1713400504
transform 1 0 2772 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_10
timestamp 1713400504
transform 1 0 2908 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_11
timestamp 1713400504
transform 1 0 2796 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_12
timestamp 1713400504
transform 1 0 2956 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_13
timestamp 1713400504
transform 1 0 2956 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_14
timestamp 1713400504
transform 1 0 340 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_15
timestamp 1713400504
transform 1 0 332 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_16
timestamp 1713400504
transform 1 0 468 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_17
timestamp 1713400504
transform 1 0 428 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_18
timestamp 1713400504
transform 1 0 428 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_19
timestamp 1713400504
transform 1 0 300 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_20
timestamp 1713400504
transform 1 0 260 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_21
timestamp 1713400504
transform 1 0 164 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_22
timestamp 1713400504
transform 1 0 164 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_23
timestamp 1713400504
transform 1 0 132 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_24
timestamp 1713400504
transform 1 0 124 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_25
timestamp 1713400504
transform 1 0 172 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_26
timestamp 1713400504
transform 1 0 156 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_27
timestamp 1713400504
transform 1 0 84 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_28
timestamp 1713400504
transform 1 0 84 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_29
timestamp 1713400504
transform 1 0 76 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_30
timestamp 1713400504
transform 1 0 76 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_31
timestamp 1713400504
transform 1 0 452 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_32
timestamp 1713400504
transform 1 0 260 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_33
timestamp 1713400504
transform 1 0 260 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_34
timestamp 1713400504
transform 1 0 252 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_35
timestamp 1713400504
transform 1 0 244 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_36
timestamp 1713400504
transform 1 0 244 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_37
timestamp 1713400504
transform 1 0 956 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_38
timestamp 1713400504
transform 1 0 780 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_39
timestamp 1713400504
transform 1 0 620 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_40
timestamp 1713400504
transform 1 0 468 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_41
timestamp 1713400504
transform 1 0 468 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_42
timestamp 1713400504
transform 1 0 468 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_43
timestamp 1713400504
transform 1 0 980 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_44
timestamp 1713400504
transform 1 0 916 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_45
timestamp 1713400504
transform 1 0 884 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_46
timestamp 1713400504
transform 1 0 756 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_47
timestamp 1713400504
transform 1 0 668 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_48
timestamp 1713400504
transform 1 0 620 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_49
timestamp 1713400504
transform 1 0 2620 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_50
timestamp 1713400504
transform 1 0 2564 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_51
timestamp 1713400504
transform 1 0 2484 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_52
timestamp 1713400504
transform 1 0 2220 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_53
timestamp 1713400504
transform 1 0 2220 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_54
timestamp 1713400504
transform 1 0 2204 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_55
timestamp 1713400504
transform 1 0 2516 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_56
timestamp 1713400504
transform 1 0 2476 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_57
timestamp 1713400504
transform 1 0 2420 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_58
timestamp 1713400504
transform 1 0 2332 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_59
timestamp 1713400504
transform 1 0 2332 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_60
timestamp 1713400504
transform 1 0 2564 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_61
timestamp 1713400504
transform 1 0 2500 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_62
timestamp 1713400504
transform 1 0 2396 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_63
timestamp 1713400504
transform 1 0 2260 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_64
timestamp 1713400504
transform 1 0 2260 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_65
timestamp 1713400504
transform 1 0 2244 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_66
timestamp 1713400504
transform 1 0 2852 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_67
timestamp 1713400504
transform 1 0 2596 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_68
timestamp 1713400504
transform 1 0 2444 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_69
timestamp 1713400504
transform 1 0 2396 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_70
timestamp 1713400504
transform 1 0 204 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_71
timestamp 1713400504
transform 1 0 100 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_72
timestamp 1713400504
transform 1 0 188 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_73
timestamp 1713400504
transform 1 0 188 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_74
timestamp 1713400504
transform 1 0 404 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_75
timestamp 1713400504
transform 1 0 396 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_76
timestamp 1713400504
transform 1 0 628 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_77
timestamp 1713400504
transform 1 0 612 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_78
timestamp 1713400504
transform 1 0 580 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_79
timestamp 1713400504
transform 1 0 556 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_80
timestamp 1713400504
transform 1 0 844 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_81
timestamp 1713400504
transform 1 0 812 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_82
timestamp 1713400504
transform 1 0 756 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_83
timestamp 1713400504
transform 1 0 972 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_84
timestamp 1713400504
transform 1 0 892 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_85
timestamp 1713400504
transform 1 0 1052 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_86
timestamp 1713400504
transform 1 0 964 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_87
timestamp 1713400504
transform 1 0 964 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_88
timestamp 1713400504
transform 1 0 1036 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_89
timestamp 1713400504
transform 1 0 1004 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_90
timestamp 1713400504
transform 1 0 940 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_91
timestamp 1713400504
transform 1 0 868 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_92
timestamp 1713400504
transform 1 0 820 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_93
timestamp 1713400504
transform 1 0 740 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_94
timestamp 1713400504
transform 1 0 700 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_95
timestamp 1713400504
transform 1 0 588 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_96
timestamp 1713400504
transform 1 0 580 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_97
timestamp 1713400504
transform 1 0 564 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_98
timestamp 1713400504
transform 1 0 660 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_99
timestamp 1713400504
transform 1 0 620 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_100
timestamp 1713400504
transform 1 0 812 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_101
timestamp 1713400504
transform 1 0 492 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_102
timestamp 1713400504
transform 1 0 652 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_103
timestamp 1713400504
transform 1 0 508 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_104
timestamp 1713400504
transform 1 0 516 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_105
timestamp 1713400504
transform 1 0 444 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_106
timestamp 1713400504
transform 1 0 500 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_107
timestamp 1713400504
transform 1 0 428 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_108
timestamp 1713400504
transform 1 0 340 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_109
timestamp 1713400504
transform 1 0 324 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_110
timestamp 1713400504
transform 1 0 508 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_111
timestamp 1713400504
transform 1 0 420 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_112
timestamp 1713400504
transform 1 0 284 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_113
timestamp 1713400504
transform 1 0 196 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_114
timestamp 1713400504
transform 1 0 316 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_115
timestamp 1713400504
transform 1 0 244 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_116
timestamp 1713400504
transform 1 0 300 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_117
timestamp 1713400504
transform 1 0 228 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_118
timestamp 1713400504
transform 1 0 276 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_119
timestamp 1713400504
transform 1 0 204 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_120
timestamp 1713400504
transform 1 0 100 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_121
timestamp 1713400504
transform 1 0 84 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_122
timestamp 1713400504
transform 1 0 340 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_123
timestamp 1713400504
transform 1 0 244 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_124
timestamp 1713400504
transform 1 0 116 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_125
timestamp 1713400504
transform 1 0 68 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_126
timestamp 1713400504
transform 1 0 124 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_127
timestamp 1713400504
transform 1 0 116 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_128
timestamp 1713400504
transform 1 0 140 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_129
timestamp 1713400504
transform 1 0 132 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_130
timestamp 1713400504
transform 1 0 172 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_131
timestamp 1713400504
transform 1 0 140 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_132
timestamp 1713400504
transform 1 0 116 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_133
timestamp 1713400504
transform 1 0 84 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_134
timestamp 1713400504
transform 1 0 212 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_135
timestamp 1713400504
transform 1 0 196 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_136
timestamp 1713400504
transform 1 0 244 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_137
timestamp 1713400504
transform 1 0 236 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_138
timestamp 1713400504
transform 1 0 172 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_139
timestamp 1713400504
transform 1 0 100 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_140
timestamp 1713400504
transform 1 0 100 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_141
timestamp 1713400504
transform 1 0 268 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_142
timestamp 1713400504
transform 1 0 268 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_143
timestamp 1713400504
transform 1 0 236 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_144
timestamp 1713400504
transform 1 0 236 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_145
timestamp 1713400504
transform 1 0 196 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_146
timestamp 1713400504
transform 1 0 180 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_147
timestamp 1713400504
transform 1 0 180 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_148
timestamp 1713400504
transform 1 0 340 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_149
timestamp 1713400504
transform 1 0 332 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_150
timestamp 1713400504
transform 1 0 324 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_151
timestamp 1713400504
transform 1 0 316 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_152
timestamp 1713400504
transform 1 0 308 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_153
timestamp 1713400504
transform 1 0 156 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_154
timestamp 1713400504
transform 1 0 356 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_155
timestamp 1713400504
transform 1 0 340 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_156
timestamp 1713400504
transform 1 0 324 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_157
timestamp 1713400504
transform 1 0 324 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_158
timestamp 1713400504
transform 1 0 324 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_159
timestamp 1713400504
transform 1 0 324 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_160
timestamp 1713400504
transform 1 0 620 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_161
timestamp 1713400504
transform 1 0 540 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_162
timestamp 1713400504
transform 1 0 468 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_163
timestamp 1713400504
transform 1 0 428 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_164
timestamp 1713400504
transform 1 0 396 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_165
timestamp 1713400504
transform 1 0 388 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_166
timestamp 1713400504
transform 1 0 380 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_167
timestamp 1713400504
transform 1 0 1412 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_168
timestamp 1713400504
transform 1 0 1356 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_169
timestamp 1713400504
transform 1 0 1332 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_170
timestamp 1713400504
transform 1 0 1332 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_171
timestamp 1713400504
transform 1 0 1316 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_172
timestamp 1713400504
transform 1 0 1252 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_173
timestamp 1713400504
transform 1 0 1252 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_174
timestamp 1713400504
transform 1 0 1196 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_175
timestamp 1713400504
transform 1 0 1196 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_176
timestamp 1713400504
transform 1 0 1124 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_177
timestamp 1713400504
transform 1 0 1084 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_178
timestamp 1713400504
transform 1 0 1084 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_179
timestamp 1713400504
transform 1 0 1036 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_180
timestamp 1713400504
transform 1 0 1020 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_181
timestamp 1713400504
transform 1 0 1948 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_182
timestamp 1713400504
transform 1 0 1948 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_183
timestamp 1713400504
transform 1 0 1948 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_184
timestamp 1713400504
transform 1 0 1916 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_185
timestamp 1713400504
transform 1 0 2340 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_186
timestamp 1713400504
transform 1 0 2260 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_187
timestamp 1713400504
transform 1 0 2196 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_188
timestamp 1713400504
transform 1 0 2092 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_189
timestamp 1713400504
transform 1 0 2028 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_190
timestamp 1713400504
transform 1 0 2020 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_191
timestamp 1713400504
transform 1 0 2012 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_192
timestamp 1713400504
transform 1 0 2004 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_193
timestamp 1713400504
transform 1 0 2268 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_194
timestamp 1713400504
transform 1 0 2236 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_195
timestamp 1713400504
transform 1 0 2228 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_196
timestamp 1713400504
transform 1 0 2124 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_197
timestamp 1713400504
transform 1 0 2356 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_198
timestamp 1713400504
transform 1 0 2268 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_199
timestamp 1713400504
transform 1 0 2236 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_200
timestamp 1713400504
transform 1 0 2236 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_201
timestamp 1713400504
transform 1 0 1980 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_202
timestamp 1713400504
transform 1 0 2340 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_203
timestamp 1713400504
transform 1 0 2252 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_204
timestamp 1713400504
transform 1 0 2252 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_205
timestamp 1713400504
transform 1 0 1964 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_206
timestamp 1713400504
transform 1 0 1964 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_207
timestamp 1713400504
transform 1 0 1964 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_208
timestamp 1713400504
transform 1 0 1924 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_209
timestamp 1713400504
transform 1 0 1924 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_210
timestamp 1713400504
transform 1 0 2260 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_211
timestamp 1713400504
transform 1 0 2260 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_212
timestamp 1713400504
transform 1 0 2156 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_213
timestamp 1713400504
transform 1 0 2012 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_214
timestamp 1713400504
transform 1 0 1932 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_215
timestamp 1713400504
transform 1 0 1892 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_216
timestamp 1713400504
transform 1 0 1884 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_217
timestamp 1713400504
transform 1 0 2308 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_218
timestamp 1713400504
transform 1 0 2300 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_219
timestamp 1713400504
transform 1 0 2284 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_220
timestamp 1713400504
transform 1 0 2220 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_221
timestamp 1713400504
transform 1 0 2140 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_222
timestamp 1713400504
transform 1 0 2076 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_223
timestamp 1713400504
transform 1 0 2020 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_224
timestamp 1713400504
transform 1 0 2020 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_225
timestamp 1713400504
transform 1 0 1980 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_226
timestamp 1713400504
transform 1 0 1900 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_227
timestamp 1713400504
transform 1 0 2060 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_228
timestamp 1713400504
transform 1 0 1980 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_229
timestamp 1713400504
transform 1 0 1924 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_230
timestamp 1713400504
transform 1 0 1924 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_231
timestamp 1713400504
transform 1 0 1916 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_232
timestamp 1713400504
transform 1 0 2020 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_233
timestamp 1713400504
transform 1 0 2004 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_234
timestamp 1713400504
transform 1 0 1964 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_235
timestamp 1713400504
transform 1 0 1956 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_236
timestamp 1713400504
transform 1 0 1932 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_237
timestamp 1713400504
transform 1 0 1900 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_238
timestamp 1713400504
transform 1 0 1892 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_239
timestamp 1713400504
transform 1 0 2180 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_240
timestamp 1713400504
transform 1 0 2124 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_241
timestamp 1713400504
transform 1 0 2068 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_242
timestamp 1713400504
transform 1 0 2044 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_243
timestamp 1713400504
transform 1 0 2036 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_244
timestamp 1713400504
transform 1 0 1396 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_245
timestamp 1713400504
transform 1 0 1372 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_246
timestamp 1713400504
transform 1 0 668 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_247
timestamp 1713400504
transform 1 0 660 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_248
timestamp 1713400504
transform 1 0 660 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_249
timestamp 1713400504
transform 1 0 660 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_250
timestamp 1713400504
transform 1 0 396 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_251
timestamp 1713400504
transform 1 0 356 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_252
timestamp 1713400504
transform 1 0 348 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_253
timestamp 1713400504
transform 1 0 316 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_254
timestamp 1713400504
transform 1 0 476 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_255
timestamp 1713400504
transform 1 0 476 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_256
timestamp 1713400504
transform 1 0 476 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_257
timestamp 1713400504
transform 1 0 348 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_258
timestamp 1713400504
transform 1 0 564 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_259
timestamp 1713400504
transform 1 0 548 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_260
timestamp 1713400504
transform 1 0 532 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_261
timestamp 1713400504
transform 1 0 532 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_262
timestamp 1713400504
transform 1 0 700 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_263
timestamp 1713400504
transform 1 0 668 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_264
timestamp 1713400504
transform 1 0 644 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_265
timestamp 1713400504
transform 1 0 644 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_266
timestamp 1713400504
transform 1 0 596 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_267
timestamp 1713400504
transform 1 0 548 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_268
timestamp 1713400504
transform 1 0 2860 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_269
timestamp 1713400504
transform 1 0 2860 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_270
timestamp 1713400504
transform 1 0 2572 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_271
timestamp 1713400504
transform 1 0 2564 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_272
timestamp 1713400504
transform 1 0 2508 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_273
timestamp 1713400504
transform 1 0 1500 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_274
timestamp 1713400504
transform 1 0 2980 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_275
timestamp 1713400504
transform 1 0 2804 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_276
timestamp 1713400504
transform 1 0 2804 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_277
timestamp 1713400504
transform 1 0 2508 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_278
timestamp 1713400504
transform 1 0 2124 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_279
timestamp 1713400504
transform 1 0 1828 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_280
timestamp 1713400504
transform 1 0 2868 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_281
timestamp 1713400504
transform 1 0 2708 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_282
timestamp 1713400504
transform 1 0 2692 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_283
timestamp 1713400504
transform 1 0 1404 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_284
timestamp 1713400504
transform 1 0 2916 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_285
timestamp 1713400504
transform 1 0 2828 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_286
timestamp 1713400504
transform 1 0 2772 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_287
timestamp 1713400504
transform 1 0 1812 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_288
timestamp 1713400504
transform 1 0 1164 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_289
timestamp 1713400504
transform 1 0 1164 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_290
timestamp 1713400504
transform 1 0 1708 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_291
timestamp 1713400504
transform 1 0 1700 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_292
timestamp 1713400504
transform 1 0 1948 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_293
timestamp 1713400504
transform 1 0 1844 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_294
timestamp 1713400504
transform 1 0 1844 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_295
timestamp 1713400504
transform 1 0 1748 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_296
timestamp 1713400504
transform 1 0 1732 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_297
timestamp 1713400504
transform 1 0 1732 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_298
timestamp 1713400504
transform 1 0 1676 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_299
timestamp 1713400504
transform 1 0 2796 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_300
timestamp 1713400504
transform 1 0 2772 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_301
timestamp 1713400504
transform 1 0 2644 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_302
timestamp 1713400504
transform 1 0 2220 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_303
timestamp 1713400504
transform 1 0 2652 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_304
timestamp 1713400504
transform 1 0 2636 0 1 2835
box -2 -2 2 2
use M2_M1  M2_M1_305
timestamp 1713400504
transform 1 0 2460 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_306
timestamp 1713400504
transform 1 0 1516 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_307
timestamp 1713400504
transform 1 0 1660 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_308
timestamp 1713400504
transform 1 0 1652 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_309
timestamp 1713400504
transform 1 0 1548 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_310
timestamp 1713400504
transform 1 0 1556 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_311
timestamp 1713400504
transform 1 0 1556 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_312
timestamp 1713400504
transform 1 0 1556 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_313
timestamp 1713400504
transform 1 0 1556 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_314
timestamp 1713400504
transform 1 0 1644 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_315
timestamp 1713400504
transform 1 0 1644 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_316
timestamp 1713400504
transform 1 0 1644 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_317
timestamp 1713400504
transform 1 0 1644 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_318
timestamp 1713400504
transform 1 0 1556 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_319
timestamp 1713400504
transform 1 0 1492 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_320
timestamp 1713400504
transform 1 0 1460 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_321
timestamp 1713400504
transform 1 0 1612 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_322
timestamp 1713400504
transform 1 0 1396 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_323
timestamp 1713400504
transform 1 0 1340 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_324
timestamp 1713400504
transform 1 0 1260 0 1 2705
box -2 -2 2 2
use M2_M1  M2_M1_325
timestamp 1713400504
transform 1 0 1252 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_326
timestamp 1713400504
transform 1 0 1548 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_327
timestamp 1713400504
transform 1 0 1468 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_328
timestamp 1713400504
transform 1 0 1436 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_329
timestamp 1713400504
transform 1 0 1412 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_330
timestamp 1713400504
transform 1 0 1348 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_331
timestamp 1713400504
transform 1 0 1348 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_332
timestamp 1713400504
transform 1 0 1284 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_333
timestamp 1713400504
transform 1 0 1236 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_334
timestamp 1713400504
transform 1 0 204 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_335
timestamp 1713400504
transform 1 0 196 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_336
timestamp 1713400504
transform 1 0 196 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_337
timestamp 1713400504
transform 1 0 172 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_338
timestamp 1713400504
transform 1 0 100 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_339
timestamp 1713400504
transform 1 0 380 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_340
timestamp 1713400504
transform 1 0 364 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_341
timestamp 1713400504
transform 1 0 308 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_342
timestamp 1713400504
transform 1 0 284 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_343
timestamp 1713400504
transform 1 0 1492 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_344
timestamp 1713400504
transform 1 0 1476 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_345
timestamp 1713400504
transform 1 0 1452 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_346
timestamp 1713400504
transform 1 0 1452 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_347
timestamp 1713400504
transform 1 0 1212 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_348
timestamp 1713400504
transform 1 0 1188 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_349
timestamp 1713400504
transform 1 0 2428 0 1 2835
box -2 -2 2 2
use M2_M1  M2_M1_350
timestamp 1713400504
transform 1 0 2180 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_351
timestamp 1713400504
transform 1 0 1692 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_352
timestamp 1713400504
transform 1 0 2636 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_353
timestamp 1713400504
transform 1 0 2596 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_354
timestamp 1713400504
transform 1 0 2612 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_355
timestamp 1713400504
transform 1 0 2604 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_356
timestamp 1713400504
transform 1 0 2564 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_357
timestamp 1713400504
transform 1 0 2028 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_358
timestamp 1713400504
transform 1 0 1988 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_359
timestamp 1713400504
transform 1 0 1988 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_360
timestamp 1713400504
transform 1 0 1964 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_361
timestamp 1713400504
transform 1 0 1964 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_362
timestamp 1713400504
transform 1 0 1876 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_363
timestamp 1713400504
transform 1 0 1876 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_364
timestamp 1713400504
transform 1 0 1836 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_365
timestamp 1713400504
transform 1 0 1812 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_366
timestamp 1713400504
transform 1 0 1812 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_367
timestamp 1713400504
transform 1 0 1756 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_368
timestamp 1713400504
transform 1 0 1740 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_369
timestamp 1713400504
transform 1 0 1740 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_370
timestamp 1713400504
transform 1 0 1604 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_371
timestamp 1713400504
transform 1 0 1548 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_372
timestamp 1713400504
transform 1 0 1548 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_373
timestamp 1713400504
transform 1 0 1532 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_374
timestamp 1713400504
transform 1 0 1500 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_375
timestamp 1713400504
transform 1 0 1492 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_376
timestamp 1713400504
transform 1 0 1492 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_377
timestamp 1713400504
transform 1 0 1700 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_378
timestamp 1713400504
transform 1 0 1700 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_379
timestamp 1713400504
transform 1 0 1692 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_380
timestamp 1713400504
transform 1 0 1532 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_381
timestamp 1713400504
transform 1 0 1444 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_382
timestamp 1713400504
transform 1 0 1444 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_383
timestamp 1713400504
transform 1 0 1444 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_384
timestamp 1713400504
transform 1 0 1436 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_385
timestamp 1713400504
transform 1 0 2012 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_386
timestamp 1713400504
transform 1 0 2012 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_387
timestamp 1713400504
transform 1 0 1932 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_388
timestamp 1713400504
transform 1 0 1924 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_389
timestamp 1713400504
transform 1 0 1924 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_390
timestamp 1713400504
transform 1 0 1908 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_391
timestamp 1713400504
transform 1 0 1908 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_392
timestamp 1713400504
transform 1 0 1892 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_393
timestamp 1713400504
transform 1 0 1884 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_394
timestamp 1713400504
transform 1 0 1884 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_395
timestamp 1713400504
transform 1 0 1804 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_396
timestamp 1713400504
transform 1 0 1668 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_397
timestamp 1713400504
transform 1 0 1508 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_398
timestamp 1713400504
transform 1 0 1508 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_399
timestamp 1713400504
transform 1 0 1412 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_400
timestamp 1713400504
transform 1 0 1316 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_401
timestamp 1713400504
transform 1 0 1260 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_402
timestamp 1713400504
transform 1 0 1228 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_403
timestamp 1713400504
transform 1 0 1468 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_404
timestamp 1713400504
transform 1 0 1468 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_405
timestamp 1713400504
transform 1 0 1972 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_406
timestamp 1713400504
transform 1 0 1932 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_407
timestamp 1713400504
transform 1 0 1932 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_408
timestamp 1713400504
transform 1 0 1876 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_409
timestamp 1713400504
transform 1 0 1764 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_410
timestamp 1713400504
transform 1 0 1708 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_411
timestamp 1713400504
transform 1 0 1708 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_412
timestamp 1713400504
transform 1 0 1692 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_413
timestamp 1713400504
transform 1 0 1652 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_414
timestamp 1713400504
transform 1 0 1652 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_415
timestamp 1713400504
transform 1 0 1212 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_416
timestamp 1713400504
transform 1 0 1140 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_417
timestamp 1713400504
transform 1 0 1132 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_418
timestamp 1713400504
transform 1 0 1036 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_419
timestamp 1713400504
transform 1 0 1164 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_420
timestamp 1713400504
transform 1 0 1076 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_421
timestamp 1713400504
transform 1 0 996 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_422
timestamp 1713400504
transform 1 0 996 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_423
timestamp 1713400504
transform 1 0 1220 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_424
timestamp 1713400504
transform 1 0 1220 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_425
timestamp 1713400504
transform 1 0 1004 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_426
timestamp 1713400504
transform 1 0 988 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_427
timestamp 1713400504
transform 1 0 1100 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_428
timestamp 1713400504
transform 1 0 964 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_429
timestamp 1713400504
transform 1 0 780 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_430
timestamp 1713400504
transform 1 0 780 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_431
timestamp 1713400504
transform 1 0 1268 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_432
timestamp 1713400504
transform 1 0 1268 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_433
timestamp 1713400504
transform 1 0 2228 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_434
timestamp 1713400504
transform 1 0 2036 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_435
timestamp 1713400504
transform 1 0 1956 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_436
timestamp 1713400504
transform 1 0 1956 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_437
timestamp 1713400504
transform 1 0 1636 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_438
timestamp 1713400504
transform 1 0 1636 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_439
timestamp 1713400504
transform 1 0 1948 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_440
timestamp 1713400504
transform 1 0 1948 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_441
timestamp 1713400504
transform 1 0 1860 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_442
timestamp 1713400504
transform 1 0 1900 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_443
timestamp 1713400504
transform 1 0 1900 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_444
timestamp 1713400504
transform 1 0 2276 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_445
timestamp 1713400504
transform 1 0 2260 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_446
timestamp 1713400504
transform 1 0 2236 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_447
timestamp 1713400504
transform 1 0 2220 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_448
timestamp 1713400504
transform 1 0 2196 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_449
timestamp 1713400504
transform 1 0 2092 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_450
timestamp 1713400504
transform 1 0 2044 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_451
timestamp 1713400504
transform 1 0 1820 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_452
timestamp 1713400504
transform 1 0 1812 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_453
timestamp 1713400504
transform 1 0 2324 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_454
timestamp 1713400504
transform 1 0 2308 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_455
timestamp 1713400504
transform 1 0 2276 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_456
timestamp 1713400504
transform 1 0 2268 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_457
timestamp 1713400504
transform 1 0 2068 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_458
timestamp 1713400504
transform 1 0 2052 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_459
timestamp 1713400504
transform 1 0 2036 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_460
timestamp 1713400504
transform 1 0 2036 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_461
timestamp 1713400504
transform 1 0 1260 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_462
timestamp 1713400504
transform 1 0 1260 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_463
timestamp 1713400504
transform 1 0 1100 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_464
timestamp 1713400504
transform 1 0 1092 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_465
timestamp 1713400504
transform 1 0 948 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_466
timestamp 1713400504
transform 1 0 948 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_467
timestamp 1713400504
transform 1 0 1076 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_468
timestamp 1713400504
transform 1 0 1036 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_469
timestamp 1713400504
transform 1 0 2284 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_470
timestamp 1713400504
transform 1 0 2228 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_471
timestamp 1713400504
transform 1 0 2156 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_472
timestamp 1713400504
transform 1 0 2100 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_473
timestamp 1713400504
transform 1 0 1932 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_474
timestamp 1713400504
transform 1 0 1916 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_475
timestamp 1713400504
transform 1 0 1876 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_476
timestamp 1713400504
transform 1 0 2116 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_477
timestamp 1713400504
transform 1 0 2116 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_478
timestamp 1713400504
transform 1 0 2060 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_479
timestamp 1713400504
transform 1 0 2036 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_480
timestamp 1713400504
transform 1 0 2180 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_481
timestamp 1713400504
transform 1 0 2124 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_482
timestamp 1713400504
transform 1 0 2004 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_483
timestamp 1713400504
transform 1 0 1980 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_484
timestamp 1713400504
transform 1 0 1948 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_485
timestamp 1713400504
transform 1 0 1684 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_486
timestamp 1713400504
transform 1 0 1644 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_487
timestamp 1713400504
transform 1 0 2444 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_488
timestamp 1713400504
transform 1 0 2444 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_489
timestamp 1713400504
transform 1 0 1932 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_490
timestamp 1713400504
transform 1 0 1924 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_491
timestamp 1713400504
transform 1 0 1908 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_492
timestamp 1713400504
transform 1 0 1764 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_493
timestamp 1713400504
transform 1 0 1540 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_494
timestamp 1713400504
transform 1 0 1804 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_495
timestamp 1713400504
transform 1 0 1804 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_496
timestamp 1713400504
transform 1 0 1628 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_497
timestamp 1713400504
transform 1 0 1612 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_498
timestamp 1713400504
transform 1 0 2116 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_499
timestamp 1713400504
transform 1 0 1604 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_500
timestamp 1713400504
transform 1 0 1500 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_501
timestamp 1713400504
transform 1 0 1556 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_502
timestamp 1713400504
transform 1 0 1396 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_503
timestamp 1713400504
transform 1 0 1316 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_504
timestamp 1713400504
transform 1 0 1268 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_505
timestamp 1713400504
transform 1 0 1548 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_506
timestamp 1713400504
transform 1 0 1532 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_507
timestamp 1713400504
transform 1 0 1460 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_508
timestamp 1713400504
transform 1 0 1396 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_509
timestamp 1713400504
transform 1 0 1252 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_510
timestamp 1713400504
transform 1 0 1252 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_511
timestamp 1713400504
transform 1 0 1492 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_512
timestamp 1713400504
transform 1 0 1476 0 1 2705
box -2 -2 2 2
use M2_M1  M2_M1_513
timestamp 1713400504
transform 1 0 1444 0 1 2705
box -2 -2 2 2
use M2_M1  M2_M1_514
timestamp 1713400504
transform 1 0 1364 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_515
timestamp 1713400504
transform 1 0 1364 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_516
timestamp 1713400504
transform 1 0 2436 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_517
timestamp 1713400504
transform 1 0 1644 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_518
timestamp 1713400504
transform 1 0 1460 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_519
timestamp 1713400504
transform 1 0 1252 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_520
timestamp 1713400504
transform 1 0 1188 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_521
timestamp 1713400504
transform 1 0 2092 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_522
timestamp 1713400504
transform 1 0 1996 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_523
timestamp 1713400504
transform 1 0 1980 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_524
timestamp 1713400504
transform 1 0 1956 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_525
timestamp 1713400504
transform 1 0 1924 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_526
timestamp 1713400504
transform 1 0 1820 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_527
timestamp 1713400504
transform 1 0 2140 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_528
timestamp 1713400504
transform 1 0 2084 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_529
timestamp 1713400504
transform 1 0 2020 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_530
timestamp 1713400504
transform 1 0 1980 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_531
timestamp 1713400504
transform 1 0 2188 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_532
timestamp 1713400504
transform 1 0 2180 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_533
timestamp 1713400504
transform 1 0 2140 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_534
timestamp 1713400504
transform 1 0 2468 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_535
timestamp 1713400504
transform 1 0 2372 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_536
timestamp 1713400504
transform 1 0 2308 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_537
timestamp 1713400504
transform 1 0 2148 0 1 2835
box -2 -2 2 2
use M2_M1  M2_M1_538
timestamp 1713400504
transform 1 0 2780 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_539
timestamp 1713400504
transform 1 0 2508 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_540
timestamp 1713400504
transform 1 0 2396 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_541
timestamp 1713400504
transform 1 0 2356 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_542
timestamp 1713400504
transform 1 0 2740 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_543
timestamp 1713400504
transform 1 0 2644 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_544
timestamp 1713400504
transform 1 0 2420 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_545
timestamp 1713400504
transform 1 0 2300 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_546
timestamp 1713400504
transform 1 0 2300 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_547
timestamp 1713400504
transform 1 0 2436 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_548
timestamp 1713400504
transform 1 0 2428 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_549
timestamp 1713400504
transform 1 0 2932 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_550
timestamp 1713400504
transform 1 0 2844 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_551
timestamp 1713400504
transform 1 0 2764 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_552
timestamp 1713400504
transform 1 0 2700 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_553
timestamp 1713400504
transform 1 0 2636 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_554
timestamp 1713400504
transform 1 0 2628 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_555
timestamp 1713400504
transform 1 0 2988 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_556
timestamp 1713400504
transform 1 0 2892 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_557
timestamp 1713400504
transform 1 0 2692 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_558
timestamp 1713400504
transform 1 0 2660 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_559
timestamp 1713400504
transform 1 0 2660 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_560
timestamp 1713400504
transform 1 0 2580 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_561
timestamp 1713400504
transform 1 0 2548 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_562
timestamp 1713400504
transform 1 0 2444 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_563
timestamp 1713400504
transform 1 0 2972 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_564
timestamp 1713400504
transform 1 0 2892 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_565
timestamp 1713400504
transform 1 0 2876 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_566
timestamp 1713400504
transform 1 0 2676 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_567
timestamp 1713400504
transform 1 0 2676 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_568
timestamp 1713400504
transform 1 0 2668 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_569
timestamp 1713400504
transform 1 0 2540 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_570
timestamp 1713400504
transform 1 0 2540 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_571
timestamp 1713400504
transform 1 0 2452 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_572
timestamp 1713400504
transform 1 0 2428 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_573
timestamp 1713400504
transform 1 0 2692 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_574
timestamp 1713400504
transform 1 0 2628 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_575
timestamp 1713400504
transform 1 0 2436 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_576
timestamp 1713400504
transform 1 0 2356 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_577
timestamp 1713400504
transform 1 0 2340 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_578
timestamp 1713400504
transform 1 0 2580 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_579
timestamp 1713400504
transform 1 0 2548 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_580
timestamp 1713400504
transform 1 0 2532 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_581
timestamp 1713400504
transform 1 0 2820 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_582
timestamp 1713400504
transform 1 0 2668 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_583
timestamp 1713400504
transform 1 0 2668 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_584
timestamp 1713400504
transform 1 0 2644 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_585
timestamp 1713400504
transform 1 0 2516 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_586
timestamp 1713400504
transform 1 0 2956 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_587
timestamp 1713400504
transform 1 0 2956 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_588
timestamp 1713400504
transform 1 0 2732 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_589
timestamp 1713400504
transform 1 0 2732 0 1 1855
box -2 -2 2 2
use M2_M1  M2_M1_590
timestamp 1713400504
transform 1 0 2716 0 1 1855
box -2 -2 2 2
use M2_M1  M2_M1_591
timestamp 1713400504
transform 1 0 2716 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_592
timestamp 1713400504
transform 1 0 2956 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_593
timestamp 1713400504
transform 1 0 2956 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_594
timestamp 1713400504
transform 1 0 2900 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_595
timestamp 1713400504
transform 1 0 2780 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_596
timestamp 1713400504
transform 1 0 2724 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_597
timestamp 1713400504
transform 1 0 2724 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_598
timestamp 1713400504
transform 1 0 2692 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_599
timestamp 1713400504
transform 1 0 2412 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_600
timestamp 1713400504
transform 1 0 2412 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_601
timestamp 1713400504
transform 1 0 2828 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_602
timestamp 1713400504
transform 1 0 2708 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_603
timestamp 1713400504
transform 1 0 2684 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_604
timestamp 1713400504
transform 1 0 2300 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_605
timestamp 1713400504
transform 1 0 2300 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_606
timestamp 1713400504
transform 1 0 2284 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_607
timestamp 1713400504
transform 1 0 2188 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_608
timestamp 1713400504
transform 1 0 2148 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_609
timestamp 1713400504
transform 1 0 2412 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_610
timestamp 1713400504
transform 1 0 2380 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_611
timestamp 1713400504
transform 1 0 2332 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_612
timestamp 1713400504
transform 1 0 2332 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_613
timestamp 1713400504
transform 1 0 2452 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_614
timestamp 1713400504
transform 1 0 2452 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_615
timestamp 1713400504
transform 1 0 2436 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_616
timestamp 1713400504
transform 1 0 2436 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_617
timestamp 1713400504
transform 1 0 2396 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_618
timestamp 1713400504
transform 1 0 2396 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_619
timestamp 1713400504
transform 1 0 2484 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_620
timestamp 1713400504
transform 1 0 2484 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_621
timestamp 1713400504
transform 1 0 2380 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_622
timestamp 1713400504
transform 1 0 2380 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_623
timestamp 1713400504
transform 1 0 2028 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_624
timestamp 1713400504
transform 1 0 1852 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_625
timestamp 1713400504
transform 1 0 1380 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_626
timestamp 1713400504
transform 1 0 1596 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_627
timestamp 1713400504
transform 1 0 1580 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_628
timestamp 1713400504
transform 1 0 1500 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_629
timestamp 1713400504
transform 1 0 1452 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_630
timestamp 1713400504
transform 1 0 1260 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_631
timestamp 1713400504
transform 1 0 1260 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_632
timestamp 1713400504
transform 1 0 1244 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_633
timestamp 1713400504
transform 1 0 1228 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_634
timestamp 1713400504
transform 1 0 1340 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_635
timestamp 1713400504
transform 1 0 1340 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_636
timestamp 1713400504
transform 1 0 1180 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_637
timestamp 1713400504
transform 1 0 1180 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_638
timestamp 1713400504
transform 1 0 1180 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_639
timestamp 1713400504
transform 1 0 2140 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_640
timestamp 1713400504
transform 1 0 2124 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_641
timestamp 1713400504
transform 1 0 2516 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_642
timestamp 1713400504
transform 1 0 2436 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_643
timestamp 1713400504
transform 1 0 2436 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_644
timestamp 1713400504
transform 1 0 2748 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_645
timestamp 1713400504
transform 1 0 2716 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_646
timestamp 1713400504
transform 1 0 2668 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_647
timestamp 1713400504
transform 1 0 2660 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_648
timestamp 1713400504
transform 1 0 2644 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_649
timestamp 1713400504
transform 1 0 2924 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_650
timestamp 1713400504
transform 1 0 2892 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_651
timestamp 1713400504
transform 1 0 2852 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_652
timestamp 1713400504
transform 1 0 2836 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_653
timestamp 1713400504
transform 1 0 2788 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_654
timestamp 1713400504
transform 1 0 2764 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_655
timestamp 1713400504
transform 1 0 2900 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_656
timestamp 1713400504
transform 1 0 2900 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_657
timestamp 1713400504
transform 1 0 2868 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_658
timestamp 1713400504
transform 1 0 2868 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_659
timestamp 1713400504
transform 1 0 2868 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_660
timestamp 1713400504
transform 1 0 2852 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_661
timestamp 1713400504
transform 1 0 2964 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_662
timestamp 1713400504
transform 1 0 2884 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_663
timestamp 1713400504
transform 1 0 2852 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_664
timestamp 1713400504
transform 1 0 2836 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_665
timestamp 1713400504
transform 1 0 2836 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_666
timestamp 1713400504
transform 1 0 2596 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_667
timestamp 1713400504
transform 1 0 2588 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_668
timestamp 1713400504
transform 1 0 2580 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_669
timestamp 1713400504
transform 1 0 2700 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_670
timestamp 1713400504
transform 1 0 2668 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_671
timestamp 1713400504
transform 1 0 2612 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_672
timestamp 1713400504
transform 1 0 2580 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_673
timestamp 1713400504
transform 1 0 2580 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_674
timestamp 1713400504
transform 1 0 2860 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_675
timestamp 1713400504
transform 1 0 2796 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_676
timestamp 1713400504
transform 1 0 2620 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_677
timestamp 1713400504
transform 1 0 2596 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_678
timestamp 1713400504
transform 1 0 2940 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_679
timestamp 1713400504
transform 1 0 2900 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_680
timestamp 1713400504
transform 1 0 2900 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_681
timestamp 1713400504
transform 1 0 2980 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_682
timestamp 1713400504
transform 1 0 2876 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_683
timestamp 1713400504
transform 1 0 2876 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_684
timestamp 1713400504
transform 1 0 2844 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_685
timestamp 1713400504
transform 1 0 2860 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_686
timestamp 1713400504
transform 1 0 2860 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_687
timestamp 1713400504
transform 1 0 2740 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_688
timestamp 1713400504
transform 1 0 2676 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_689
timestamp 1713400504
transform 1 0 2812 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_690
timestamp 1713400504
transform 1 0 2772 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_691
timestamp 1713400504
transform 1 0 2676 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_692
timestamp 1713400504
transform 1 0 2660 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_693
timestamp 1713400504
transform 1 0 2564 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_694
timestamp 1713400504
transform 1 0 2540 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_695
timestamp 1713400504
transform 1 0 2972 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_696
timestamp 1713400504
transform 1 0 2820 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_697
timestamp 1713400504
transform 1 0 2788 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_698
timestamp 1713400504
transform 1 0 2716 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_699
timestamp 1713400504
transform 1 0 2700 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_700
timestamp 1713400504
transform 1 0 2404 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_701
timestamp 1713400504
transform 1 0 2300 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_702
timestamp 1713400504
transform 1 0 2260 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_703
timestamp 1713400504
transform 1 0 2244 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_704
timestamp 1713400504
transform 1 0 2164 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_705
timestamp 1713400504
transform 1 0 2156 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_706
timestamp 1713400504
transform 1 0 2124 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_707
timestamp 1713400504
transform 1 0 2124 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_708
timestamp 1713400504
transform 1 0 2124 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_709
timestamp 1713400504
transform 1 0 2716 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_710
timestamp 1713400504
transform 1 0 2700 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_711
timestamp 1713400504
transform 1 0 2700 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_712
timestamp 1713400504
transform 1 0 2220 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_713
timestamp 1713400504
transform 1 0 2076 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_714
timestamp 1713400504
transform 1 0 2068 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_715
timestamp 1713400504
transform 1 0 2412 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_716
timestamp 1713400504
transform 1 0 2404 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_717
timestamp 1713400504
transform 1 0 2316 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_718
timestamp 1713400504
transform 1 0 2300 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_719
timestamp 1713400504
transform 1 0 2876 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_720
timestamp 1713400504
transform 1 0 2860 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_721
timestamp 1713400504
transform 1 0 2724 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_722
timestamp 1713400504
transform 1 0 2676 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_723
timestamp 1713400504
transform 1 0 2660 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_724
timestamp 1713400504
transform 1 0 2636 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_725
timestamp 1713400504
transform 1 0 2636 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_726
timestamp 1713400504
transform 1 0 2932 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_727
timestamp 1713400504
transform 1 0 2908 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_728
timestamp 1713400504
transform 1 0 2916 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_729
timestamp 1713400504
transform 1 0 2916 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_730
timestamp 1713400504
transform 1 0 2876 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_731
timestamp 1713400504
transform 1 0 2828 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_732
timestamp 1713400504
transform 1 0 2828 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_733
timestamp 1713400504
transform 1 0 2748 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_734
timestamp 1713400504
transform 1 0 2676 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_735
timestamp 1713400504
transform 1 0 2676 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_736
timestamp 1713400504
transform 1 0 2204 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_737
timestamp 1713400504
transform 1 0 2108 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_738
timestamp 1713400504
transform 1 0 2108 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_739
timestamp 1713400504
transform 1 0 2076 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_740
timestamp 1713400504
transform 1 0 1980 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_741
timestamp 1713400504
transform 1 0 2164 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_742
timestamp 1713400504
transform 1 0 2116 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_743
timestamp 1713400504
transform 1 0 2332 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_744
timestamp 1713400504
transform 1 0 2052 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_745
timestamp 1713400504
transform 1 0 1924 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_746
timestamp 1713400504
transform 1 0 1820 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_747
timestamp 1713400504
transform 1 0 1444 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_748
timestamp 1713400504
transform 1 0 2228 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_749
timestamp 1713400504
transform 1 0 2228 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_750
timestamp 1713400504
transform 1 0 2156 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_751
timestamp 1713400504
transform 1 0 2148 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_752
timestamp 1713400504
transform 1 0 2196 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_753
timestamp 1713400504
transform 1 0 2172 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_754
timestamp 1713400504
transform 1 0 2148 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_755
timestamp 1713400504
transform 1 0 2948 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_756
timestamp 1713400504
transform 1 0 2932 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_757
timestamp 1713400504
transform 1 0 596 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_758
timestamp 1713400504
transform 1 0 580 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_759
timestamp 1713400504
transform 1 0 524 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_760
timestamp 1713400504
transform 1 0 508 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_761
timestamp 1713400504
transform 1 0 468 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_762
timestamp 1713400504
transform 1 0 452 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_763
timestamp 1713400504
transform 1 0 396 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_764
timestamp 1713400504
transform 1 0 380 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_765
timestamp 1713400504
transform 1 0 348 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_766
timestamp 1713400504
transform 1 0 348 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_767
timestamp 1713400504
transform 1 0 724 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_768
timestamp 1713400504
transform 1 0 684 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_769
timestamp 1713400504
transform 1 0 564 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_770
timestamp 1713400504
transform 1 0 388 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_771
timestamp 1713400504
transform 1 0 364 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_772
timestamp 1713400504
transform 1 0 284 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_773
timestamp 1713400504
transform 1 0 772 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_774
timestamp 1713400504
transform 1 0 716 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_775
timestamp 1713400504
transform 1 0 620 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_776
timestamp 1713400504
transform 1 0 508 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_777
timestamp 1713400504
transform 1 0 356 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_778
timestamp 1713400504
transform 1 0 348 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_779
timestamp 1713400504
transform 1 0 652 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_780
timestamp 1713400504
transform 1 0 604 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_781
timestamp 1713400504
transform 1 0 884 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_782
timestamp 1713400504
transform 1 0 828 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_783
timestamp 1713400504
transform 1 0 764 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_784
timestamp 1713400504
transform 1 0 964 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_785
timestamp 1713400504
transform 1 0 932 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_786
timestamp 1713400504
transform 1 0 844 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_787
timestamp 1713400504
transform 1 0 828 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_788
timestamp 1713400504
transform 1 0 788 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_789
timestamp 1713400504
transform 1 0 724 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_790
timestamp 1713400504
transform 1 0 684 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_791
timestamp 1713400504
transform 1 0 660 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_792
timestamp 1713400504
transform 1 0 628 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_793
timestamp 1713400504
transform 1 0 524 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_794
timestamp 1713400504
transform 1 0 492 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_795
timestamp 1713400504
transform 1 0 612 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_796
timestamp 1713400504
transform 1 0 572 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_797
timestamp 1713400504
transform 1 0 508 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_798
timestamp 1713400504
transform 1 0 476 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_799
timestamp 1713400504
transform 1 0 460 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_800
timestamp 1713400504
transform 1 0 428 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_801
timestamp 1713400504
transform 1 0 508 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_802
timestamp 1713400504
transform 1 0 292 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_803
timestamp 1713400504
transform 1 0 260 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_804
timestamp 1713400504
transform 1 0 420 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_805
timestamp 1713400504
transform 1 0 364 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_806
timestamp 1713400504
transform 1 0 284 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_807
timestamp 1713400504
transform 1 0 252 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_808
timestamp 1713400504
transform 1 0 420 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_809
timestamp 1713400504
transform 1 0 324 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_810
timestamp 1713400504
transform 1 0 292 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_811
timestamp 1713400504
transform 1 0 308 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_812
timestamp 1713400504
transform 1 0 276 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_813
timestamp 1713400504
transform 1 0 180 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_814
timestamp 1713400504
transform 1 0 148 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_815
timestamp 1713400504
transform 1 0 220 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_816
timestamp 1713400504
transform 1 0 124 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_817
timestamp 1713400504
transform 1 0 92 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_818
timestamp 1713400504
transform 1 0 108 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_819
timestamp 1713400504
transform 1 0 100 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_820
timestamp 1713400504
transform 1 0 220 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_821
timestamp 1713400504
transform 1 0 196 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_822
timestamp 1713400504
transform 1 0 180 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_823
timestamp 1713400504
transform 1 0 164 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_824
timestamp 1713400504
transform 1 0 148 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_825
timestamp 1713400504
transform 1 0 220 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_826
timestamp 1713400504
transform 1 0 140 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_827
timestamp 1713400504
transform 1 0 92 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_828
timestamp 1713400504
transform 1 0 92 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_829
timestamp 1713400504
transform 1 0 92 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_830
timestamp 1713400504
transform 1 0 188 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_831
timestamp 1713400504
transform 1 0 124 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_832
timestamp 1713400504
transform 1 0 84 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_833
timestamp 1713400504
transform 1 0 196 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_834
timestamp 1713400504
transform 1 0 156 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_835
timestamp 1713400504
transform 1 0 84 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_836
timestamp 1713400504
transform 1 0 132 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_837
timestamp 1713400504
transform 1 0 108 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_838
timestamp 1713400504
transform 1 0 268 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_839
timestamp 1713400504
transform 1 0 220 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_840
timestamp 1713400504
transform 1 0 204 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_841
timestamp 1713400504
transform 1 0 196 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_842
timestamp 1713400504
transform 1 0 228 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_843
timestamp 1713400504
transform 1 0 148 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_844
timestamp 1713400504
transform 1 0 132 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_845
timestamp 1713400504
transform 1 0 140 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_846
timestamp 1713400504
transform 1 0 132 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_847
timestamp 1713400504
transform 1 0 332 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_848
timestamp 1713400504
transform 1 0 316 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_849
timestamp 1713400504
transform 1 0 372 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_850
timestamp 1713400504
transform 1 0 348 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_851
timestamp 1713400504
transform 1 0 516 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_852
timestamp 1713400504
transform 1 0 508 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_853
timestamp 1713400504
transform 1 0 500 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_854
timestamp 1713400504
transform 1 0 564 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_855
timestamp 1713400504
transform 1 0 468 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_856
timestamp 1713400504
transform 1 0 452 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_857
timestamp 1713400504
transform 1 0 420 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_858
timestamp 1713400504
transform 1 0 404 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_859
timestamp 1713400504
transform 1 0 372 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_860
timestamp 1713400504
transform 1 0 348 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_861
timestamp 1713400504
transform 1 0 340 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_862
timestamp 1713400504
transform 1 0 324 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_863
timestamp 1713400504
transform 1 0 2636 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_864
timestamp 1713400504
transform 1 0 2636 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_865
timestamp 1713400504
transform 1 0 2492 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_866
timestamp 1713400504
transform 1 0 2116 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_867
timestamp 1713400504
transform 1 0 2116 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_868
timestamp 1713400504
transform 1 0 1916 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_869
timestamp 1713400504
transform 1 0 1868 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_870
timestamp 1713400504
transform 1 0 1780 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_871
timestamp 1713400504
transform 1 0 1556 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_872
timestamp 1713400504
transform 1 0 1348 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_873
timestamp 1713400504
transform 1 0 1300 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_874
timestamp 1713400504
transform 1 0 1300 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_875
timestamp 1713400504
transform 1 0 2892 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_876
timestamp 1713400504
transform 1 0 2892 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_877
timestamp 1713400504
transform 1 0 2860 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_878
timestamp 1713400504
transform 1 0 2796 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_879
timestamp 1713400504
transform 1 0 2796 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_880
timestamp 1713400504
transform 1 0 2788 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_881
timestamp 1713400504
transform 1 0 2780 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_882
timestamp 1713400504
transform 1 0 2780 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_883
timestamp 1713400504
transform 1 0 2756 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_884
timestamp 1713400504
transform 1 0 2756 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_885
timestamp 1713400504
transform 1 0 2716 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_886
timestamp 1713400504
transform 1 0 2540 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_887
timestamp 1713400504
transform 1 0 2956 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_888
timestamp 1713400504
transform 1 0 2916 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_889
timestamp 1713400504
transform 1 0 2892 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_890
timestamp 1713400504
transform 1 0 2852 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_891
timestamp 1713400504
transform 1 0 2644 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_892
timestamp 1713400504
transform 1 0 2604 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_893
timestamp 1713400504
transform 1 0 2732 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_894
timestamp 1713400504
transform 1 0 2684 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_895
timestamp 1713400504
transform 1 0 2956 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_896
timestamp 1713400504
transform 1 0 2916 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_897
timestamp 1713400504
transform 1 0 2772 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_898
timestamp 1713400504
transform 1 0 2732 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_899
timestamp 1713400504
transform 1 0 2956 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_900
timestamp 1713400504
transform 1 0 2916 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_901
timestamp 1713400504
transform 1 0 2948 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_902
timestamp 1713400504
transform 1 0 2900 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_903
timestamp 1713400504
transform 1 0 1892 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_904
timestamp 1713400504
transform 1 0 1860 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_905
timestamp 1713400504
transform 1 0 1860 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_906
timestamp 1713400504
transform 1 0 1860 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_907
timestamp 1713400504
transform 1 0 1812 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_908
timestamp 1713400504
transform 1 0 1812 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_909
timestamp 1713400504
transform 1 0 1772 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_910
timestamp 1713400504
transform 1 0 1772 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_911
timestamp 1713400504
transform 1 0 476 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_912
timestamp 1713400504
transform 1 0 476 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_913
timestamp 1713400504
transform 1 0 396 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_914
timestamp 1713400504
transform 1 0 668 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_915
timestamp 1713400504
transform 1 0 668 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_916
timestamp 1713400504
transform 1 0 652 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_917
timestamp 1713400504
transform 1 0 572 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_918
timestamp 1713400504
transform 1 0 484 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_919
timestamp 1713400504
transform 1 0 204 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_920
timestamp 1713400504
transform 1 0 148 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_921
timestamp 1713400504
transform 1 0 148 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_922
timestamp 1713400504
transform 1 0 572 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_923
timestamp 1713400504
transform 1 0 532 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_924
timestamp 1713400504
transform 1 0 532 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_925
timestamp 1713400504
transform 1 0 700 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_926
timestamp 1713400504
transform 1 0 620 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_927
timestamp 1713400504
transform 1 0 236 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_928
timestamp 1713400504
transform 1 0 220 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_929
timestamp 1713400504
transform 1 0 220 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_930
timestamp 1713400504
transform 1 0 748 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_931
timestamp 1713400504
transform 1 0 684 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_932
timestamp 1713400504
transform 1 0 684 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_933
timestamp 1713400504
transform 1 0 620 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_934
timestamp 1713400504
transform 1 0 548 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_935
timestamp 1713400504
transform 1 0 548 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_936
timestamp 1713400504
transform 1 0 620 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_937
timestamp 1713400504
transform 1 0 516 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_938
timestamp 1713400504
transform 1 0 516 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_939
timestamp 1713400504
transform 1 0 908 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_940
timestamp 1713400504
transform 1 0 868 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_941
timestamp 1713400504
transform 1 0 868 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_942
timestamp 1713400504
transform 1 0 620 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_943
timestamp 1713400504
transform 1 0 532 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_944
timestamp 1713400504
transform 1 0 276 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_945
timestamp 1713400504
transform 1 0 204 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_946
timestamp 1713400504
transform 1 0 204 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_947
timestamp 1713400504
transform 1 0 756 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_948
timestamp 1713400504
transform 1 0 756 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_949
timestamp 1713400504
transform 1 0 740 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_950
timestamp 1713400504
transform 1 0 820 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_951
timestamp 1713400504
transform 1 0 820 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_952
timestamp 1713400504
transform 1 0 804 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_953
timestamp 1713400504
transform 1 0 636 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_954
timestamp 1713400504
transform 1 0 636 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_955
timestamp 1713400504
transform 1 0 636 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_956
timestamp 1713400504
transform 1 0 1092 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_957
timestamp 1713400504
transform 1 0 972 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_958
timestamp 1713400504
transform 1 0 284 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_959
timestamp 1713400504
transform 1 0 196 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_960
timestamp 1713400504
transform 1 0 212 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_961
timestamp 1713400504
transform 1 0 204 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_962
timestamp 1713400504
transform 1 0 116 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_963
timestamp 1713400504
transform 1 0 92 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_964
timestamp 1713400504
transform 1 0 92 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_965
timestamp 1713400504
transform 1 0 508 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_966
timestamp 1713400504
transform 1 0 508 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_967
timestamp 1713400504
transform 1 0 364 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_968
timestamp 1713400504
transform 1 0 348 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_969
timestamp 1713400504
transform 1 0 348 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_970
timestamp 1713400504
transform 1 0 260 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_971
timestamp 1713400504
transform 1 0 252 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_972
timestamp 1713400504
transform 1 0 252 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_973
timestamp 1713400504
transform 1 0 180 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_974
timestamp 1713400504
transform 1 0 140 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_975
timestamp 1713400504
transform 1 0 924 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_976
timestamp 1713400504
transform 1 0 924 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_977
timestamp 1713400504
transform 1 0 876 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_978
timestamp 1713400504
transform 1 0 772 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_979
timestamp 1713400504
transform 1 0 756 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_980
timestamp 1713400504
transform 1 0 1148 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_981
timestamp 1713400504
transform 1 0 1036 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_982
timestamp 1713400504
transform 1 0 1124 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_983
timestamp 1713400504
transform 1 0 1124 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_984
timestamp 1713400504
transform 1 0 1092 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_985
timestamp 1713400504
transform 1 0 996 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_986
timestamp 1713400504
transform 1 0 1028 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_987
timestamp 1713400504
transform 1 0 932 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_988
timestamp 1713400504
transform 1 0 644 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_989
timestamp 1713400504
transform 1 0 804 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_990
timestamp 1713400504
transform 1 0 724 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_991
timestamp 1713400504
transform 1 0 2932 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_992
timestamp 1713400504
transform 1 0 2932 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_993
timestamp 1713400504
transform 1 0 2932 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_994
timestamp 1713400504
transform 1 0 2868 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_995
timestamp 1713400504
transform 1 0 2772 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_996
timestamp 1713400504
transform 1 0 2684 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_997
timestamp 1713400504
transform 1 0 2684 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_998
timestamp 1713400504
transform 1 0 2636 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_999
timestamp 1713400504
transform 1 0 2556 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1000
timestamp 1713400504
transform 1 0 2540 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1001
timestamp 1713400504
transform 1 0 2532 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1002
timestamp 1713400504
transform 1 0 2500 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1003
timestamp 1713400504
transform 1 0 2484 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1004
timestamp 1713400504
transform 1 0 2436 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1005
timestamp 1713400504
transform 1 0 2932 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1006
timestamp 1713400504
transform 1 0 2932 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1007
timestamp 1713400504
transform 1 0 2924 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1008
timestamp 1713400504
transform 1 0 2924 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1009
timestamp 1713400504
transform 1 0 2924 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1010
timestamp 1713400504
transform 1 0 2924 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1011
timestamp 1713400504
transform 1 0 2924 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1012
timestamp 1713400504
transform 1 0 2876 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1013
timestamp 1713400504
transform 1 0 2820 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1014
timestamp 1713400504
transform 1 0 2772 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1015
timestamp 1713400504
transform 1 0 2684 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1016
timestamp 1713400504
transform 1 0 2628 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1017
timestamp 1713400504
transform 1 0 2588 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1018
timestamp 1713400504
transform 1 0 2572 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1019
timestamp 1713400504
transform 1 0 2604 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1020
timestamp 1713400504
transform 1 0 2508 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1021
timestamp 1713400504
transform 1 0 2212 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1022
timestamp 1713400504
transform 1 0 2052 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1023
timestamp 1713400504
transform 1 0 1852 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1024
timestamp 1713400504
transform 1 0 1660 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1025
timestamp 1713400504
transform 1 0 1620 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1026
timestamp 1713400504
transform 1 0 1612 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1027
timestamp 1713400504
transform 1 0 1372 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1028
timestamp 1713400504
transform 1 0 1300 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1029
timestamp 1713400504
transform 1 0 1172 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1030
timestamp 1713400504
transform 1 0 1076 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1031
timestamp 1713400504
transform 1 0 1068 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1032
timestamp 1713400504
transform 1 0 980 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1033
timestamp 1713400504
transform 1 0 2780 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1034
timestamp 1713400504
transform 1 0 2780 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1035
timestamp 1713400504
transform 1 0 2764 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1036
timestamp 1713400504
transform 1 0 2732 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1037
timestamp 1713400504
transform 1 0 2724 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1038
timestamp 1713400504
transform 1 0 2556 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1039
timestamp 1713400504
transform 1 0 2460 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1040
timestamp 1713400504
transform 1 0 2412 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1041
timestamp 1713400504
transform 1 0 2412 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1042
timestamp 1713400504
transform 1 0 2220 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1043
timestamp 1713400504
transform 1 0 2220 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1044
timestamp 1713400504
transform 1 0 2212 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1045
timestamp 1713400504
transform 1 0 2212 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1046
timestamp 1713400504
transform 1 0 2164 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1047
timestamp 1713400504
transform 1 0 2324 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1048
timestamp 1713400504
transform 1 0 2228 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1049
timestamp 1713400504
transform 1 0 2180 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1050
timestamp 1713400504
transform 1 0 2084 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1051
timestamp 1713400504
transform 1 0 1996 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1052
timestamp 1713400504
transform 1 0 1996 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1053
timestamp 1713400504
transform 1 0 1812 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1054
timestamp 1713400504
transform 1 0 1716 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1055
timestamp 1713400504
transform 1 0 1708 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1056
timestamp 1713400504
transform 1 0 1564 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1057
timestamp 1713400504
transform 1 0 1548 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1058
timestamp 1713400504
transform 1 0 1516 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1059
timestamp 1713400504
transform 1 0 1468 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1060
timestamp 1713400504
transform 1 0 1444 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1061
timestamp 1713400504
transform 1 0 1988 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1062
timestamp 1713400504
transform 1 0 1876 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1063
timestamp 1713400504
transform 1 0 1852 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1064
timestamp 1713400504
transform 1 0 1708 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1065
timestamp 1713400504
transform 1 0 1652 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1066
timestamp 1713400504
transform 1 0 1580 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1067
timestamp 1713400504
transform 1 0 1140 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1068
timestamp 1713400504
transform 1 0 1068 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1069
timestamp 1713400504
transform 1 0 1044 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1070
timestamp 1713400504
transform 1 0 1036 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1071
timestamp 1713400504
transform 1 0 844 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1072
timestamp 1713400504
transform 1 0 796 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1073
timestamp 1713400504
transform 1 0 724 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1074
timestamp 1713400504
transform 1 0 436 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1075
timestamp 1713400504
transform 1 0 964 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1076
timestamp 1713400504
transform 1 0 940 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1077
timestamp 1713400504
transform 1 0 892 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1078
timestamp 1713400504
transform 1 0 804 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1079
timestamp 1713400504
transform 1 0 716 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1080
timestamp 1713400504
transform 1 0 652 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1081
timestamp 1713400504
transform 1 0 628 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1082
timestamp 1713400504
transform 1 0 612 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1083
timestamp 1713400504
transform 1 0 580 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1084
timestamp 1713400504
transform 1 0 508 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1085
timestamp 1713400504
transform 1 0 476 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1086
timestamp 1713400504
transform 1 0 396 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1087
timestamp 1713400504
transform 1 0 140 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1088
timestamp 1713400504
transform 1 0 92 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1089
timestamp 1713400504
transform 1 0 604 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1090
timestamp 1713400504
transform 1 0 596 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1091
timestamp 1713400504
transform 1 0 468 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1092
timestamp 1713400504
transform 1 0 420 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1093
timestamp 1713400504
transform 1 0 412 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1094
timestamp 1713400504
transform 1 0 388 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1095
timestamp 1713400504
transform 1 0 252 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1096
timestamp 1713400504
transform 1 0 236 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1097
timestamp 1713400504
transform 1 0 92 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1098
timestamp 1713400504
transform 1 0 92 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1099
timestamp 1713400504
transform 1 0 92 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1100
timestamp 1713400504
transform 1 0 84 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1101
timestamp 1713400504
transform 1 0 84 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1102
timestamp 1713400504
transform 1 0 84 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1103
timestamp 1713400504
transform 1 0 2708 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1104
timestamp 1713400504
transform 1 0 2660 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1105
timestamp 1713400504
transform 1 0 2660 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1106
timestamp 1713400504
transform 1 0 2196 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1107
timestamp 1713400504
transform 1 0 2196 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1108
timestamp 1713400504
transform 1 0 2188 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1109
timestamp 1713400504
transform 1 0 2188 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1110
timestamp 1713400504
transform 1 0 2164 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1111
timestamp 1713400504
transform 1 0 756 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1112
timestamp 1713400504
transform 1 0 708 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1113
timestamp 1713400504
transform 1 0 636 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1114
timestamp 1713400504
transform 1 0 612 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1115
timestamp 1713400504
transform 1 0 588 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1116
timestamp 1713400504
transform 1 0 2412 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1117
timestamp 1713400504
transform 1 0 2412 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_1118
timestamp 1713400504
transform 1 0 2396 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1119
timestamp 1713400504
transform 1 0 2388 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1120
timestamp 1713400504
transform 1 0 2380 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1121
timestamp 1713400504
transform 1 0 2380 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1122
timestamp 1713400504
transform 1 0 2380 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_1123
timestamp 1713400504
transform 1 0 2372 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1124
timestamp 1713400504
transform 1 0 2340 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1125
timestamp 1713400504
transform 1 0 2316 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_1126
timestamp 1713400504
transform 1 0 2316 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1127
timestamp 1713400504
transform 1 0 2268 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_1128
timestamp 1713400504
transform 1 0 2252 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_1129
timestamp 1713400504
transform 1 0 2188 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1130
timestamp 1713400504
transform 1 0 2124 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_1131
timestamp 1713400504
transform 1 0 2116 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1132
timestamp 1713400504
transform 1 0 2100 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1133
timestamp 1713400504
transform 1 0 2084 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1134
timestamp 1713400504
transform 1 0 2076 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1135
timestamp 1713400504
transform 1 0 2036 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_1136
timestamp 1713400504
transform 1 0 2004 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1137
timestamp 1713400504
transform 1 0 1940 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_1138
timestamp 1713400504
transform 1 0 1924 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1139
timestamp 1713400504
transform 1 0 1892 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_1140
timestamp 1713400504
transform 1 0 1892 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1141
timestamp 1713400504
transform 1 0 1876 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1142
timestamp 1713400504
transform 1 0 1868 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_1143
timestamp 1713400504
transform 1 0 1860 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1144
timestamp 1713400504
transform 1 0 1844 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1145
timestamp 1713400504
transform 1 0 2716 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1146
timestamp 1713400504
transform 1 0 2716 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1147
timestamp 1713400504
transform 1 0 2700 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1148
timestamp 1713400504
transform 1 0 2684 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1149
timestamp 1713400504
transform 1 0 2668 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1150
timestamp 1713400504
transform 1 0 2668 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1151
timestamp 1713400504
transform 1 0 2508 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1152
timestamp 1713400504
transform 1 0 2436 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1153
timestamp 1713400504
transform 1 0 2364 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1154
timestamp 1713400504
transform 1 0 2364 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1155
timestamp 1713400504
transform 1 0 2316 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1156
timestamp 1713400504
transform 1 0 2316 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1157
timestamp 1713400504
transform 1 0 2308 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1158
timestamp 1713400504
transform 1 0 2236 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1159
timestamp 1713400504
transform 1 0 2116 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1160
timestamp 1713400504
transform 1 0 2084 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1161
timestamp 1713400504
transform 1 0 2052 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1162
timestamp 1713400504
transform 1 0 2044 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1163
timestamp 1713400504
transform 1 0 2036 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1164
timestamp 1713400504
transform 1 0 1908 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_1165
timestamp 1713400504
transform 1 0 1828 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1166
timestamp 1713400504
transform 1 0 1788 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1167
timestamp 1713400504
transform 1 0 1652 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1168
timestamp 1713400504
transform 1 0 1636 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1169
timestamp 1713400504
transform 1 0 1604 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1170
timestamp 1713400504
transform 1 0 1588 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1171
timestamp 1713400504
transform 1 0 1556 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1172
timestamp 1713400504
transform 1 0 1540 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1173
timestamp 1713400504
transform 1 0 1524 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1174
timestamp 1713400504
transform 1 0 2156 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1175
timestamp 1713400504
transform 1 0 2148 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1176
timestamp 1713400504
transform 1 0 2148 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1177
timestamp 1713400504
transform 1 0 1988 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1178
timestamp 1713400504
transform 1 0 1788 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1179
timestamp 1713400504
transform 1 0 1716 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1180
timestamp 1713400504
transform 1 0 1604 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1181
timestamp 1713400504
transform 1 0 1452 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1182
timestamp 1713400504
transform 1 0 1396 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1183
timestamp 1713400504
transform 1 0 1316 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1184
timestamp 1713400504
transform 1 0 1268 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1185
timestamp 1713400504
transform 1 0 1220 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1186
timestamp 1713400504
transform 1 0 1220 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1187
timestamp 1713400504
transform 1 0 2884 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1188
timestamp 1713400504
transform 1 0 2884 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1189
timestamp 1713400504
transform 1 0 2884 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1190
timestamp 1713400504
transform 1 0 2868 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1191
timestamp 1713400504
transform 1 0 2860 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1192
timestamp 1713400504
transform 1 0 2844 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1193
timestamp 1713400504
transform 1 0 2788 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1194
timestamp 1713400504
transform 1 0 2788 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1195
timestamp 1713400504
transform 1 0 2740 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1196
timestamp 1713400504
transform 1 0 2724 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1197
timestamp 1713400504
transform 1 0 2708 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1198
timestamp 1713400504
transform 1 0 2660 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1199
timestamp 1713400504
transform 1 0 2604 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1200
timestamp 1713400504
transform 1 0 2492 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1201
timestamp 1713400504
transform 1 0 2436 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1202
timestamp 1713400504
transform 1 0 2540 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1203
timestamp 1713400504
transform 1 0 2516 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1204
timestamp 1713400504
transform 1 0 2532 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1205
timestamp 1713400504
transform 1 0 2532 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_1206
timestamp 1713400504
transform 1 0 2436 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1207
timestamp 1713400504
transform 1 0 2436 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_1208
timestamp 1713400504
transform 1 0 2428 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1209
timestamp 1713400504
transform 1 0 2908 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1210
timestamp 1713400504
transform 1 0 2820 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1211
timestamp 1713400504
transform 1 0 2772 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1212
timestamp 1713400504
transform 1 0 2732 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1213
timestamp 1713400504
transform 1 0 2484 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1214
timestamp 1713400504
transform 1 0 2460 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1215
timestamp 1713400504
transform 1 0 2180 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1216
timestamp 1713400504
transform 1 0 2172 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1217
timestamp 1713400504
transform 1 0 2108 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1218
timestamp 1713400504
transform 1 0 2012 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1219
timestamp 1713400504
transform 1 0 1812 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1220
timestamp 1713400504
transform 1 0 1756 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1221
timestamp 1713400504
transform 1 0 1676 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1222
timestamp 1713400504
transform 1 0 1476 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1223
timestamp 1713400504
transform 1 0 1436 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1224
timestamp 1713400504
transform 1 0 1356 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1225
timestamp 1713400504
transform 1 0 1308 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1226
timestamp 1713400504
transform 1 0 1244 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1227
timestamp 1713400504
transform 1 0 1244 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1228
timestamp 1713400504
transform 1 0 1788 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1229
timestamp 1713400504
transform 1 0 1732 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1230
timestamp 1713400504
transform 1 0 1732 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1231
timestamp 1713400504
transform 1 0 1716 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1232
timestamp 1713400504
transform 1 0 1652 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1233
timestamp 1713400504
transform 1 0 1652 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1234
timestamp 1713400504
transform 1 0 1612 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1235
timestamp 1713400504
transform 1 0 1612 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1236
timestamp 1713400504
transform 1 0 1604 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_1237
timestamp 1713400504
transform 1 0 1268 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1238
timestamp 1713400504
transform 1 0 1108 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1239
timestamp 1713400504
transform 1 0 1100 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1240
timestamp 1713400504
transform 1 0 1100 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1241
timestamp 1713400504
transform 1 0 1060 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_1242
timestamp 1713400504
transform 1 0 1052 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1243
timestamp 1713400504
transform 1 0 1052 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1244
timestamp 1713400504
transform 1 0 1020 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1245
timestamp 1713400504
transform 1 0 980 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1246
timestamp 1713400504
transform 1 0 980 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1247
timestamp 1713400504
transform 1 0 364 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1248
timestamp 1713400504
transform 1 0 340 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1249
timestamp 1713400504
transform 1 0 308 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1250
timestamp 1713400504
transform 1 0 292 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1251
timestamp 1713400504
transform 1 0 356 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1252
timestamp 1713400504
transform 1 0 324 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1253
timestamp 1713400504
transform 1 0 180 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1254
timestamp 1713400504
transform 1 0 180 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_1255
timestamp 1713400504
transform 1 0 980 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1256
timestamp 1713400504
transform 1 0 964 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1257
timestamp 1713400504
transform 1 0 964 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1258
timestamp 1713400504
transform 1 0 884 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1259
timestamp 1713400504
transform 1 0 884 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1260
timestamp 1713400504
transform 1 0 884 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_1261
timestamp 1713400504
transform 1 0 828 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1262
timestamp 1713400504
transform 1 0 788 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1263
timestamp 1713400504
transform 1 0 700 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1264
timestamp 1713400504
transform 1 0 652 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1265
timestamp 1713400504
transform 1 0 580 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1266
timestamp 1713400504
transform 1 0 540 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1267
timestamp 1713400504
transform 1 0 540 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1268
timestamp 1713400504
transform 1 0 532 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1269
timestamp 1713400504
transform 1 0 508 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1270
timestamp 1713400504
transform 1 0 396 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1271
timestamp 1713400504
transform 1 0 380 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1272
timestamp 1713400504
transform 1 0 380 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_1273
timestamp 1713400504
transform 1 0 340 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1274
timestamp 1713400504
transform 1 0 332 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1275
timestamp 1713400504
transform 1 0 300 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1276
timestamp 1713400504
transform 1 0 268 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1277
timestamp 1713400504
transform 1 0 236 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1278
timestamp 1713400504
transform 1 0 228 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1279
timestamp 1713400504
transform 1 0 180 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1280
timestamp 1713400504
transform 1 0 180 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1281
timestamp 1713400504
transform 1 0 156 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1282
timestamp 1713400504
transform 1 0 1988 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1283
timestamp 1713400504
transform 1 0 1964 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1284
timestamp 1713400504
transform 1 0 1924 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1285
timestamp 1713400504
transform 1 0 1916 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1286
timestamp 1713400504
transform 1 0 1892 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1287
timestamp 1713400504
transform 1 0 1892 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1288
timestamp 1713400504
transform 1 0 1860 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1289
timestamp 1713400504
transform 1 0 1828 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1290
timestamp 1713400504
transform 1 0 1788 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1291
timestamp 1713400504
transform 1 0 1780 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1292
timestamp 1713400504
transform 1 0 3004 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1293
timestamp 1713400504
transform 1 0 2948 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_1294
timestamp 1713400504
transform 1 0 2644 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_1295
timestamp 1713400504
transform 1 0 2596 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_1296
timestamp 1713400504
transform 1 0 2596 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_1297
timestamp 1713400504
transform 1 0 2388 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_1298
timestamp 1713400504
transform 1 0 2084 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1299
timestamp 1713400504
transform 1 0 1980 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_1300
timestamp 1713400504
transform 1 0 940 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1301
timestamp 1713400504
transform 1 0 924 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_1302
timestamp 1713400504
transform 1 0 924 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1303
timestamp 1713400504
transform 1 0 2572 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1304
timestamp 1713400504
transform 1 0 2540 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1305
timestamp 1713400504
transform 1 0 2476 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1306
timestamp 1713400504
transform 1 0 2460 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1307
timestamp 1713400504
transform 1 0 2444 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1308
timestamp 1713400504
transform 1 0 2356 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1309
timestamp 1713400504
transform 1 0 2324 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1310
timestamp 1713400504
transform 1 0 2324 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1311
timestamp 1713400504
transform 1 0 1988 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1312
timestamp 1713400504
transform 1 0 1940 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1313
timestamp 1713400504
transform 1 0 1940 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1314
timestamp 1713400504
transform 1 0 1716 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1315
timestamp 1713400504
transform 1 0 1564 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1316
timestamp 1713400504
transform 1 0 1476 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1317
timestamp 1713400504
transform 1 0 1604 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1318
timestamp 1713400504
transform 1 0 1588 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1319
timestamp 1713400504
transform 1 0 1508 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1320
timestamp 1713400504
transform 1 0 1468 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1321
timestamp 1713400504
transform 1 0 1444 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1322
timestamp 1713400504
transform 1 0 1372 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1323
timestamp 1713400504
transform 1 0 1372 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1324
timestamp 1713400504
transform 1 0 1684 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1325
timestamp 1713400504
transform 1 0 1596 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1326
timestamp 1713400504
transform 1 0 1420 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1327
timestamp 1713400504
transform 1 0 1340 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1328
timestamp 1713400504
transform 1 0 1324 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1329
timestamp 1713400504
transform 1 0 828 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1330
timestamp 1713400504
transform 1 0 796 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1331
timestamp 1713400504
transform 1 0 740 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1332
timestamp 1713400504
transform 1 0 684 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1333
timestamp 1713400504
transform 1 0 684 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1334
timestamp 1713400504
transform 1 0 604 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1335
timestamp 1713400504
transform 1 0 572 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1336
timestamp 1713400504
transform 1 0 300 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1337
timestamp 1713400504
transform 1 0 244 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1338
timestamp 1713400504
transform 1 0 1380 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1339
timestamp 1713400504
transform 1 0 1380 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1340
timestamp 1713400504
transform 1 0 1324 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1341
timestamp 1713400504
transform 1 0 1332 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1342
timestamp 1713400504
transform 1 0 1268 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1343
timestamp 1713400504
transform 1 0 908 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1344
timestamp 1713400504
transform 1 0 908 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1345
timestamp 1713400504
transform 1 0 852 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1346
timestamp 1713400504
transform 1 0 1340 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1347
timestamp 1713400504
transform 1 0 820 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_1348
timestamp 1713400504
transform 1 0 796 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1349
timestamp 1713400504
transform 1 0 788 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1350
timestamp 1713400504
transform 1 0 732 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_1351
timestamp 1713400504
transform 1 0 732 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1352
timestamp 1713400504
transform 1 0 732 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1353
timestamp 1713400504
transform 1 0 708 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1354
timestamp 1713400504
transform 1 0 652 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1355
timestamp 1713400504
transform 1 0 620 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1356
timestamp 1713400504
transform 1 0 596 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_1357
timestamp 1713400504
transform 1 0 596 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1358
timestamp 1713400504
transform 1 0 540 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1359
timestamp 1713400504
transform 1 0 524 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1360
timestamp 1713400504
transform 1 0 524 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_1361
timestamp 1713400504
transform 1 0 484 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_1362
timestamp 1713400504
transform 1 0 484 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1363
timestamp 1713400504
transform 1 0 452 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_1364
timestamp 1713400504
transform 1 0 444 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1365
timestamp 1713400504
transform 1 0 444 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1366
timestamp 1713400504
transform 1 0 396 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1367
timestamp 1713400504
transform 1 0 396 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_1368
timestamp 1713400504
transform 1 0 380 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1369
timestamp 1713400504
transform 1 0 356 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_1370
timestamp 1713400504
transform 1 0 332 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_1371
timestamp 1713400504
transform 1 0 324 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_1372
timestamp 1713400504
transform 1 0 252 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1373
timestamp 1713400504
transform 1 0 1700 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1374
timestamp 1713400504
transform 1 0 1692 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1375
timestamp 1713400504
transform 1 0 1500 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1376
timestamp 1713400504
transform 1 0 1444 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1377
timestamp 1713400504
transform 1 0 1340 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1378
timestamp 1713400504
transform 1 0 1324 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1379
timestamp 1713400504
transform 1 0 1268 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1380
timestamp 1713400504
transform 1 0 1396 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1381
timestamp 1713400504
transform 1 0 1396 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1382
timestamp 1713400504
transform 1 0 796 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1383
timestamp 1713400504
transform 1 0 724 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1384
timestamp 1713400504
transform 1 0 700 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1385
timestamp 1713400504
transform 1 0 676 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1386
timestamp 1713400504
transform 1 0 628 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1387
timestamp 1713400504
transform 1 0 548 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1388
timestamp 1713400504
transform 1 0 532 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1389
timestamp 1713400504
transform 1 0 508 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1390
timestamp 1713400504
transform 1 0 452 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1391
timestamp 1713400504
transform 1 0 380 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1392
timestamp 1713400504
transform 1 0 756 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_1393
timestamp 1713400504
transform 1 0 708 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1394
timestamp 1713400504
transform 1 0 788 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_1395
timestamp 1713400504
transform 1 0 684 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1396
timestamp 1713400504
transform 1 0 820 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1397
timestamp 1713400504
transform 1 0 692 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1398
timestamp 1713400504
transform 1 0 812 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_1399
timestamp 1713400504
transform 1 0 540 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1400
timestamp 1713400504
transform 1 0 644 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1401
timestamp 1713400504
transform 1 0 532 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1402
timestamp 1713400504
transform 1 0 628 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_1403
timestamp 1713400504
transform 1 0 524 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1404
timestamp 1713400504
transform 1 0 516 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1405
timestamp 1713400504
transform 1 0 420 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1406
timestamp 1713400504
transform 1 0 460 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1407
timestamp 1713400504
transform 1 0 388 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1408
timestamp 1713400504
transform 1 0 676 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1409
timestamp 1713400504
transform 1 0 660 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1410
timestamp 1713400504
transform 1 0 732 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1411
timestamp 1713400504
transform 1 0 732 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1412
timestamp 1713400504
transform 1 0 716 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1413
timestamp 1713400504
transform 1 0 668 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1414
timestamp 1713400504
transform 1 0 500 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1415
timestamp 1713400504
transform 1 0 500 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1416
timestamp 1713400504
transform 1 0 692 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1417
timestamp 1713400504
transform 1 0 692 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1418
timestamp 1713400504
transform 1 0 724 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1419
timestamp 1713400504
transform 1 0 708 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1420
timestamp 1713400504
transform 1 0 540 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1421
timestamp 1713400504
transform 1 0 540 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_1422
timestamp 1713400504
transform 1 0 708 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1423
timestamp 1713400504
transform 1 0 700 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1424
timestamp 1713400504
transform 1 0 524 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1425
timestamp 1713400504
transform 1 0 516 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1426
timestamp 1713400504
transform 1 0 468 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1427
timestamp 1713400504
transform 1 0 388 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1428
timestamp 1713400504
transform 1 0 444 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1429
timestamp 1713400504
transform 1 0 436 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1430
timestamp 1713400504
transform 1 0 292 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1431
timestamp 1713400504
transform 1 0 252 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1432
timestamp 1713400504
transform 1 0 188 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1433
timestamp 1713400504
transform 1 0 180 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1434
timestamp 1713400504
transform 1 0 220 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1435
timestamp 1713400504
transform 1 0 180 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1436
timestamp 1713400504
transform 1 0 212 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1437
timestamp 1713400504
transform 1 0 172 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1438
timestamp 1713400504
transform 1 0 252 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1439
timestamp 1713400504
transform 1 0 220 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1440
timestamp 1713400504
transform 1 0 180 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1441
timestamp 1713400504
transform 1 0 180 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1442
timestamp 1713400504
transform 1 0 212 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_1443
timestamp 1713400504
transform 1 0 148 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1444
timestamp 1713400504
transform 1 0 212 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_1445
timestamp 1713400504
transform 1 0 148 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1446
timestamp 1713400504
transform 1 0 340 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1447
timestamp 1713400504
transform 1 0 308 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1448
timestamp 1713400504
transform 1 0 388 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1449
timestamp 1713400504
transform 1 0 300 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1450
timestamp 1713400504
transform 1 0 412 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_1451
timestamp 1713400504
transform 1 0 316 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1452
timestamp 1713400504
transform 1 0 388 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_1453
timestamp 1713400504
transform 1 0 324 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1454
timestamp 1713400504
transform 1 0 548 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1455
timestamp 1713400504
transform 1 0 516 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1456
timestamp 1713400504
transform 1 0 612 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1457
timestamp 1713400504
transform 1 0 516 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1458
timestamp 1713400504
transform 1 0 748 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_1459
timestamp 1713400504
transform 1 0 652 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1460
timestamp 1713400504
transform 1 0 908 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_1461
timestamp 1713400504
transform 1 0 812 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1462
timestamp 1713400504
transform 1 0 716 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1463
timestamp 1713400504
transform 1 0 716 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1464
timestamp 1713400504
transform 1 0 836 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1465
timestamp 1713400504
transform 1 0 820 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1466
timestamp 1713400504
transform 1 0 948 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1467
timestamp 1713400504
transform 1 0 948 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1468
timestamp 1713400504
transform 1 0 1044 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1469
timestamp 1713400504
transform 1 0 1044 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1470
timestamp 1713400504
transform 1 0 660 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1471
timestamp 1713400504
transform 1 0 612 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1472
timestamp 1713400504
transform 1 0 820 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1473
timestamp 1713400504
transform 1 0 716 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_1474
timestamp 1713400504
transform 1 0 916 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1475
timestamp 1713400504
transform 1 0 876 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_1476
timestamp 1713400504
transform 1 0 420 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1477
timestamp 1713400504
transform 1 0 356 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1478
timestamp 1713400504
transform 1 0 372 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_1479
timestamp 1713400504
transform 1 0 332 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1480
timestamp 1713400504
transform 1 0 396 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1481
timestamp 1713400504
transform 1 0 356 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_1482
timestamp 1713400504
transform 1 0 172 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_1483
timestamp 1713400504
transform 1 0 156 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1484
timestamp 1713400504
transform 1 0 180 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_1485
timestamp 1713400504
transform 1 0 156 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1486
timestamp 1713400504
transform 1 0 172 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_1487
timestamp 1713400504
transform 1 0 156 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1488
timestamp 1713400504
transform 1 0 92 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1489
timestamp 1713400504
transform 1 0 92 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1490
timestamp 1713400504
transform 1 0 108 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1491
timestamp 1713400504
transform 1 0 92 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1492
timestamp 1713400504
transform 1 0 116 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1493
timestamp 1713400504
transform 1 0 100 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1494
timestamp 1713400504
transform 1 0 1556 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1495
timestamp 1713400504
transform 1 0 1428 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_1496
timestamp 1713400504
transform 1 0 1428 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1497
timestamp 1713400504
transform 1 0 388 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1498
timestamp 1713400504
transform 1 0 356 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1499
timestamp 1713400504
transform 1 0 324 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1500
timestamp 1713400504
transform 1 0 252 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1501
timestamp 1713400504
transform 1 0 244 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1502
timestamp 1713400504
transform 1 0 332 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_1503
timestamp 1713400504
transform 1 0 268 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1504
timestamp 1713400504
transform 1 0 268 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1505
timestamp 1713400504
transform 1 0 220 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1506
timestamp 1713400504
transform 1 0 212 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1507
timestamp 1713400504
transform 1 0 188 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1508
timestamp 1713400504
transform 1 0 420 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_1509
timestamp 1713400504
transform 1 0 404 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1510
timestamp 1713400504
transform 1 0 388 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1511
timestamp 1713400504
transform 1 0 356 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1512
timestamp 1713400504
transform 1 0 348 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1513
timestamp 1713400504
transform 1 0 316 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1514
timestamp 1713400504
transform 1 0 604 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1515
timestamp 1713400504
transform 1 0 564 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1516
timestamp 1713400504
transform 1 0 540 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1517
timestamp 1713400504
transform 1 0 484 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1518
timestamp 1713400504
transform 1 0 460 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1519
timestamp 1713400504
transform 1 0 708 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1520
timestamp 1713400504
transform 1 0 628 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1521
timestamp 1713400504
transform 1 0 596 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1522
timestamp 1713400504
transform 1 0 588 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1523
timestamp 1713400504
transform 1 0 732 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1524
timestamp 1713400504
transform 1 0 732 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1525
timestamp 1713400504
transform 1 0 676 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1526
timestamp 1713400504
transform 1 0 660 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1527
timestamp 1713400504
transform 1 0 820 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1528
timestamp 1713400504
transform 1 0 820 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1529
timestamp 1713400504
transform 1 0 796 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1530
timestamp 1713400504
transform 1 0 940 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1531
timestamp 1713400504
transform 1 0 916 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1532
timestamp 1713400504
transform 1 0 916 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1533
timestamp 1713400504
transform 1 0 1012 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1534
timestamp 1713400504
transform 1 0 996 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1535
timestamp 1713400504
transform 1 0 932 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1536
timestamp 1713400504
transform 1 0 900 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1537
timestamp 1713400504
transform 1 0 844 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1538
timestamp 1713400504
transform 1 0 868 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1539
timestamp 1713400504
transform 1 0 844 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1540
timestamp 1713400504
transform 1 0 812 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_1541
timestamp 1713400504
transform 1 0 788 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_1542
timestamp 1713400504
transform 1 0 756 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1543
timestamp 1713400504
transform 1 0 732 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1544
timestamp 1713400504
transform 1 0 652 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1545
timestamp 1713400504
transform 1 0 636 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_1546
timestamp 1713400504
transform 1 0 620 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1547
timestamp 1713400504
transform 1 0 620 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_1548
timestamp 1713400504
transform 1 0 516 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1549
timestamp 1713400504
transform 1 0 484 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1550
timestamp 1713400504
transform 1 0 476 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_1551
timestamp 1713400504
transform 1 0 316 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1552
timestamp 1713400504
transform 1 0 492 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1553
timestamp 1713400504
transform 1 0 228 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1554
timestamp 1713400504
transform 1 0 348 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1555
timestamp 1713400504
transform 1 0 340 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1556
timestamp 1713400504
transform 1 0 284 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1557
timestamp 1713400504
transform 1 0 1660 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_1558
timestamp 1713400504
transform 1 0 1652 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1559
timestamp 1713400504
transform 1 0 1684 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_1560
timestamp 1713400504
transform 1 0 1276 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1561
timestamp 1713400504
transform 1 0 940 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1562
timestamp 1713400504
transform 1 0 1476 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_1563
timestamp 1713400504
transform 1 0 1044 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1564
timestamp 1713400504
transform 1 0 932 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1565
timestamp 1713400504
transform 1 0 740 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1566
timestamp 1713400504
transform 1 0 732 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1567
timestamp 1713400504
transform 1 0 524 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1568
timestamp 1713400504
transform 1 0 492 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1569
timestamp 1713400504
transform 1 0 364 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1570
timestamp 1713400504
transform 1 0 276 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1571
timestamp 1713400504
transform 1 0 212 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1572
timestamp 1713400504
transform 1 0 204 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1573
timestamp 1713400504
transform 1 0 164 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1574
timestamp 1713400504
transform 1 0 124 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1575
timestamp 1713400504
transform 1 0 180 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_1576
timestamp 1713400504
transform 1 0 156 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1577
timestamp 1713400504
transform 1 0 284 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1578
timestamp 1713400504
transform 1 0 220 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1579
timestamp 1713400504
transform 1 0 260 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1580
timestamp 1713400504
transform 1 0 260 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1581
timestamp 1713400504
transform 1 0 492 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1582
timestamp 1713400504
transform 1 0 420 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1583
timestamp 1713400504
transform 1 0 380 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_1584
timestamp 1713400504
transform 1 0 268 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1585
timestamp 1713400504
transform 1 0 244 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1586
timestamp 1713400504
transform 1 0 620 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1587
timestamp 1713400504
transform 1 0 612 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1588
timestamp 1713400504
transform 1 0 572 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1589
timestamp 1713400504
transform 1 0 548 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_1590
timestamp 1713400504
transform 1 0 548 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1591
timestamp 1713400504
transform 1 0 540 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1592
timestamp 1713400504
transform 1 0 676 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1593
timestamp 1713400504
transform 1 0 676 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1594
timestamp 1713400504
transform 1 0 660 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1595
timestamp 1713400504
transform 1 0 556 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1596
timestamp 1713400504
transform 1 0 460 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1597
timestamp 1713400504
transform 1 0 436 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1598
timestamp 1713400504
transform 1 0 300 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1599
timestamp 1713400504
transform 1 0 300 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1600
timestamp 1713400504
transform 1 0 692 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1601
timestamp 1713400504
transform 1 0 676 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1602
timestamp 1713400504
transform 1 0 500 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1603
timestamp 1713400504
transform 1 0 444 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1604
timestamp 1713400504
transform 1 0 844 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_1605
timestamp 1713400504
transform 1 0 820 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1606
timestamp 1713400504
transform 1 0 660 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1607
timestamp 1713400504
transform 1 0 652 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1608
timestamp 1713400504
transform 1 0 740 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1609
timestamp 1713400504
transform 1 0 620 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1610
timestamp 1713400504
transform 1 0 596 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1611
timestamp 1713400504
transform 1 0 460 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1612
timestamp 1713400504
transform 1 0 372 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1613
timestamp 1713400504
transform 1 0 340 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1614
timestamp 1713400504
transform 1 0 900 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1615
timestamp 1713400504
transform 1 0 876 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1616
timestamp 1713400504
transform 1 0 980 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_1617
timestamp 1713400504
transform 1 0 956 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1618
timestamp 1713400504
transform 1 0 812 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1619
timestamp 1713400504
transform 1 0 684 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1620
timestamp 1713400504
transform 1 0 772 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1621
timestamp 1713400504
transform 1 0 764 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1622
timestamp 1713400504
transform 1 0 724 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1623
timestamp 1713400504
transform 1 0 700 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1624
timestamp 1713400504
transform 1 0 652 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1625
timestamp 1713400504
transform 1 0 628 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1626
timestamp 1713400504
transform 1 0 540 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1627
timestamp 1713400504
transform 1 0 348 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1628
timestamp 1713400504
transform 1 0 348 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1629
timestamp 1713400504
transform 1 0 516 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_1630
timestamp 1713400504
transform 1 0 452 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1631
timestamp 1713400504
transform 1 0 268 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1632
timestamp 1713400504
transform 1 0 156 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1633
timestamp 1713400504
transform 1 0 844 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_1634
timestamp 1713400504
transform 1 0 764 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1635
timestamp 1713400504
transform 1 0 716 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1636
timestamp 1713400504
transform 1 0 692 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1637
timestamp 1713400504
transform 1 0 428 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1638
timestamp 1713400504
transform 1 0 396 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1639
timestamp 1713400504
transform 1 0 444 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1640
timestamp 1713400504
transform 1 0 388 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1641
timestamp 1713400504
transform 1 0 364 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_1642
timestamp 1713400504
transform 1 0 356 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1643
timestamp 1713400504
transform 1 0 564 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1644
timestamp 1713400504
transform 1 0 564 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1645
timestamp 1713400504
transform 1 0 484 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1646
timestamp 1713400504
transform 1 0 484 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1647
timestamp 1713400504
transform 1 0 708 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1648
timestamp 1713400504
transform 1 0 524 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_1649
timestamp 1713400504
transform 1 0 524 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1650
timestamp 1713400504
transform 1 0 484 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1651
timestamp 1713400504
transform 1 0 468 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1652
timestamp 1713400504
transform 1 0 900 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1653
timestamp 1713400504
transform 1 0 900 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1654
timestamp 1713400504
transform 1 0 812 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1655
timestamp 1713400504
transform 1 0 764 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1656
timestamp 1713400504
transform 1 0 748 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1657
timestamp 1713400504
transform 1 0 748 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1658
timestamp 1713400504
transform 1 0 620 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1659
timestamp 1713400504
transform 1 0 612 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1660
timestamp 1713400504
transform 1 0 668 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_1661
timestamp 1713400504
transform 1 0 644 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1662
timestamp 1713400504
transform 1 0 628 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1663
timestamp 1713400504
transform 1 0 572 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1664
timestamp 1713400504
transform 1 0 932 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1665
timestamp 1713400504
transform 1 0 804 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1666
timestamp 1713400504
transform 1 0 564 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1667
timestamp 1713400504
transform 1 0 556 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1668
timestamp 1713400504
transform 1 0 548 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1669
timestamp 1713400504
transform 1 0 220 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1670
timestamp 1713400504
transform 1 0 1164 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1671
timestamp 1713400504
transform 1 0 804 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1672
timestamp 1713400504
transform 1 0 756 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_1673
timestamp 1713400504
transform 1 0 732 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1674
timestamp 1713400504
transform 1 0 572 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1675
timestamp 1713400504
transform 1 0 548 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1676
timestamp 1713400504
transform 1 0 732 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1677
timestamp 1713400504
transform 1 0 660 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1678
timestamp 1713400504
transform 1 0 676 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1679
timestamp 1713400504
transform 1 0 580 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1680
timestamp 1713400504
transform 1 0 412 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1681
timestamp 1713400504
transform 1 0 412 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1682
timestamp 1713400504
transform 1 0 324 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1683
timestamp 1713400504
transform 1 0 228 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1684
timestamp 1713400504
transform 1 0 356 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1685
timestamp 1713400504
transform 1 0 348 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1686
timestamp 1713400504
transform 1 0 324 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1687
timestamp 1713400504
transform 1 0 308 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1688
timestamp 1713400504
transform 1 0 308 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1689
timestamp 1713400504
transform 1 0 348 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_1690
timestamp 1713400504
transform 1 0 276 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_1691
timestamp 1713400504
transform 1 0 268 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1692
timestamp 1713400504
transform 1 0 444 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1693
timestamp 1713400504
transform 1 0 316 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1694
timestamp 1713400504
transform 1 0 364 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1695
timestamp 1713400504
transform 1 0 220 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1696
timestamp 1713400504
transform 1 0 372 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1697
timestamp 1713400504
transform 1 0 348 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1698
timestamp 1713400504
transform 1 0 348 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1699
timestamp 1713400504
transform 1 0 204 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1700
timestamp 1713400504
transform 1 0 652 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1701
timestamp 1713400504
transform 1 0 452 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1702
timestamp 1713400504
transform 1 0 436 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1703
timestamp 1713400504
transform 1 0 420 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1704
timestamp 1713400504
transform 1 0 372 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1705
timestamp 1713400504
transform 1 0 356 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_1706
timestamp 1713400504
transform 1 0 292 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_1707
timestamp 1713400504
transform 1 0 268 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1708
timestamp 1713400504
transform 1 0 332 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1709
timestamp 1713400504
transform 1 0 244 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1710
timestamp 1713400504
transform 1 0 372 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_1711
timestamp 1713400504
transform 1 0 364 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1712
timestamp 1713400504
transform 1 0 212 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_1713
timestamp 1713400504
transform 1 0 212 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1714
timestamp 1713400504
transform 1 0 276 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1715
timestamp 1713400504
transform 1 0 204 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1716
timestamp 1713400504
transform 1 0 556 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1717
timestamp 1713400504
transform 1 0 532 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1718
timestamp 1713400504
transform 1 0 364 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1719
timestamp 1713400504
transform 1 0 356 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1720
timestamp 1713400504
transform 1 0 244 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1721
timestamp 1713400504
transform 1 0 244 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1722
timestamp 1713400504
transform 1 0 196 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1723
timestamp 1713400504
transform 1 0 196 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1724
timestamp 1713400504
transform 1 0 164 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1725
timestamp 1713400504
transform 1 0 316 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1726
timestamp 1713400504
transform 1 0 292 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1727
timestamp 1713400504
transform 1 0 380 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_1728
timestamp 1713400504
transform 1 0 348 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_1729
timestamp 1713400504
transform 1 0 252 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_1730
timestamp 1713400504
transform 1 0 172 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1731
timestamp 1713400504
transform 1 0 92 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1732
timestamp 1713400504
transform 1 0 188 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_1733
timestamp 1713400504
transform 1 0 172 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_1734
timestamp 1713400504
transform 1 0 1508 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1735
timestamp 1713400504
transform 1 0 1404 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_1736
timestamp 1713400504
transform 1 0 1324 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1737
timestamp 1713400504
transform 1 0 884 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1738
timestamp 1713400504
transform 1 0 380 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_1739
timestamp 1713400504
transform 1 0 428 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1740
timestamp 1713400504
transform 1 0 356 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_1741
timestamp 1713400504
transform 1 0 372 0 1 105
box -2 -2 2 2
use M2_M1  M2_M1_1742
timestamp 1713400504
transform 1 0 276 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1743
timestamp 1713400504
transform 1 0 1740 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1744
timestamp 1713400504
transform 1 0 1692 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1745
timestamp 1713400504
transform 1 0 188 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1746
timestamp 1713400504
transform 1 0 188 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1747
timestamp 1713400504
transform 1 0 716 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1748
timestamp 1713400504
transform 1 0 628 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1749
timestamp 1713400504
transform 1 0 572 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1750
timestamp 1713400504
transform 1 0 524 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1751
timestamp 1713400504
transform 1 0 844 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1752
timestamp 1713400504
transform 1 0 764 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1753
timestamp 1713400504
transform 1 0 916 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1754
timestamp 1713400504
transform 1 0 916 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1755
timestamp 1713400504
transform 1 0 1060 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1756
timestamp 1713400504
transform 1 0 1020 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1757
timestamp 1713400504
transform 1 0 844 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1758
timestamp 1713400504
transform 1 0 844 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1759
timestamp 1713400504
transform 1 0 420 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1760
timestamp 1713400504
transform 1 0 420 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1761
timestamp 1713400504
transform 1 0 556 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1762
timestamp 1713400504
transform 1 0 548 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1763
timestamp 1713400504
transform 1 0 556 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1764
timestamp 1713400504
transform 1 0 460 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1765
timestamp 1713400504
transform 1 0 964 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1766
timestamp 1713400504
transform 1 0 924 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1767
timestamp 1713400504
transform 1 0 668 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1768
timestamp 1713400504
transform 1 0 660 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1769
timestamp 1713400504
transform 1 0 1004 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1770
timestamp 1713400504
transform 1 0 1004 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1771
timestamp 1713400504
transform 1 0 1068 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1772
timestamp 1713400504
transform 1 0 1068 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1773
timestamp 1713400504
transform 1 0 1164 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1774
timestamp 1713400504
transform 1 0 1060 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1775
timestamp 1713400504
transform 1 0 836 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1776
timestamp 1713400504
transform 1 0 772 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1777
timestamp 1713400504
transform 1 0 652 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1778
timestamp 1713400504
transform 1 0 652 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1779
timestamp 1713400504
transform 1 0 556 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1780
timestamp 1713400504
transform 1 0 468 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1781
timestamp 1713400504
transform 1 0 228 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1782
timestamp 1713400504
transform 1 0 140 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1783
timestamp 1713400504
transform 1 0 220 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1784
timestamp 1713400504
transform 1 0 132 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1785
timestamp 1713400504
transform 1 0 140 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1786
timestamp 1713400504
transform 1 0 132 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1787
timestamp 1713400504
transform 1 0 1092 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1788
timestamp 1713400504
transform 1 0 1004 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1789
timestamp 1713400504
transform 1 0 868 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1790
timestamp 1713400504
transform 1 0 780 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1791
timestamp 1713400504
transform 1 0 508 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1792
timestamp 1713400504
transform 1 0 508 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1793
timestamp 1713400504
transform 1 0 292 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1794
timestamp 1713400504
transform 1 0 292 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1795
timestamp 1713400504
transform 1 0 204 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1796
timestamp 1713400504
transform 1 0 132 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1797
timestamp 1713400504
transform 1 0 284 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1798
timestamp 1713400504
transform 1 0 284 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1799
timestamp 1713400504
transform 1 0 620 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1800
timestamp 1713400504
transform 1 0 556 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1801
timestamp 1713400504
transform 1 0 412 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1802
timestamp 1713400504
transform 1 0 372 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1803
timestamp 1713400504
transform 1 0 460 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1804
timestamp 1713400504
transform 1 0 380 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1805
timestamp 1713400504
transform 1 0 116 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1806
timestamp 1713400504
transform 1 0 116 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1807
timestamp 1713400504
transform 1 0 172 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1808
timestamp 1713400504
transform 1 0 140 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1809
timestamp 1713400504
transform 1 0 1500 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1810
timestamp 1713400504
transform 1 0 1420 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1811
timestamp 1713400504
transform 1 0 2140 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1812
timestamp 1713400504
transform 1 0 2140 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1813
timestamp 1713400504
transform 1 0 2364 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1814
timestamp 1713400504
transform 1 0 2292 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1815
timestamp 1713400504
transform 1 0 2300 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1816
timestamp 1713400504
transform 1 0 2276 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1817
timestamp 1713400504
transform 1 0 2340 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1818
timestamp 1713400504
transform 1 0 2292 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1819
timestamp 1713400504
transform 1 0 2316 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1820
timestamp 1713400504
transform 1 0 2292 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1821
timestamp 1713400504
transform 1 0 2340 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1822
timestamp 1713400504
transform 1 0 2324 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1823
timestamp 1713400504
transform 1 0 2228 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1824
timestamp 1713400504
transform 1 0 2228 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1825
timestamp 1713400504
transform 1 0 2300 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1826
timestamp 1713400504
transform 1 0 2300 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1827
timestamp 1713400504
transform 1 0 2308 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1828
timestamp 1713400504
transform 1 0 2300 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1829
timestamp 1713400504
transform 1 0 2180 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1830
timestamp 1713400504
transform 1 0 2180 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_1831
timestamp 1713400504
transform 1 0 2116 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1832
timestamp 1713400504
transform 1 0 2108 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1833
timestamp 1713400504
transform 1 0 2060 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1834
timestamp 1713400504
transform 1 0 2060 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1835
timestamp 1713400504
transform 1 0 1972 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1836
timestamp 1713400504
transform 1 0 1844 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1837
timestamp 1713400504
transform 1 0 1948 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1838
timestamp 1713400504
transform 1 0 1876 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1839
timestamp 1713400504
transform 1 0 1972 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1840
timestamp 1713400504
transform 1 0 1924 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1841
timestamp 1713400504
transform 1 0 1852 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1842
timestamp 1713400504
transform 1 0 1820 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1843
timestamp 1713400504
transform 1 0 1908 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1844
timestamp 1713400504
transform 1 0 1908 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1845
timestamp 1713400504
transform 1 0 1860 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1846
timestamp 1713400504
transform 1 0 1844 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1847
timestamp 1713400504
transform 1 0 2004 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1848
timestamp 1713400504
transform 1 0 1988 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1849
timestamp 1713400504
transform 1 0 1876 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1850
timestamp 1713400504
transform 1 0 1860 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1851
timestamp 1713400504
transform 1 0 1988 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1852
timestamp 1713400504
transform 1 0 1988 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1853
timestamp 1713400504
transform 1 0 1244 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1854
timestamp 1713400504
transform 1 0 1076 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_1855
timestamp 1713400504
transform 1 0 996 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1856
timestamp 1713400504
transform 1 0 980 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1857
timestamp 1713400504
transform 1 0 1300 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1858
timestamp 1713400504
transform 1 0 1244 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1859
timestamp 1713400504
transform 1 0 1188 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1860
timestamp 1713400504
transform 1 0 1076 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_1861
timestamp 1713400504
transform 1 0 1244 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1862
timestamp 1713400504
transform 1 0 1108 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1863
timestamp 1713400504
transform 1 0 1060 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1864
timestamp 1713400504
transform 1 0 1044 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1865
timestamp 1713400504
transform 1 0 1292 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1866
timestamp 1713400504
transform 1 0 1260 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1867
timestamp 1713400504
transform 1 0 1204 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1868
timestamp 1713400504
transform 1 0 868 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1869
timestamp 1713400504
transform 1 0 756 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1870
timestamp 1713400504
transform 1 0 740 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1871
timestamp 1713400504
transform 1 0 1356 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1872
timestamp 1713400504
transform 1 0 1300 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1873
timestamp 1713400504
transform 1 0 1292 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1874
timestamp 1713400504
transform 1 0 1260 0 1 1585
box -2 -2 2 2
use M2_M1  M2_M1_1875
timestamp 1713400504
transform 1 0 1252 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_1876
timestamp 1713400504
transform 1 0 1556 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1877
timestamp 1713400504
transform 1 0 1452 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1878
timestamp 1713400504
transform 1 0 1420 0 1 555
box -2 -2 2 2
use M2_M1  M2_M1_1879
timestamp 1713400504
transform 1 0 1412 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_1880
timestamp 1713400504
transform 1 0 1244 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1881
timestamp 1713400504
transform 1 0 1156 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_1882
timestamp 1713400504
transform 1 0 932 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1883
timestamp 1713400504
transform 1 0 892 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1884
timestamp 1713400504
transform 1 0 892 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1885
timestamp 1713400504
transform 1 0 1316 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1886
timestamp 1713400504
transform 1 0 1308 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1887
timestamp 1713400504
transform 1 0 1196 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_1888
timestamp 1713400504
transform 1 0 1188 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1889
timestamp 1713400504
transform 1 0 2012 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1890
timestamp 1713400504
transform 1 0 1956 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1891
timestamp 1713400504
transform 1 0 2204 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1892
timestamp 1713400504
transform 1 0 2100 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1893
timestamp 1713400504
transform 1 0 1964 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1894
timestamp 1713400504
transform 1 0 1940 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1895
timestamp 1713400504
transform 1 0 2220 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1896
timestamp 1713400504
transform 1 0 2212 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1897
timestamp 1713400504
transform 1 0 2196 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1898
timestamp 1713400504
transform 1 0 2164 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1899
timestamp 1713400504
transform 1 0 2140 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1900
timestamp 1713400504
transform 1 0 1884 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1901
timestamp 1713400504
transform 1 0 2180 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1902
timestamp 1713400504
transform 1 0 2172 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1903
timestamp 1713400504
transform 1 0 1924 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1904
timestamp 1713400504
transform 1 0 2364 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1905
timestamp 1713400504
transform 1 0 2260 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1906
timestamp 1713400504
transform 1 0 2428 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1907
timestamp 1713400504
transform 1 0 2396 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1908
timestamp 1713400504
transform 1 0 2444 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1909
timestamp 1713400504
transform 1 0 2340 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1910
timestamp 1713400504
transform 1 0 2380 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1911
timestamp 1713400504
transform 1 0 2356 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1912
timestamp 1713400504
transform 1 0 2268 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1913
timestamp 1713400504
transform 1 0 2236 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1914
timestamp 1713400504
transform 1 0 2380 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1915
timestamp 1713400504
transform 1 0 2324 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1916
timestamp 1713400504
transform 1 0 2876 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_1917
timestamp 1713400504
transform 1 0 2740 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1918
timestamp 1713400504
transform 1 0 2980 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1919
timestamp 1713400504
transform 1 0 2836 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1920
timestamp 1713400504
transform 1 0 2876 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_1921
timestamp 1713400504
transform 1 0 2732 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1922
timestamp 1713400504
transform 1 0 2884 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_1923
timestamp 1713400504
transform 1 0 2756 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1924
timestamp 1713400504
transform 1 0 2828 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_1925
timestamp 1713400504
transform 1 0 2692 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1926
timestamp 1713400504
transform 1 0 2996 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_1927
timestamp 1713400504
transform 1 0 2868 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1928
timestamp 1713400504
transform 1 0 2980 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1929
timestamp 1713400504
transform 1 0 2868 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1930
timestamp 1713400504
transform 1 0 2244 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1931
timestamp 1713400504
transform 1 0 2012 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1932
timestamp 1713400504
transform 1 0 2228 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1933
timestamp 1713400504
transform 1 0 2116 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1934
timestamp 1713400504
transform 1 0 2404 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1935
timestamp 1713400504
transform 1 0 2116 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1936
timestamp 1713400504
transform 1 0 2372 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1937
timestamp 1713400504
transform 1 0 2372 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1938
timestamp 1713400504
transform 1 0 2260 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1939
timestamp 1713400504
transform 1 0 2244 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1940
timestamp 1713400504
transform 1 0 2236 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1941
timestamp 1713400504
transform 1 0 2236 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1942
timestamp 1713400504
transform 1 0 2052 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1943
timestamp 1713400504
transform 1 0 2292 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1944
timestamp 1713400504
transform 1 0 2292 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1945
timestamp 1713400504
transform 1 0 2180 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1946
timestamp 1713400504
transform 1 0 2284 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1947
timestamp 1713400504
transform 1 0 1932 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1948
timestamp 1713400504
transform 1 0 2180 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1949
timestamp 1713400504
transform 1 0 2092 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1950
timestamp 1713400504
transform 1 0 2084 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1951
timestamp 1713400504
transform 1 0 2492 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1952
timestamp 1713400504
transform 1 0 2476 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1953
timestamp 1713400504
transform 1 0 2452 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1954
timestamp 1713400504
transform 1 0 2300 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1955
timestamp 1713400504
transform 1 0 2292 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_1956
timestamp 1713400504
transform 1 0 2972 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1957
timestamp 1713400504
transform 1 0 2948 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1958
timestamp 1713400504
transform 1 0 2924 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1959
timestamp 1713400504
transform 1 0 2868 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1960
timestamp 1713400504
transform 1 0 2812 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1961
timestamp 1713400504
transform 1 0 2740 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_1962
timestamp 1713400504
transform 1 0 2684 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1963
timestamp 1713400504
transform 1 0 2660 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1964
timestamp 1713400504
transform 1 0 2580 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1965
timestamp 1713400504
transform 1 0 2548 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_1966
timestamp 1713400504
transform 1 0 2540 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1967
timestamp 1713400504
transform 1 0 2500 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1968
timestamp 1713400504
transform 1 0 2468 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1969
timestamp 1713400504
transform 1 0 2212 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1970
timestamp 1713400504
transform 1 0 2300 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1971
timestamp 1713400504
transform 1 0 2284 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1972
timestamp 1713400504
transform 1 0 2236 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1973
timestamp 1713400504
transform 1 0 2236 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_1974
timestamp 1713400504
transform 1 0 2204 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_1975
timestamp 1713400504
transform 1 0 2076 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1976
timestamp 1713400504
transform 1 0 2068 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1977
timestamp 1713400504
transform 1 0 2268 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1978
timestamp 1713400504
transform 1 0 2252 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_1979
timestamp 1713400504
transform 1 0 2484 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1980
timestamp 1713400504
transform 1 0 2484 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1981
timestamp 1713400504
transform 1 0 2540 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_1982
timestamp 1713400504
transform 1 0 2452 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1983
timestamp 1713400504
transform 1 0 2436 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1984
timestamp 1713400504
transform 1 0 2604 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1985
timestamp 1713400504
transform 1 0 2508 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_1986
timestamp 1713400504
transform 1 0 2636 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_1987
timestamp 1713400504
transform 1 0 2460 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_1988
timestamp 1713400504
transform 1 0 2460 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1989
timestamp 1713400504
transform 1 0 2356 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1990
timestamp 1713400504
transform 1 0 2324 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1991
timestamp 1713400504
transform 1 0 2460 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1992
timestamp 1713400504
transform 1 0 2436 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1993
timestamp 1713400504
transform 1 0 2396 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1994
timestamp 1713400504
transform 1 0 2348 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1995
timestamp 1713400504
transform 1 0 2444 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1996
timestamp 1713400504
transform 1 0 2348 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1997
timestamp 1713400504
transform 1 0 2460 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_1998
timestamp 1713400504
transform 1 0 2460 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1999
timestamp 1713400504
transform 1 0 2532 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2000
timestamp 1713400504
transform 1 0 2516 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2001
timestamp 1713400504
transform 1 0 2516 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2002
timestamp 1713400504
transform 1 0 2524 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2003
timestamp 1713400504
transform 1 0 2524 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2004
timestamp 1713400504
transform 1 0 2524 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_2005
timestamp 1713400504
transform 1 0 2508 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2006
timestamp 1713400504
transform 1 0 2508 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2007
timestamp 1713400504
transform 1 0 2468 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_2008
timestamp 1713400504
transform 1 0 2468 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2009
timestamp 1713400504
transform 1 0 2332 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2010
timestamp 1713400504
transform 1 0 2420 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2011
timestamp 1713400504
transform 1 0 2380 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2012
timestamp 1713400504
transform 1 0 2428 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2013
timestamp 1713400504
transform 1 0 2340 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2014
timestamp 1713400504
transform 1 0 2404 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2015
timestamp 1713400504
transform 1 0 2404 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2016
timestamp 1713400504
transform 1 0 2364 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_2017
timestamp 1713400504
transform 1 0 2348 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2018
timestamp 1713400504
transform 1 0 2452 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_2019
timestamp 1713400504
transform 1 0 2316 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_2020
timestamp 1713400504
transform 1 0 2316 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_2021
timestamp 1713400504
transform 1 0 2356 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2022
timestamp 1713400504
transform 1 0 2340 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2023
timestamp 1713400504
transform 1 0 2428 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2024
timestamp 1713400504
transform 1 0 2420 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_2025
timestamp 1713400504
transform 1 0 2284 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2026
timestamp 1713400504
transform 1 0 2372 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2027
timestamp 1713400504
transform 1 0 2372 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2028
timestamp 1713400504
transform 1 0 2324 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2029
timestamp 1713400504
transform 1 0 2324 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_2030
timestamp 1713400504
transform 1 0 2412 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2031
timestamp 1713400504
transform 1 0 2396 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2032
timestamp 1713400504
transform 1 0 2340 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2033
timestamp 1713400504
transform 1 0 2132 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2034
timestamp 1713400504
transform 1 0 2436 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_2035
timestamp 1713400504
transform 1 0 2436 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2036
timestamp 1713400504
transform 1 0 2420 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2037
timestamp 1713400504
transform 1 0 2420 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_2038
timestamp 1713400504
transform 1 0 2140 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2039
timestamp 1713400504
transform 1 0 2124 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_2040
timestamp 1713400504
transform 1 0 2732 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2041
timestamp 1713400504
transform 1 0 2716 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2042
timestamp 1713400504
transform 1 0 2300 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2043
timestamp 1713400504
transform 1 0 2196 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2044
timestamp 1713400504
transform 1 0 2332 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2045
timestamp 1713400504
transform 1 0 2308 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2046
timestamp 1713400504
transform 1 0 2684 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2047
timestamp 1713400504
transform 1 0 2348 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_2048
timestamp 1713400504
transform 1 0 2364 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2049
timestamp 1713400504
transform 1 0 2020 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2050
timestamp 1713400504
transform 1 0 2148 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_2051
timestamp 1713400504
transform 1 0 1508 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_2052
timestamp 1713400504
transform 1 0 2172 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_2053
timestamp 1713400504
transform 1 0 2172 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2054
timestamp 1713400504
transform 1 0 2892 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2055
timestamp 1713400504
transform 1 0 2884 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2056
timestamp 1713400504
transform 1 0 2852 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2057
timestamp 1713400504
transform 1 0 2852 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2058
timestamp 1713400504
transform 1 0 2804 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2059
timestamp 1713400504
transform 1 0 2748 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2060
timestamp 1713400504
transform 1 0 2748 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2061
timestamp 1713400504
transform 1 0 2716 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2062
timestamp 1713400504
transform 1 0 2716 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2063
timestamp 1713400504
transform 1 0 2716 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2064
timestamp 1713400504
transform 1 0 2700 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2065
timestamp 1713400504
transform 1 0 2700 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2066
timestamp 1713400504
transform 1 0 2884 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2067
timestamp 1713400504
transform 1 0 2820 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2068
timestamp 1713400504
transform 1 0 2708 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2069
timestamp 1713400504
transform 1 0 2660 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2070
timestamp 1713400504
transform 1 0 2772 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2071
timestamp 1713400504
transform 1 0 2724 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2072
timestamp 1713400504
transform 1 0 2884 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2073
timestamp 1713400504
transform 1 0 2748 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2074
timestamp 1713400504
transform 1 0 2852 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2075
timestamp 1713400504
transform 1 0 2788 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2076
timestamp 1713400504
transform 1 0 2884 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2077
timestamp 1713400504
transform 1 0 2756 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2078
timestamp 1713400504
transform 1 0 2884 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2079
timestamp 1713400504
transform 1 0 2788 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2080
timestamp 1713400504
transform 1 0 2556 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2081
timestamp 1713400504
transform 1 0 2556 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2082
timestamp 1713400504
transform 1 0 2620 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2083
timestamp 1713400504
transform 1 0 2588 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2084
timestamp 1713400504
transform 1 0 2492 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2085
timestamp 1713400504
transform 1 0 2388 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2086
timestamp 1713400504
transform 1 0 2620 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_2087
timestamp 1713400504
transform 1 0 2572 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2088
timestamp 1713400504
transform 1 0 2548 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2089
timestamp 1713400504
transform 1 0 2524 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_2090
timestamp 1713400504
transform 1 0 2596 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2091
timestamp 1713400504
transform 1 0 2556 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2092
timestamp 1713400504
transform 1 0 2564 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_2093
timestamp 1713400504
transform 1 0 2516 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2094
timestamp 1713400504
transform 1 0 2484 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2095
timestamp 1713400504
transform 1 0 2444 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_2096
timestamp 1713400504
transform 1 0 2420 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2097
timestamp 1713400504
transform 1 0 2492 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2098
timestamp 1713400504
transform 1 0 2428 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2099
timestamp 1713400504
transform 1 0 1860 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2100
timestamp 1713400504
transform 1 0 2732 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2101
timestamp 1713400504
transform 1 0 2532 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2102
timestamp 1713400504
transform 1 0 2524 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2103
timestamp 1713400504
transform 1 0 2540 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2104
timestamp 1713400504
transform 1 0 2540 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_2105
timestamp 1713400504
transform 1 0 2556 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_2106
timestamp 1713400504
transform 1 0 2540 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_2107
timestamp 1713400504
transform 1 0 2516 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_2108
timestamp 1713400504
transform 1 0 1996 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2109
timestamp 1713400504
transform 1 0 2556 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2110
timestamp 1713400504
transform 1 0 2500 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_2111
timestamp 1713400504
transform 1 0 1452 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2112
timestamp 1713400504
transform 1 0 2524 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2113
timestamp 1713400504
transform 1 0 2476 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2114
timestamp 1713400504
transform 1 0 1652 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2115
timestamp 1713400504
transform 1 0 2268 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2116
timestamp 1713400504
transform 1 0 1540 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2117
timestamp 1713400504
transform 1 0 2316 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2118
timestamp 1713400504
transform 1 0 1828 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2119
timestamp 1713400504
transform 1 0 2604 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2120
timestamp 1713400504
transform 1 0 2308 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_2121
timestamp 1713400504
transform 1 0 2652 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2122
timestamp 1713400504
transform 1 0 2636 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_2123
timestamp 1713400504
transform 1 0 2660 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2124
timestamp 1713400504
transform 1 0 2652 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2125
timestamp 1713400504
transform 1 0 2596 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2126
timestamp 1713400504
transform 1 0 2596 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2127
timestamp 1713400504
transform 1 0 2756 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2128
timestamp 1713400504
transform 1 0 2604 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2129
timestamp 1713400504
transform 1 0 2580 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_2130
timestamp 1713400504
transform 1 0 2580 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2131
timestamp 1713400504
transform 1 0 2556 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_2132
timestamp 1713400504
transform 1 0 2548 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2133
timestamp 1713400504
transform 1 0 2572 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2134
timestamp 1713400504
transform 1 0 2468 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2135
timestamp 1713400504
transform 1 0 1756 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2136
timestamp 1713400504
transform 1 0 1756 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2137
timestamp 1713400504
transform 1 0 1836 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2138
timestamp 1713400504
transform 1 0 1740 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2139
timestamp 1713400504
transform 1 0 2668 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2140
timestamp 1713400504
transform 1 0 2620 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2141
timestamp 1713400504
transform 1 0 2740 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2142
timestamp 1713400504
transform 1 0 2716 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2143
timestamp 1713400504
transform 1 0 2492 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_2144
timestamp 1713400504
transform 1 0 2396 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2145
timestamp 1713400504
transform 1 0 2508 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2146
timestamp 1713400504
transform 1 0 2508 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_2147
timestamp 1713400504
transform 1 0 1628 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2148
timestamp 1713400504
transform 1 0 1372 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2149
timestamp 1713400504
transform 1 0 1428 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2150
timestamp 1713400504
transform 1 0 1428 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_2151
timestamp 1713400504
transform 1 0 2764 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2152
timestamp 1713400504
transform 1 0 2740 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_2153
timestamp 1713400504
transform 1 0 2588 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2154
timestamp 1713400504
transform 1 0 2572 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2155
timestamp 1713400504
transform 1 0 2588 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2156
timestamp 1713400504
transform 1 0 2500 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2157
timestamp 1713400504
transform 1 0 2908 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2158
timestamp 1713400504
transform 1 0 2764 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_2159
timestamp 1713400504
transform 1 0 2852 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2160
timestamp 1713400504
transform 1 0 2828 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2161
timestamp 1713400504
transform 1 0 2852 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2162
timestamp 1713400504
transform 1 0 2820 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_2163
timestamp 1713400504
transform 1 0 2876 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2164
timestamp 1713400504
transform 1 0 2876 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2165
timestamp 1713400504
transform 1 0 2988 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2166
timestamp 1713400504
transform 1 0 2972 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_2167
timestamp 1713400504
transform 1 0 2844 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2168
timestamp 1713400504
transform 1 0 2652 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2169
timestamp 1713400504
transform 1 0 1996 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_2170
timestamp 1713400504
transform 1 0 1940 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2171
timestamp 1713400504
transform 1 0 2812 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2172
timestamp 1713400504
transform 1 0 2628 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2173
timestamp 1713400504
transform 1 0 2636 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2174
timestamp 1713400504
transform 1 0 2612 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_2175
timestamp 1713400504
transform 1 0 2644 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2176
timestamp 1713400504
transform 1 0 2644 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_2177
timestamp 1713400504
transform 1 0 2596 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_2178
timestamp 1713400504
transform 1 0 2596 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_2179
timestamp 1713400504
transform 1 0 2676 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2180
timestamp 1713400504
transform 1 0 2652 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2181
timestamp 1713400504
transform 1 0 2676 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_2182
timestamp 1713400504
transform 1 0 2548 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2183
timestamp 1713400504
transform 1 0 2660 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_2184
timestamp 1713400504
transform 1 0 2572 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_2185
timestamp 1713400504
transform 1 0 2580 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2186
timestamp 1713400504
transform 1 0 2492 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_2187
timestamp 1713400504
transform 1 0 2628 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2188
timestamp 1713400504
transform 1 0 2588 0 1 2835
box -2 -2 2 2
use M2_M1  M2_M1_2189
timestamp 1713400504
transform 1 0 2644 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2190
timestamp 1713400504
transform 1 0 2540 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2191
timestamp 1713400504
transform 1 0 2604 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_2192
timestamp 1713400504
transform 1 0 2588 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2193
timestamp 1713400504
transform 1 0 2644 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2194
timestamp 1713400504
transform 1 0 2628 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2195
timestamp 1713400504
transform 1 0 2700 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2196
timestamp 1713400504
transform 1 0 2620 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2197
timestamp 1713400504
transform 1 0 2892 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2198
timestamp 1713400504
transform 1 0 2804 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_2199
timestamp 1713400504
transform 1 0 2852 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2200
timestamp 1713400504
transform 1 0 2852 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2201
timestamp 1713400504
transform 1 0 2892 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2202
timestamp 1713400504
transform 1 0 2876 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2203
timestamp 1713400504
transform 1 0 2924 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2204
timestamp 1713400504
transform 1 0 2924 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2205
timestamp 1713400504
transform 1 0 1764 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_2206
timestamp 1713400504
transform 1 0 1396 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_2207
timestamp 1713400504
transform 1 0 1804 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2208
timestamp 1713400504
transform 1 0 1788 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2209
timestamp 1713400504
transform 1 0 1764 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2210
timestamp 1713400504
transform 1 0 1724 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_2211
timestamp 1713400504
transform 1 0 1852 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2212
timestamp 1713400504
transform 1 0 1740 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2213
timestamp 1713400504
transform 1 0 1732 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_2214
timestamp 1713400504
transform 1 0 1732 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2215
timestamp 1713400504
transform 1 0 1700 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2216
timestamp 1713400504
transform 1 0 1676 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2217
timestamp 1713400504
transform 1 0 1700 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_2218
timestamp 1713400504
transform 1 0 1652 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2219
timestamp 1713400504
transform 1 0 1588 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2220
timestamp 1713400504
transform 1 0 1572 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2221
timestamp 1713400504
transform 1 0 1628 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2222
timestamp 1713400504
transform 1 0 1596 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2223
timestamp 1713400504
transform 1 0 1828 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2224
timestamp 1713400504
transform 1 0 1828 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2225
timestamp 1713400504
transform 1 0 1692 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2226
timestamp 1713400504
transform 1 0 1364 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_2227
timestamp 1713400504
transform 1 0 1372 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2228
timestamp 1713400504
transform 1 0 1108 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2229
timestamp 1713400504
transform 1 0 1308 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2230
timestamp 1713400504
transform 1 0 1308 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_2231
timestamp 1713400504
transform 1 0 1324 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2232
timestamp 1713400504
transform 1 0 1236 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2233
timestamp 1713400504
transform 1 0 1268 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_2234
timestamp 1713400504
transform 1 0 1252 0 1 2705
box -2 -2 2 2
use M2_M1  M2_M1_2235
timestamp 1713400504
transform 1 0 1292 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2236
timestamp 1713400504
transform 1 0 1268 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2237
timestamp 1713400504
transform 1 0 1292 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_2238
timestamp 1713400504
transform 1 0 1260 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_2239
timestamp 1713400504
transform 1 0 1852 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2240
timestamp 1713400504
transform 1 0 1676 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2241
timestamp 1713400504
transform 1 0 1548 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2242
timestamp 1713400504
transform 1 0 1484 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_2243
timestamp 1713400504
transform 1 0 1556 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2244
timestamp 1713400504
transform 1 0 1556 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2245
timestamp 1713400504
transform 1 0 1484 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2246
timestamp 1713400504
transform 1 0 1452 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2247
timestamp 1713400504
transform 1 0 1476 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_2248
timestamp 1713400504
transform 1 0 1468 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2249
timestamp 1713400504
transform 1 0 2556 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2250
timestamp 1713400504
transform 1 0 1548 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_2251
timestamp 1713400504
transform 1 0 2516 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2252
timestamp 1713400504
transform 1 0 2500 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2253
timestamp 1713400504
transform 1 0 2548 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_2254
timestamp 1713400504
transform 1 0 2548 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2255
timestamp 1713400504
transform 1 0 2540 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2256
timestamp 1713400504
transform 1 0 2524 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2257
timestamp 1713400504
transform 1 0 2684 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2258
timestamp 1713400504
transform 1 0 2572 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2259
timestamp 1713400504
transform 1 0 1508 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2260
timestamp 1713400504
transform 1 0 1452 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2261
timestamp 1713400504
transform 1 0 1636 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2262
timestamp 1713400504
transform 1 0 1524 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2263
timestamp 1713400504
transform 1 0 1532 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2264
timestamp 1713400504
transform 1 0 1524 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2265
timestamp 1713400504
transform 1 0 1412 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2266
timestamp 1713400504
transform 1 0 1412 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2267
timestamp 1713400504
transform 1 0 1476 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_2268
timestamp 1713400504
transform 1 0 1444 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2269
timestamp 1713400504
transform 1 0 1396 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2270
timestamp 1713400504
transform 1 0 1348 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2271
timestamp 1713400504
transform 1 0 1836 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2272
timestamp 1713400504
transform 1 0 1508 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2273
timestamp 1713400504
transform 1 0 2444 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2274
timestamp 1713400504
transform 1 0 2444 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2275
timestamp 1713400504
transform 1 0 2084 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2276
timestamp 1713400504
transform 1 0 2084 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2277
timestamp 1713400504
transform 1 0 2180 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2278
timestamp 1713400504
transform 1 0 2172 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2279
timestamp 1713400504
transform 1 0 2124 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2280
timestamp 1713400504
transform 1 0 2100 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2281
timestamp 1713400504
transform 1 0 2100 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_2282
timestamp 1713400504
transform 1 0 2084 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_2283
timestamp 1713400504
transform 1 0 2172 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2284
timestamp 1713400504
transform 1 0 2164 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2285
timestamp 1713400504
transform 1 0 2172 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2286
timestamp 1713400504
transform 1 0 2172 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2287
timestamp 1713400504
transform 1 0 2100 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2288
timestamp 1713400504
transform 1 0 2084 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2289
timestamp 1713400504
transform 1 0 2748 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2290
timestamp 1713400504
transform 1 0 2428 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2291
timestamp 1713400504
transform 1 0 2764 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2292
timestamp 1713400504
transform 1 0 2420 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2293
timestamp 1713400504
transform 1 0 2540 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2294
timestamp 1713400504
transform 1 0 2396 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2295
timestamp 1713400504
transform 1 0 2380 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2296
timestamp 1713400504
transform 1 0 2356 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2297
timestamp 1713400504
transform 1 0 2452 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2298
timestamp 1713400504
transform 1 0 2436 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2299
timestamp 1713400504
transform 1 0 2716 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2300
timestamp 1713400504
transform 1 0 2428 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2301
timestamp 1713400504
transform 1 0 2684 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_2302
timestamp 1713400504
transform 1 0 2412 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2303
timestamp 1713400504
transform 1 0 2724 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_2304
timestamp 1713400504
transform 1 0 2420 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2305
timestamp 1713400504
transform 1 0 2332 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_2306
timestamp 1713400504
transform 1 0 2300 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2307
timestamp 1713400504
transform 1 0 2380 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_2308
timestamp 1713400504
transform 1 0 2372 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2309
timestamp 1713400504
transform 1 0 2356 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_2310
timestamp 1713400504
transform 1 0 2348 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2311
timestamp 1713400504
transform 1 0 2260 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_2312
timestamp 1713400504
transform 1 0 2244 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2313
timestamp 1713400504
transform 1 0 2132 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_2314
timestamp 1713400504
transform 1 0 2132 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2315
timestamp 1713400504
transform 1 0 2084 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_2316
timestamp 1713400504
transform 1 0 2084 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2317
timestamp 1713400504
transform 1 0 1852 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2318
timestamp 1713400504
transform 1 0 1668 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_2319
timestamp 1713400504
transform 1 0 1860 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2320
timestamp 1713400504
transform 1 0 1572 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_2321
timestamp 1713400504
transform 1 0 1900 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2322
timestamp 1713400504
transform 1 0 1620 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_2323
timestamp 1713400504
transform 1 0 1812 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2324
timestamp 1713400504
transform 1 0 1604 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_2325
timestamp 1713400504
transform 1 0 1868 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2326
timestamp 1713400504
transform 1 0 1660 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_2327
timestamp 1713400504
transform 1 0 1868 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2328
timestamp 1713400504
transform 1 0 1868 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2329
timestamp 1713400504
transform 1 0 2076 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2330
timestamp 1713400504
transform 1 0 2068 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2331
timestamp 1713400504
transform 1 0 2092 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2332
timestamp 1713400504
transform 1 0 2092 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2333
timestamp 1713400504
transform 1 0 2132 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2334
timestamp 1713400504
transform 1 0 2076 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2335
timestamp 1713400504
transform 1 0 2076 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2336
timestamp 1713400504
transform 1 0 1788 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2337
timestamp 1713400504
transform 1 0 1788 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2338
timestamp 1713400504
transform 1 0 1764 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2339
timestamp 1713400504
transform 1 0 1756 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2340
timestamp 1713400504
transform 1 0 1740 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2341
timestamp 1713400504
transform 1 0 1716 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2342
timestamp 1713400504
transform 1 0 1716 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2343
timestamp 1713400504
transform 1 0 1700 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2344
timestamp 1713400504
transform 1 0 1796 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2345
timestamp 1713400504
transform 1 0 1796 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2346
timestamp 1713400504
transform 1 0 1772 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2347
timestamp 1713400504
transform 1 0 1772 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2348
timestamp 1713400504
transform 1 0 1732 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2349
timestamp 1713400504
transform 1 0 1732 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2350
timestamp 1713400504
transform 1 0 1836 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2351
timestamp 1713400504
transform 1 0 1828 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2352
timestamp 1713400504
transform 1 0 1892 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2353
timestamp 1713400504
transform 1 0 1852 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2354
timestamp 1713400504
transform 1 0 1940 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2355
timestamp 1713400504
transform 1 0 1852 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2356
timestamp 1713400504
transform 1 0 2316 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2357
timestamp 1713400504
transform 1 0 2212 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2358
timestamp 1713400504
transform 1 0 2148 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2359
timestamp 1713400504
transform 1 0 2148 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2360
timestamp 1713400504
transform 1 0 2108 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2361
timestamp 1713400504
transform 1 0 2028 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2362
timestamp 1713400504
transform 1 0 1988 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2363
timestamp 1713400504
transform 1 0 2052 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2364
timestamp 1713400504
transform 1 0 2052 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2365
timestamp 1713400504
transform 1 0 1948 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2366
timestamp 1713400504
transform 1 0 1868 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2367
timestamp 1713400504
transform 1 0 1404 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2368
timestamp 1713400504
transform 1 0 2164 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2369
timestamp 1713400504
transform 1 0 2060 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2370
timestamp 1713400504
transform 1 0 2044 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_2371
timestamp 1713400504
transform 1 0 2044 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2372
timestamp 1713400504
transform 1 0 1388 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2373
timestamp 1713400504
transform 1 0 2132 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2374
timestamp 1713400504
transform 1 0 2044 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2375
timestamp 1713400504
transform 1 0 2020 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2376
timestamp 1713400504
transform 1 0 1948 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2377
timestamp 1713400504
transform 1 0 1524 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2378
timestamp 1713400504
transform 1 0 2316 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2379
timestamp 1713400504
transform 1 0 2292 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2380
timestamp 1713400504
transform 1 0 2060 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2381
timestamp 1713400504
transform 1 0 2004 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2382
timestamp 1713400504
transform 1 0 1964 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2383
timestamp 1713400504
transform 1 0 1940 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2384
timestamp 1713400504
transform 1 0 1612 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2385
timestamp 1713400504
transform 1 0 2140 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2386
timestamp 1713400504
transform 1 0 2124 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2387
timestamp 1713400504
transform 1 0 2028 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2388
timestamp 1713400504
transform 1 0 2204 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2389
timestamp 1713400504
transform 1 0 2196 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2390
timestamp 1713400504
transform 1 0 2300 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2391
timestamp 1713400504
transform 1 0 2292 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2392
timestamp 1713400504
transform 1 0 2268 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2393
timestamp 1713400504
transform 1 0 2324 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2394
timestamp 1713400504
transform 1 0 2220 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2395
timestamp 1713400504
transform 1 0 2340 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2396
timestamp 1713400504
transform 1 0 2164 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2397
timestamp 1713400504
transform 1 0 2196 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2398
timestamp 1713400504
transform 1 0 2148 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2399
timestamp 1713400504
transform 1 0 2148 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2400
timestamp 1713400504
transform 1 0 2100 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2401
timestamp 1713400504
transform 1 0 1980 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2402
timestamp 1713400504
transform 1 0 1916 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2403
timestamp 1713400504
transform 1 0 2244 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2404
timestamp 1713400504
transform 1 0 2188 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2405
timestamp 1713400504
transform 1 0 2076 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2406
timestamp 1713400504
transform 1 0 2076 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2407
timestamp 1713400504
transform 1 0 1940 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2408
timestamp 1713400504
transform 1 0 1916 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2409
timestamp 1713400504
transform 1 0 1836 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2410
timestamp 1713400504
transform 1 0 1636 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2411
timestamp 1713400504
transform 1 0 1636 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2412
timestamp 1713400504
transform 1 0 1572 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2413
timestamp 1713400504
transform 1 0 1564 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2414
timestamp 1713400504
transform 1 0 1564 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2415
timestamp 1713400504
transform 1 0 1620 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2416
timestamp 1713400504
transform 1 0 1620 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2417
timestamp 1713400504
transform 1 0 1716 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2418
timestamp 1713400504
transform 1 0 1604 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2419
timestamp 1713400504
transform 1 0 1684 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2420
timestamp 1713400504
transform 1 0 1684 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2421
timestamp 1713400504
transform 1 0 1628 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2422
timestamp 1713400504
transform 1 0 1588 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2423
timestamp 1713400504
transform 1 0 1588 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_2424
timestamp 1713400504
transform 1 0 1804 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2425
timestamp 1713400504
transform 1 0 1740 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2426
timestamp 1713400504
transform 1 0 1740 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2427
timestamp 1713400504
transform 1 0 1708 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2428
timestamp 1713400504
transform 1 0 1820 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2429
timestamp 1713400504
transform 1 0 1796 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2430
timestamp 1713400504
transform 1 0 1796 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_2431
timestamp 1713400504
transform 1 0 1756 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2432
timestamp 1713400504
transform 1 0 1740 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2433
timestamp 1713400504
transform 1 0 1724 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2434
timestamp 1713400504
transform 1 0 1852 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2435
timestamp 1713400504
transform 1 0 1852 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2436
timestamp 1713400504
transform 1 0 1724 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2437
timestamp 1713400504
transform 1 0 1908 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2438
timestamp 1713400504
transform 1 0 1724 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2439
timestamp 1713400504
transform 1 0 1716 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2440
timestamp 1713400504
transform 1 0 1716 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2441
timestamp 1713400504
transform 1 0 1556 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2442
timestamp 1713400504
transform 1 0 1732 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2443
timestamp 1713400504
transform 1 0 1500 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2444
timestamp 1713400504
transform 1 0 1948 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2445
timestamp 1713400504
transform 1 0 1940 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2446
timestamp 1713400504
transform 1 0 1868 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2447
timestamp 1713400504
transform 1 0 1852 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2448
timestamp 1713400504
transform 1 0 1812 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2449
timestamp 1713400504
transform 1 0 1724 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2450
timestamp 1713400504
transform 1 0 1604 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2451
timestamp 1713400504
transform 1 0 1596 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_2452
timestamp 1713400504
transform 1 0 1596 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2453
timestamp 1713400504
transform 1 0 1684 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_2454
timestamp 1713400504
transform 1 0 1604 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2455
timestamp 1713400504
transform 1 0 1804 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2456
timestamp 1713400504
transform 1 0 1772 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2457
timestamp 1713400504
transform 1 0 1812 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2458
timestamp 1713400504
transform 1 0 1716 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2459
timestamp 1713400504
transform 1 0 1852 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2460
timestamp 1713400504
transform 1 0 1852 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2461
timestamp 1713400504
transform 1 0 1804 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2462
timestamp 1713400504
transform 1 0 1668 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2463
timestamp 1713400504
transform 1 0 1668 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2464
timestamp 1713400504
transform 1 0 1620 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2465
timestamp 1713400504
transform 1 0 1508 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2466
timestamp 1713400504
transform 1 0 1508 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2467
timestamp 1713400504
transform 1 0 1508 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2468
timestamp 1713400504
transform 1 0 1700 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2469
timestamp 1713400504
transform 1 0 1612 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2470
timestamp 1713400504
transform 1 0 1612 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2471
timestamp 1713400504
transform 1 0 1732 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2472
timestamp 1713400504
transform 1 0 1708 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2473
timestamp 1713400504
transform 1 0 1812 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2474
timestamp 1713400504
transform 1 0 1788 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2475
timestamp 1713400504
transform 1 0 1692 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2476
timestamp 1713400504
transform 1 0 1588 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2477
timestamp 1713400504
transform 1 0 1708 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2478
timestamp 1713400504
transform 1 0 1708 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2479
timestamp 1713400504
transform 1 0 1716 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2480
timestamp 1713400504
transform 1 0 1468 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2481
timestamp 1713400504
transform 1 0 1708 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2482
timestamp 1713400504
transform 1 0 1708 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2483
timestamp 1713400504
transform 1 0 1692 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2484
timestamp 1713400504
transform 1 0 1716 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2485
timestamp 1713400504
transform 1 0 1620 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2486
timestamp 1713400504
transform 1 0 1580 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2487
timestamp 1713400504
transform 1 0 1564 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2488
timestamp 1713400504
transform 1 0 1924 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2489
timestamp 1713400504
transform 1 0 1892 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2490
timestamp 1713400504
transform 1 0 1836 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2491
timestamp 1713400504
transform 1 0 1828 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2492
timestamp 1713400504
transform 1 0 1780 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2493
timestamp 1713400504
transform 1 0 1772 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_2494
timestamp 1713400504
transform 1 0 1708 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2495
timestamp 1713400504
transform 1 0 1580 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2496
timestamp 1713400504
transform 1 0 1700 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2497
timestamp 1713400504
transform 1 0 1684 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2498
timestamp 1713400504
transform 1 0 1628 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2499
timestamp 1713400504
transform 1 0 1620 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2500
timestamp 1713400504
transform 1 0 1620 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2501
timestamp 1713400504
transform 1 0 1524 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2502
timestamp 1713400504
transform 1 0 1524 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2503
timestamp 1713400504
transform 1 0 1708 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2504
timestamp 1713400504
transform 1 0 1692 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2505
timestamp 1713400504
transform 1 0 1532 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2506
timestamp 1713400504
transform 1 0 1468 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2507
timestamp 1713400504
transform 1 0 1468 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2508
timestamp 1713400504
transform 1 0 1636 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2509
timestamp 1713400504
transform 1 0 1572 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2510
timestamp 1713400504
transform 1 0 1572 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2511
timestamp 1713400504
transform 1 0 1436 0 1 1055
box -2 -2 2 2
use M2_M1  M2_M1_2512
timestamp 1713400504
transform 1 0 1436 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2513
timestamp 1713400504
transform 1 0 1396 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2514
timestamp 1713400504
transform 1 0 1396 0 1 1055
box -2 -2 2 2
use M2_M1  M2_M1_2515
timestamp 1713400504
transform 1 0 1588 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2516
timestamp 1713400504
transform 1 0 1588 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2517
timestamp 1713400504
transform 1 0 1580 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2518
timestamp 1713400504
transform 1 0 1404 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2519
timestamp 1713400504
transform 1 0 1308 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2520
timestamp 1713400504
transform 1 0 1508 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2521
timestamp 1713400504
transform 1 0 1492 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2522
timestamp 1713400504
transform 1 0 1508 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2523
timestamp 1713400504
transform 1 0 1420 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2524
timestamp 1713400504
transform 1 0 1484 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2525
timestamp 1713400504
transform 1 0 1420 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2526
timestamp 1713400504
transform 1 0 1436 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2527
timestamp 1713400504
transform 1 0 1324 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2528
timestamp 1713400504
transform 1 0 1612 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2529
timestamp 1713400504
transform 1 0 1596 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2530
timestamp 1713400504
transform 1 0 1676 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2531
timestamp 1713400504
transform 1 0 1620 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2532
timestamp 1713400504
transform 1 0 1692 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2533
timestamp 1713400504
transform 1 0 1588 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2534
timestamp 1713400504
transform 1 0 1588 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2535
timestamp 1713400504
transform 1 0 1476 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2536
timestamp 1713400504
transform 1 0 1532 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2537
timestamp 1713400504
transform 1 0 1484 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2538
timestamp 1713400504
transform 1 0 1588 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2539
timestamp 1713400504
transform 1 0 1468 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2540
timestamp 1713400504
transform 1 0 1300 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2541
timestamp 1713400504
transform 1 0 1292 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2542
timestamp 1713400504
transform 1 0 1356 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2543
timestamp 1713400504
transform 1 0 1324 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2544
timestamp 1713400504
transform 1 0 1244 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2545
timestamp 1713400504
transform 1 0 1244 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2546
timestamp 1713400504
transform 1 0 1148 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2547
timestamp 1713400504
transform 1 0 892 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2548
timestamp 1713400504
transform 1 0 1100 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2549
timestamp 1713400504
transform 1 0 1100 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2550
timestamp 1713400504
transform 1 0 1004 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2551
timestamp 1713400504
transform 1 0 860 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2552
timestamp 1713400504
transform 1 0 1084 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2553
timestamp 1713400504
transform 1 0 1076 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2554
timestamp 1713400504
transform 1 0 1044 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2555
timestamp 1713400504
transform 1 0 1044 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2556
timestamp 1713400504
transform 1 0 1036 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2557
timestamp 1713400504
transform 1 0 964 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2558
timestamp 1713400504
transform 1 0 964 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2559
timestamp 1713400504
transform 1 0 964 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2560
timestamp 1713400504
transform 1 0 916 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2561
timestamp 1713400504
transform 1 0 916 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2562
timestamp 1713400504
transform 1 0 916 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2563
timestamp 1713400504
transform 1 0 1148 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2564
timestamp 1713400504
transform 1 0 1116 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2565
timestamp 1713400504
transform 1 0 1084 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2566
timestamp 1713400504
transform 1 0 1020 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2567
timestamp 1713400504
transform 1 0 980 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2568
timestamp 1713400504
transform 1 0 980 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2569
timestamp 1713400504
transform 1 0 980 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2570
timestamp 1713400504
transform 1 0 980 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2571
timestamp 1713400504
transform 1 0 964 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2572
timestamp 1713400504
transform 1 0 1004 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2573
timestamp 1713400504
transform 1 0 964 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2574
timestamp 1713400504
transform 1 0 924 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2575
timestamp 1713400504
transform 1 0 876 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2576
timestamp 1713400504
transform 1 0 860 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2577
timestamp 1713400504
transform 1 0 772 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2578
timestamp 1713400504
transform 1 0 724 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2579
timestamp 1713400504
transform 1 0 724 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2580
timestamp 1713400504
transform 1 0 1036 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2581
timestamp 1713400504
transform 1 0 972 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2582
timestamp 1713400504
transform 1 0 884 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2583
timestamp 1713400504
transform 1 0 876 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2584
timestamp 1713400504
transform 1 0 868 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2585
timestamp 1713400504
transform 1 0 756 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2586
timestamp 1713400504
transform 1 0 748 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2587
timestamp 1713400504
transform 1 0 868 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2588
timestamp 1713400504
transform 1 0 748 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2589
timestamp 1713400504
transform 1 0 972 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2590
timestamp 1713400504
transform 1 0 876 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2591
timestamp 1713400504
transform 1 0 1156 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2592
timestamp 1713400504
transform 1 0 1156 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2593
timestamp 1713400504
transform 1 0 996 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2594
timestamp 1713400504
transform 1 0 964 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2595
timestamp 1713400504
transform 1 0 1012 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2596
timestamp 1713400504
transform 1 0 1012 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2597
timestamp 1713400504
transform 1 0 1124 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2598
timestamp 1713400504
transform 1 0 1028 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2599
timestamp 1713400504
transform 1 0 1108 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2600
timestamp 1713400504
transform 1 0 1108 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2601
timestamp 1713400504
transform 1 0 1268 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2602
timestamp 1713400504
transform 1 0 868 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2603
timestamp 1713400504
transform 1 0 860 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2604
timestamp 1713400504
transform 1 0 852 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2605
timestamp 1713400504
transform 1 0 892 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2606
timestamp 1713400504
transform 1 0 884 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2607
timestamp 1713400504
transform 1 0 868 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2608
timestamp 1713400504
transform 1 0 860 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2609
timestamp 1713400504
transform 1 0 972 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2610
timestamp 1713400504
transform 1 0 868 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2611
timestamp 1713400504
transform 1 0 764 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2612
timestamp 1713400504
transform 1 0 740 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2613
timestamp 1713400504
transform 1 0 956 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2614
timestamp 1713400504
transform 1 0 844 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2615
timestamp 1713400504
transform 1 0 1540 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_2616
timestamp 1713400504
transform 1 0 1540 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2617
timestamp 1713400504
transform 1 0 1620 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2618
timestamp 1713400504
transform 1 0 1564 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2619
timestamp 1713400504
transform 1 0 1492 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2620
timestamp 1713400504
transform 1 0 1492 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2621
timestamp 1713400504
transform 1 0 1468 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2622
timestamp 1713400504
transform 1 0 1420 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2623
timestamp 1713400504
transform 1 0 1308 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2624
timestamp 1713400504
transform 1 0 1300 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2625
timestamp 1713400504
transform 1 0 1316 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2626
timestamp 1713400504
transform 1 0 1268 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2627
timestamp 1713400504
transform 1 0 1300 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2628
timestamp 1713400504
transform 1 0 1276 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2629
timestamp 1713400504
transform 1 0 1236 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2630
timestamp 1713400504
transform 1 0 1236 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2631
timestamp 1713400504
transform 1 0 1236 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2632
timestamp 1713400504
transform 1 0 1172 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2633
timestamp 1713400504
transform 1 0 1172 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2634
timestamp 1713400504
transform 1 0 1172 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2635
timestamp 1713400504
transform 1 0 1164 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2636
timestamp 1713400504
transform 1 0 1164 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2637
timestamp 1713400504
transform 1 0 1308 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2638
timestamp 1713400504
transform 1 0 1292 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2639
timestamp 1713400504
transform 1 0 1252 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2640
timestamp 1713400504
transform 1 0 1212 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2641
timestamp 1713400504
transform 1 0 1188 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2642
timestamp 1713400504
transform 1 0 1188 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2643
timestamp 1713400504
transform 1 0 1116 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2644
timestamp 1713400504
transform 1 0 1356 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2645
timestamp 1713400504
transform 1 0 1284 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2646
timestamp 1713400504
transform 1 0 1284 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2647
timestamp 1713400504
transform 1 0 1284 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2648
timestamp 1713400504
transform 1 0 1164 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2649
timestamp 1713400504
transform 1 0 1164 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2650
timestamp 1713400504
transform 1 0 1164 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2651
timestamp 1713400504
transform 1 0 1412 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2652
timestamp 1713400504
transform 1 0 1380 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2653
timestamp 1713400504
transform 1 0 1324 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2654
timestamp 1713400504
transform 1 0 1300 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2655
timestamp 1713400504
transform 1 0 1268 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2656
timestamp 1713400504
transform 1 0 1212 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2657
timestamp 1713400504
transform 1 0 1188 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2658
timestamp 1713400504
transform 1 0 1252 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2659
timestamp 1713400504
transform 1 0 1204 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2660
timestamp 1713400504
transform 1 0 1188 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2661
timestamp 1713400504
transform 1 0 1180 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2662
timestamp 1713400504
transform 1 0 1428 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2663
timestamp 1713400504
transform 1 0 1428 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2664
timestamp 1713400504
transform 1 0 1332 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2665
timestamp 1713400504
transform 1 0 1260 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2666
timestamp 1713400504
transform 1 0 1268 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2667
timestamp 1713400504
transform 1 0 1244 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2668
timestamp 1713400504
transform 1 0 1380 0 1 755
box -2 -2 2 2
use M2_M1  M2_M1_2669
timestamp 1713400504
transform 1 0 1380 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2670
timestamp 1713400504
transform 1 0 1292 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2671
timestamp 1713400504
transform 1 0 1292 0 1 755
box -2 -2 2 2
use M2_M1  M2_M1_2672
timestamp 1713400504
transform 1 0 1324 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2673
timestamp 1713400504
transform 1 0 1204 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2674
timestamp 1713400504
transform 1 0 1524 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2675
timestamp 1713400504
transform 1 0 1524 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2676
timestamp 1713400504
transform 1 0 1540 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2677
timestamp 1713400504
transform 1 0 1436 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2678
timestamp 1713400504
transform 1 0 1372 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2679
timestamp 1713400504
transform 1 0 1356 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2680
timestamp 1713400504
transform 1 0 1308 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2681
timestamp 1713400504
transform 1 0 1284 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2682
timestamp 1713400504
transform 1 0 1444 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2683
timestamp 1713400504
transform 1 0 1404 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2684
timestamp 1713400504
transform 1 0 1388 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2685
timestamp 1713400504
transform 1 0 1180 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2686
timestamp 1713400504
transform 1 0 1460 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2687
timestamp 1713400504
transform 1 0 1276 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2688
timestamp 1713400504
transform 1 0 1484 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2689
timestamp 1713400504
transform 1 0 1460 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2690
timestamp 1713400504
transform 1 0 1292 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2691
timestamp 1713400504
transform 1 0 1292 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2692
timestamp 1713400504
transform 1 0 1300 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2693
timestamp 1713400504
transform 1 0 1236 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2694
timestamp 1713400504
transform 1 0 1156 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2695
timestamp 1713400504
transform 1 0 932 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2696
timestamp 1713400504
transform 1 0 1084 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_2697
timestamp 1713400504
transform 1 0 1036 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2698
timestamp 1713400504
transform 1 0 860 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2699
timestamp 1713400504
transform 1 0 724 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2700
timestamp 1713400504
transform 1 0 1060 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2701
timestamp 1713400504
transform 1 0 948 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2702
timestamp 1713400504
transform 1 0 1076 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2703
timestamp 1713400504
transform 1 0 1076 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2704
timestamp 1713400504
transform 1 0 1076 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2705
timestamp 1713400504
transform 1 0 1020 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2706
timestamp 1713400504
transform 1 0 1020 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2707
timestamp 1713400504
transform 1 0 836 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2708
timestamp 1713400504
transform 1 0 836 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2709
timestamp 1713400504
transform 1 0 828 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2710
timestamp 1713400504
transform 1 0 1148 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2711
timestamp 1713400504
transform 1 0 1148 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2712
timestamp 1713400504
transform 1 0 1092 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2713
timestamp 1713400504
transform 1 0 1068 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2714
timestamp 1713400504
transform 1 0 852 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2715
timestamp 1713400504
transform 1 0 852 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2716
timestamp 1713400504
transform 1 0 844 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2717
timestamp 1713400504
transform 1 0 988 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2718
timestamp 1713400504
transform 1 0 948 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2719
timestamp 1713400504
transform 1 0 948 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2720
timestamp 1713400504
transform 1 0 724 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2721
timestamp 1713400504
transform 1 0 716 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2722
timestamp 1713400504
transform 1 0 628 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2723
timestamp 1713400504
transform 1 0 628 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2724
timestamp 1713400504
transform 1 0 572 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2725
timestamp 1713400504
transform 1 0 540 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2726
timestamp 1713400504
transform 1 0 972 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2727
timestamp 1713400504
transform 1 0 972 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2728
timestamp 1713400504
transform 1 0 964 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2729
timestamp 1713400504
transform 1 0 740 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2730
timestamp 1713400504
transform 1 0 732 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2731
timestamp 1713400504
transform 1 0 660 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2732
timestamp 1713400504
transform 1 0 556 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2733
timestamp 1713400504
transform 1 0 820 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2734
timestamp 1713400504
transform 1 0 732 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2735
timestamp 1713400504
transform 1 0 836 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2736
timestamp 1713400504
transform 1 0 836 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2737
timestamp 1713400504
transform 1 0 1212 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2738
timestamp 1713400504
transform 1 0 1212 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2739
timestamp 1713400504
transform 1 0 1164 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2740
timestamp 1713400504
transform 1 0 1092 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2741
timestamp 1713400504
transform 1 0 980 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2742
timestamp 1713400504
transform 1 0 956 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2743
timestamp 1713400504
transform 1 0 1140 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2744
timestamp 1713400504
transform 1 0 1028 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2745
timestamp 1713400504
transform 1 0 1124 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2746
timestamp 1713400504
transform 1 0 964 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2747
timestamp 1713400504
transform 1 0 1132 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2748
timestamp 1713400504
transform 1 0 1084 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2749
timestamp 1713400504
transform 1 0 1244 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2750
timestamp 1713400504
transform 1 0 828 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2751
timestamp 1713400504
transform 1 0 756 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2752
timestamp 1713400504
transform 1 0 756 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2753
timestamp 1713400504
transform 1 0 676 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2754
timestamp 1713400504
transform 1 0 548 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2755
timestamp 1713400504
transform 1 0 844 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2756
timestamp 1713400504
transform 1 0 740 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2757
timestamp 1713400504
transform 1 0 652 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2758
timestamp 1713400504
transform 1 0 644 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2759
timestamp 1713400504
transform 1 0 844 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2760
timestamp 1713400504
transform 1 0 652 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2761
timestamp 1713400504
transform 1 0 1380 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2762
timestamp 1713400504
transform 1 0 1228 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2763
timestamp 1713400504
transform 1 0 1404 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2764
timestamp 1713400504
transform 1 0 1372 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2765
timestamp 1713400504
transform 1 0 1268 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2766
timestamp 1713400504
transform 1 0 1148 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2767
timestamp 1713400504
transform 1 0 1252 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2768
timestamp 1713400504
transform 1 0 1092 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2769
timestamp 1713400504
transform 1 0 972 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2770
timestamp 1713400504
transform 1 0 972 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2771
timestamp 1713400504
transform 1 0 1100 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2772
timestamp 1713400504
transform 1 0 1044 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2773
timestamp 1713400504
transform 1 0 1044 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2774
timestamp 1713400504
transform 1 0 764 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2775
timestamp 1713400504
transform 1 0 988 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2776
timestamp 1713400504
transform 1 0 980 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2777
timestamp 1713400504
transform 1 0 1100 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2778
timestamp 1713400504
transform 1 0 1020 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2779
timestamp 1713400504
transform 1 0 940 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2780
timestamp 1713400504
transform 1 0 900 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2781
timestamp 1713400504
transform 1 0 852 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2782
timestamp 1713400504
transform 1 0 844 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2783
timestamp 1713400504
transform 1 0 844 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2784
timestamp 1713400504
transform 1 0 820 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2785
timestamp 1713400504
transform 1 0 820 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2786
timestamp 1713400504
transform 1 0 1108 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2787
timestamp 1713400504
transform 1 0 996 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2788
timestamp 1713400504
transform 1 0 996 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2789
timestamp 1713400504
transform 1 0 956 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2790
timestamp 1713400504
transform 1 0 884 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2791
timestamp 1713400504
transform 1 0 884 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2792
timestamp 1713400504
transform 1 0 836 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2793
timestamp 1713400504
transform 1 0 1148 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2794
timestamp 1713400504
transform 1 0 1140 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2795
timestamp 1713400504
transform 1 0 972 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2796
timestamp 1713400504
transform 1 0 796 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2797
timestamp 1713400504
transform 1 0 764 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2798
timestamp 1713400504
transform 1 0 764 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2799
timestamp 1713400504
transform 1 0 756 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2800
timestamp 1713400504
transform 1 0 1164 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2801
timestamp 1713400504
transform 1 0 1100 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2802
timestamp 1713400504
transform 1 0 1012 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2803
timestamp 1713400504
transform 1 0 876 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2804
timestamp 1713400504
transform 1 0 812 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2805
timestamp 1713400504
transform 1 0 780 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2806
timestamp 1713400504
transform 1 0 772 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2807
timestamp 1713400504
transform 1 0 900 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2808
timestamp 1713400504
transform 1 0 772 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2809
timestamp 1713400504
transform 1 0 892 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2810
timestamp 1713400504
transform 1 0 876 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2811
timestamp 1713400504
transform 1 0 1100 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2812
timestamp 1713400504
transform 1 0 1092 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2813
timestamp 1713400504
transform 1 0 1180 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2814
timestamp 1713400504
transform 1 0 1132 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2815
timestamp 1713400504
transform 1 0 1156 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2816
timestamp 1713400504
transform 1 0 1140 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2817
timestamp 1713400504
transform 1 0 1108 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2818
timestamp 1713400504
transform 1 0 1100 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2819
timestamp 1713400504
transform 1 0 1004 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2820
timestamp 1713400504
transform 1 0 1004 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2821
timestamp 1713400504
transform 1 0 972 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2822
timestamp 1713400504
transform 1 0 948 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2823
timestamp 1713400504
transform 1 0 1172 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2824
timestamp 1713400504
transform 1 0 964 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2825
timestamp 1713400504
transform 1 0 924 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2826
timestamp 1713400504
transform 1 0 924 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2827
timestamp 1713400504
transform 1 0 980 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2828
timestamp 1713400504
transform 1 0 972 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2829
timestamp 1713400504
transform 1 0 892 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2830
timestamp 1713400504
transform 1 0 868 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2831
timestamp 1713400504
transform 1 0 900 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2832
timestamp 1713400504
transform 1 0 876 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2833
timestamp 1713400504
transform 1 0 828 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2834
timestamp 1713400504
transform 1 0 804 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2835
timestamp 1713400504
transform 1 0 836 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2836
timestamp 1713400504
transform 1 0 828 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2837
timestamp 1713400504
transform 1 0 2556 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2838
timestamp 1713400504
transform 1 0 2508 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2839
timestamp 1713400504
transform 1 0 2380 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2840
timestamp 1713400504
transform 1 0 2380 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2841
timestamp 1713400504
transform 1 0 2564 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2842
timestamp 1713400504
transform 1 0 2524 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2843
timestamp 1713400504
transform 1 0 2524 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2844
timestamp 1713400504
transform 1 0 2452 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2845
timestamp 1713400504
transform 1 0 2596 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2846
timestamp 1713400504
transform 1 0 2540 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2847
timestamp 1713400504
transform 1 0 2196 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2848
timestamp 1713400504
transform 1 0 2100 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2849
timestamp 1713400504
transform 1 0 2244 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2850
timestamp 1713400504
transform 1 0 2164 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2851
timestamp 1713400504
transform 1 0 1668 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2852
timestamp 1713400504
transform 1 0 1660 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2853
timestamp 1713400504
transform 1 0 1468 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2854
timestamp 1713400504
transform 1 0 1420 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2855
timestamp 1713400504
transform 1 0 1748 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2856
timestamp 1713400504
transform 1 0 1644 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2857
timestamp 1713400504
transform 1 0 1428 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2858
timestamp 1713400504
transform 1 0 1348 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2859
timestamp 1713400504
transform 1 0 1300 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2860
timestamp 1713400504
transform 1 0 1220 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2861
timestamp 1713400504
transform 1 0 1236 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2862
timestamp 1713400504
transform 1 0 1108 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2863
timestamp 1713400504
transform 1 0 1348 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2864
timestamp 1713400504
transform 1 0 1028 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2865
timestamp 1713400504
transform 1 0 1236 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2866
timestamp 1713400504
transform 1 0 1124 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2867
timestamp 1713400504
transform 1 0 1804 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2868
timestamp 1713400504
transform 1 0 1708 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2869
timestamp 1713400504
transform 1 0 2004 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2870
timestamp 1713400504
transform 1 0 1900 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2871
timestamp 1713400504
transform 1 0 2172 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2872
timestamp 1713400504
transform 1 0 2100 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2873
timestamp 1713400504
transform 1 0 2532 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2874
timestamp 1713400504
transform 1 0 2452 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2875
timestamp 1713400504
transform 1 0 2764 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2876
timestamp 1713400504
transform 1 0 2652 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2877
timestamp 1713400504
transform 1 0 2844 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2878
timestamp 1713400504
transform 1 0 2724 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2879
timestamp 1713400504
transform 1 0 2948 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2880
timestamp 1713400504
transform 1 0 2900 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2881
timestamp 1713400504
transform 1 0 2964 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2882
timestamp 1713400504
transform 1 0 2964 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2883
timestamp 1713400504
transform 1 0 2956 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2884
timestamp 1713400504
transform 1 0 2860 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2885
timestamp 1713400504
transform 1 0 2652 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2886
timestamp 1713400504
transform 1 0 2652 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2887
timestamp 1713400504
transform 1 0 2796 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2888
timestamp 1713400504
transform 1 0 2676 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2889
timestamp 1713400504
transform 1 0 2948 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2890
timestamp 1713400504
transform 1 0 2804 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2891
timestamp 1713400504
transform 1 0 2948 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2892
timestamp 1713400504
transform 1 0 2916 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2893
timestamp 1713400504
transform 1 0 2948 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2894
timestamp 1713400504
transform 1 0 2940 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2895
timestamp 1713400504
transform 1 0 2900 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2896
timestamp 1713400504
transform 1 0 2812 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2897
timestamp 1713400504
transform 1 0 2236 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2898
timestamp 1713400504
transform 1 0 2196 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2899
timestamp 1713400504
transform 1 0 2804 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2900
timestamp 1713400504
transform 1 0 2748 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2901
timestamp 1713400504
transform 1 0 2804 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2902
timestamp 1713400504
transform 1 0 2804 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2903
timestamp 1713400504
transform 1 0 2580 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2904
timestamp 1713400504
transform 1 0 2564 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2905
timestamp 1713400504
transform 1 0 2436 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2906
timestamp 1713400504
transform 1 0 2396 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2907
timestamp 1713400504
transform 1 0 2484 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2908
timestamp 1713400504
transform 1 0 2484 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2909
timestamp 1713400504
transform 1 0 2788 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2910
timestamp 1713400504
transform 1 0 2748 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2911
timestamp 1713400504
transform 1 0 2756 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2912
timestamp 1713400504
transform 1 0 2716 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2913
timestamp 1713400504
transform 1 0 2748 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2914
timestamp 1713400504
transform 1 0 2748 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2915
timestamp 1713400504
transform 1 0 2332 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2916
timestamp 1713400504
transform 1 0 2236 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2917
timestamp 1713400504
transform 1 0 2436 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2918
timestamp 1713400504
transform 1 0 2396 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2919
timestamp 1713400504
transform 1 0 2364 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2920
timestamp 1713400504
transform 1 0 2364 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2921
timestamp 1713400504
transform 1 0 2252 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2922
timestamp 1713400504
transform 1 0 2252 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2923
timestamp 1713400504
transform 1 0 2132 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2924
timestamp 1713400504
transform 1 0 2044 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2925
timestamp 1713400504
transform 1 0 2076 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2926
timestamp 1713400504
transform 1 0 2044 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2927
timestamp 1713400504
transform 1 0 1668 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2928
timestamp 1713400504
transform 1 0 1596 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2929
timestamp 1713400504
transform 1 0 1540 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2930
timestamp 1713400504
transform 1 0 1484 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2931
timestamp 1713400504
transform 1 0 1612 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2932
timestamp 1713400504
transform 1 0 1612 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2933
timestamp 1713400504
transform 1 0 1596 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2934
timestamp 1713400504
transform 1 0 1516 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2935
timestamp 1713400504
transform 1 0 1652 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2936
timestamp 1713400504
transform 1 0 1564 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2937
timestamp 1713400504
transform 1 0 1844 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2938
timestamp 1713400504
transform 1 0 1756 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2939
timestamp 1713400504
transform 1 0 1948 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2940
timestamp 1713400504
transform 1 0 1860 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2941
timestamp 1713400504
transform 1 0 1804 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2942
timestamp 1713400504
transform 1 0 1764 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2943
timestamp 1713400504
transform 1 0 2116 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2944
timestamp 1713400504
transform 1 0 2116 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2945
timestamp 1713400504
transform 1 0 2060 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2946
timestamp 1713400504
transform 1 0 2036 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2947
timestamp 1713400504
transform 1 0 1756 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2948
timestamp 1713400504
transform 1 0 1748 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2949
timestamp 1713400504
transform 1 0 1772 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2950
timestamp 1713400504
transform 1 0 1700 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2951
timestamp 1713400504
transform 1 0 1716 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2952
timestamp 1713400504
transform 1 0 1604 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2953
timestamp 1713400504
transform 1 0 1876 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2954
timestamp 1713400504
transform 1 0 1836 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2955
timestamp 1713400504
transform 1 0 1900 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2956
timestamp 1713400504
transform 1 0 1844 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2957
timestamp 1713400504
transform 1 0 2596 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2958
timestamp 1713400504
transform 1 0 2580 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2959
timestamp 1713400504
transform 1 0 2620 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2960
timestamp 1713400504
transform 1 0 2484 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2961
timestamp 1713400504
transform 1 0 2580 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2962
timestamp 1713400504
transform 1 0 2532 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2963
timestamp 1713400504
transform 1 0 2948 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2964
timestamp 1713400504
transform 1 0 2820 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2965
timestamp 1713400504
transform 1 0 1972 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2966
timestamp 1713400504
transform 1 0 1972 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2967
timestamp 1713400504
transform 1 0 2356 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2968
timestamp 1713400504
transform 1 0 2252 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2969
timestamp 1713400504
transform 1 0 2492 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2970
timestamp 1713400504
transform 1 0 2324 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2971
timestamp 1713400504
transform 1 0 2428 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_2972
timestamp 1713400504
transform 1 0 2412 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2973
timestamp 1713400504
transform 1 0 2140 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_2974
timestamp 1713400504
transform 1 0 2092 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_2975
timestamp 1713400504
transform 1 0 2052 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2976
timestamp 1713400504
transform 1 0 2380 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2977
timestamp 1713400504
transform 1 0 2380 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2978
timestamp 1713400504
transform 1 0 2356 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2979
timestamp 1713400504
transform 1 0 2340 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2980
timestamp 1713400504
transform 1 0 2028 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2981
timestamp 1713400504
transform 1 0 1932 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2982
timestamp 1713400504
transform 1 0 1956 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2983
timestamp 1713400504
transform 1 0 1940 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2984
timestamp 1713400504
transform 1 0 2196 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2985
timestamp 1713400504
transform 1 0 2092 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2986
timestamp 1713400504
transform 1 0 2020 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2987
timestamp 1713400504
transform 1 0 2108 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2988
timestamp 1713400504
transform 1 0 2076 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2989
timestamp 1713400504
transform 1 0 2316 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2990
timestamp 1713400504
transform 1 0 2196 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2991
timestamp 1713400504
transform 1 0 2156 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_2992
timestamp 1713400504
transform 1 0 2276 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2993
timestamp 1713400504
transform 1 0 2244 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2994
timestamp 1713400504
transform 1 0 2180 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_2995
timestamp 1713400504
transform 1 0 2180 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2996
timestamp 1713400504
transform 1 0 2260 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2997
timestamp 1713400504
transform 1 0 2212 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2998
timestamp 1713400504
transform 1 0 2212 0 1 105
box -2 -2 2 2
use M2_M1  M2_M1_2999
timestamp 1713400504
transform 1 0 2188 0 1 105
box -2 -2 2 2
use M2_M1  M2_M1_3000
timestamp 1713400504
transform 1 0 2140 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3001
timestamp 1713400504
transform 1 0 2140 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3002
timestamp 1713400504
transform 1 0 2180 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3003
timestamp 1713400504
transform 1 0 2164 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3004
timestamp 1713400504
transform 1 0 2084 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3005
timestamp 1713400504
transform 1 0 2180 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3006
timestamp 1713400504
transform 1 0 2076 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3007
timestamp 1713400504
transform 1 0 2276 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3008
timestamp 1713400504
transform 1 0 2148 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3009
timestamp 1713400504
transform 1 0 2132 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3010
timestamp 1713400504
transform 1 0 2068 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3011
timestamp 1713400504
transform 1 0 2932 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3012
timestamp 1713400504
transform 1 0 2924 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3013
timestamp 1713400504
transform 1 0 2988 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_3014
timestamp 1713400504
transform 1 0 2988 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3015
timestamp 1713400504
transform 1 0 2988 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3016
timestamp 1713400504
transform 1 0 2980 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_3017
timestamp 1713400504
transform 1 0 2916 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3018
timestamp 1713400504
transform 1 0 2972 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3019
timestamp 1713400504
transform 1 0 2900 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3020
timestamp 1713400504
transform 1 0 2908 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3021
timestamp 1713400504
transform 1 0 2908 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3022
timestamp 1713400504
transform 1 0 2860 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3023
timestamp 1713400504
transform 1 0 2780 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3024
timestamp 1713400504
transform 1 0 2708 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3025
timestamp 1713400504
transform 1 0 2684 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3026
timestamp 1713400504
transform 1 0 2756 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3027
timestamp 1713400504
transform 1 0 2716 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3028
timestamp 1713400504
transform 1 0 2716 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3029
timestamp 1713400504
transform 1 0 2764 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3030
timestamp 1713400504
transform 1 0 2692 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3031
timestamp 1713400504
transform 1 0 2820 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3032
timestamp 1713400504
transform 1 0 2780 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3033
timestamp 1713400504
transform 1 0 2780 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3034
timestamp 1713400504
transform 1 0 2780 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3035
timestamp 1713400504
transform 1 0 2732 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3036
timestamp 1713400504
transform 1 0 2700 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3037
timestamp 1713400504
transform 1 0 2828 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3038
timestamp 1713400504
transform 1 0 2756 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_3039
timestamp 1713400504
transform 1 0 2804 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3040
timestamp 1713400504
transform 1 0 2796 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3041
timestamp 1713400504
transform 1 0 2868 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3042
timestamp 1713400504
transform 1 0 2836 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3043
timestamp 1713400504
transform 1 0 2788 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3044
timestamp 1713400504
transform 1 0 2652 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3045
timestamp 1713400504
transform 1 0 2644 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3046
timestamp 1713400504
transform 1 0 2668 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3047
timestamp 1713400504
transform 1 0 2572 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3048
timestamp 1713400504
transform 1 0 2804 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3049
timestamp 1713400504
transform 1 0 2572 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3050
timestamp 1713400504
transform 1 0 2980 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_3051
timestamp 1713400504
transform 1 0 2980 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3052
timestamp 1713400504
transform 1 0 2740 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3053
timestamp 1713400504
transform 1 0 2708 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_3054
timestamp 1713400504
transform 1 0 2876 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3055
timestamp 1713400504
transform 1 0 2700 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3056
timestamp 1713400504
transform 1 0 2812 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3057
timestamp 1713400504
transform 1 0 2708 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3058
timestamp 1713400504
transform 1 0 2724 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3059
timestamp 1713400504
transform 1 0 2724 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_3060
timestamp 1713400504
transform 1 0 2644 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3061
timestamp 1713400504
transform 1 0 2636 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3062
timestamp 1713400504
transform 1 0 2348 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3063
timestamp 1713400504
transform 1 0 2324 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3064
timestamp 1713400504
transform 1 0 2012 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3065
timestamp 1713400504
transform 1 0 2012 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3066
timestamp 1713400504
transform 1 0 2348 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3067
timestamp 1713400504
transform 1 0 2308 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3068
timestamp 1713400504
transform 1 0 2108 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3069
timestamp 1713400504
transform 1 0 1964 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3070
timestamp 1713400504
transform 1 0 268 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3071
timestamp 1713400504
transform 1 0 268 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3072
timestamp 1713400504
transform 1 0 204 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3073
timestamp 1713400504
transform 1 0 196 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3074
timestamp 1713400504
transform 1 0 188 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3075
timestamp 1713400504
transform 1 0 164 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3076
timestamp 1713400504
transform 1 0 108 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3077
timestamp 1713400504
transform 1 0 76 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3078
timestamp 1713400504
transform 1 0 204 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3079
timestamp 1713400504
transform 1 0 188 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3080
timestamp 1713400504
transform 1 0 516 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3081
timestamp 1713400504
transform 1 0 388 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3082
timestamp 1713400504
transform 1 0 388 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3083
timestamp 1713400504
transform 1 0 676 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3084
timestamp 1713400504
transform 1 0 476 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3085
timestamp 1713400504
transform 1 0 388 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3086
timestamp 1713400504
transform 1 0 468 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3087
timestamp 1713400504
transform 1 0 428 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3088
timestamp 1713400504
transform 1 0 228 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3089
timestamp 1713400504
transform 1 0 460 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3090
timestamp 1713400504
transform 1 0 220 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3091
timestamp 1713400504
transform 1 0 172 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3092
timestamp 1713400504
transform 1 0 452 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3093
timestamp 1713400504
transform 1 0 316 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3094
timestamp 1713400504
transform 1 0 316 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3095
timestamp 1713400504
transform 1 0 508 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3096
timestamp 1713400504
transform 1 0 164 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3097
timestamp 1713400504
transform 1 0 164 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3098
timestamp 1713400504
transform 1 0 68 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3099
timestamp 1713400504
transform 1 0 2964 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3100
timestamp 1713400504
transform 1 0 2812 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3101
timestamp 1713400504
transform 1 0 2436 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3102
timestamp 1713400504
transform 1 0 2436 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3103
timestamp 1713400504
transform 1 0 2404 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3104
timestamp 1713400504
transform 1 0 2356 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3105
timestamp 1713400504
transform 1 0 2292 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_3106
timestamp 1713400504
transform 1 0 2956 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3107
timestamp 1713400504
transform 1 0 2876 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3108
timestamp 1713400504
transform 1 0 3004 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3109
timestamp 1713400504
transform 1 0 2988 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3110
timestamp 1713400504
transform 1 0 3004 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3111
timestamp 1713400504
transform 1 0 2996 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3112
timestamp 1713400504
transform 1 0 2612 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3113
timestamp 1713400504
transform 1 0 3004 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3114
timestamp 1713400504
transform 1 0 2876 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3115
timestamp 1713400504
transform 1 0 2852 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3116
timestamp 1713400504
transform 1 0 2732 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3117
timestamp 1713400504
transform 1 0 2708 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3118
timestamp 1713400504
transform 1 0 2580 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3119
timestamp 1713400504
transform 1 0 3020 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3120
timestamp 1713400504
transform 1 0 2908 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3121
timestamp 1713400504
transform 1 0 3020 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3122
timestamp 1713400504
transform 1 0 2892 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3123
timestamp 1713400504
transform 1 0 3004 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3124
timestamp 1713400504
transform 1 0 2980 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3125
timestamp 1713400504
transform 1 0 2900 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3126
timestamp 1713400504
transform 1 0 2788 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3127
timestamp 1713400504
transform 1 0 2684 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3128
timestamp 1713400504
transform 1 0 2548 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3129
timestamp 1713400504
transform 1 0 2532 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3130
timestamp 1713400504
transform 1 0 2588 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3131
timestamp 1713400504
transform 1 0 2564 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3132
timestamp 1713400504
transform 1 0 2532 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3133
timestamp 1713400504
transform 1 0 2132 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3134
timestamp 1713400504
transform 1 0 2092 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3135
timestamp 1713400504
transform 1 0 1884 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3136
timestamp 1713400504
transform 1 0 1884 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3137
timestamp 1713400504
transform 1 0 1932 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3138
timestamp 1713400504
transform 1 0 1788 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3139
timestamp 1713400504
transform 1 0 1748 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3140
timestamp 1713400504
transform 1 0 1836 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3141
timestamp 1713400504
transform 1 0 1812 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3142
timestamp 1713400504
transform 1 0 1756 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3143
timestamp 1713400504
transform 1 0 1164 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3144
timestamp 1713400504
transform 1 0 1260 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3145
timestamp 1713400504
transform 1 0 1060 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3146
timestamp 1713400504
transform 1 0 1060 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3147
timestamp 1713400504
transform 1 0 1148 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3148
timestamp 1713400504
transform 1 0 1148 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3149
timestamp 1713400504
transform 1 0 1484 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3150
timestamp 1713400504
transform 1 0 1252 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3151
timestamp 1713400504
transform 1 0 1188 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3152
timestamp 1713400504
transform 1 0 1380 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3153
timestamp 1713400504
transform 1 0 1380 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3154
timestamp 1713400504
transform 1 0 1356 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3155
timestamp 1713400504
transform 1 0 1700 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3156
timestamp 1713400504
transform 1 0 1668 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3157
timestamp 1713400504
transform 1 0 1556 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3158
timestamp 1713400504
transform 1 0 1524 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3159
timestamp 1713400504
transform 1 0 1540 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3160
timestamp 1713400504
transform 1 0 1452 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3161
timestamp 1713400504
transform 1 0 1404 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3162
timestamp 1713400504
transform 1 0 1692 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3163
timestamp 1713400504
transform 1 0 1564 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_3164
timestamp 1713400504
transform 1 0 1556 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3165
timestamp 1713400504
transform 1 0 2300 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3166
timestamp 1713400504
transform 1 0 2092 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3167
timestamp 1713400504
transform 1 0 1756 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3168
timestamp 1713400504
transform 1 0 1716 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3169
timestamp 1713400504
transform 1 0 2244 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3170
timestamp 1713400504
transform 1 0 1876 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3171
timestamp 1713400504
transform 1 0 2292 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3172
timestamp 1713400504
transform 1 0 2220 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3173
timestamp 1713400504
transform 1 0 2956 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3174
timestamp 1713400504
transform 1 0 2876 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3175
timestamp 1713400504
transform 1 0 2980 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3176
timestamp 1713400504
transform 1 0 2860 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3177
timestamp 1713400504
transform 1 0 2716 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3178
timestamp 1713400504
transform 1 0 2652 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3179
timestamp 1713400504
transform 1 0 2636 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3180
timestamp 1713400504
transform 1 0 2484 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3181
timestamp 1713400504
transform 1 0 2516 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3182
timestamp 1713400504
transform 1 0 2492 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3183
timestamp 1713400504
transform 1 0 2476 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3184
timestamp 1713400504
transform 1 0 2396 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_3185
timestamp 1713400504
transform 1 0 2548 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_3186
timestamp 1713400504
transform 1 0 2540 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3187
timestamp 1713400504
transform 1 0 2500 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3188
timestamp 1713400504
transform 1 0 2412 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_3189
timestamp 1713400504
transform 1 0 2844 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3190
timestamp 1713400504
transform 1 0 2700 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3191
timestamp 1713400504
transform 1 0 2812 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3192
timestamp 1713400504
transform 1 0 2756 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3193
timestamp 1713400504
transform 1 0 2740 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3194
timestamp 1713400504
transform 1 0 2836 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3195
timestamp 1713400504
transform 1 0 2292 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3196
timestamp 1713400504
transform 1 0 2292 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3197
timestamp 1713400504
transform 1 0 2268 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3198
timestamp 1713400504
transform 1 0 2172 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_3199
timestamp 1713400504
transform 1 0 2500 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3200
timestamp 1713400504
transform 1 0 2500 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3201
timestamp 1713400504
transform 1 0 2460 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3202
timestamp 1713400504
transform 1 0 2380 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3203
timestamp 1713400504
transform 1 0 2412 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3204
timestamp 1713400504
transform 1 0 2404 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3205
timestamp 1713400504
transform 1 0 2388 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3206
timestamp 1713400504
transform 1 0 2308 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3207
timestamp 1713400504
transform 1 0 2196 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3208
timestamp 1713400504
transform 1 0 1876 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3209
timestamp 1713400504
transform 1 0 1868 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_3210
timestamp 1713400504
transform 1 0 2076 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3211
timestamp 1713400504
transform 1 0 1956 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3212
timestamp 1713400504
transform 1 0 1948 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3213
timestamp 1713400504
transform 1 0 1764 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_3214
timestamp 1713400504
transform 1 0 2076 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3215
timestamp 1713400504
transform 1 0 1932 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3216
timestamp 1713400504
transform 1 0 1892 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3217
timestamp 1713400504
transform 1 0 1820 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_3218
timestamp 1713400504
transform 1 0 1628 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3219
timestamp 1713400504
transform 1 0 1452 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3220
timestamp 1713400504
transform 1 0 1412 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3221
timestamp 1713400504
transform 1 0 1524 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3222
timestamp 1713400504
transform 1 0 1444 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3223
timestamp 1713400504
transform 1 0 1412 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3224
timestamp 1713400504
transform 1 0 1644 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3225
timestamp 1713400504
transform 1 0 1532 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3226
timestamp 1713400504
transform 1 0 1548 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3227
timestamp 1713400504
transform 1 0 1412 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3228
timestamp 1713400504
transform 1 0 1396 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3229
timestamp 1713400504
transform 1 0 1340 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3230
timestamp 1713400504
transform 1 0 1596 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3231
timestamp 1713400504
transform 1 0 1452 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_3232
timestamp 1713400504
transform 1 0 1444 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3233
timestamp 1713400504
transform 1 0 1388 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3234
timestamp 1713400504
transform 1 0 1356 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_3235
timestamp 1713400504
transform 1 0 2444 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3236
timestamp 1713400504
transform 1 0 1788 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3237
timestamp 1713400504
transform 1 0 1660 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3238
timestamp 1713400504
transform 1 0 1540 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_3239
timestamp 1713400504
transform 1 0 1892 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3240
timestamp 1713400504
transform 1 0 1764 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3241
timestamp 1713400504
transform 1 0 1724 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3242
timestamp 1713400504
transform 1 0 1804 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3243
timestamp 1713400504
transform 1 0 1764 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3244
timestamp 1713400504
transform 1 0 1740 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3245
timestamp 1713400504
transform 1 0 2164 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3246
timestamp 1713400504
transform 1 0 2116 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3247
timestamp 1713400504
transform 1 0 1716 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_3248
timestamp 1713400504
transform 1 0 1708 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3249
timestamp 1713400504
transform 1 0 2244 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3250
timestamp 1713400504
transform 1 0 2068 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3251
timestamp 1713400504
transform 1 0 2068 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3252
timestamp 1713400504
transform 1 0 1828 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3253
timestamp 1713400504
transform 1 0 2620 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3254
timestamp 1713400504
transform 1 0 2620 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3255
timestamp 1713400504
transform 1 0 2580 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3256
timestamp 1713400504
transform 1 0 2444 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3257
timestamp 1713400504
transform 1 0 3004 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3258
timestamp 1713400504
transform 1 0 2820 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3259
timestamp 1713400504
transform 1 0 2820 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3260
timestamp 1713400504
transform 1 0 3012 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3261
timestamp 1713400504
transform 1 0 2812 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3262
timestamp 1713400504
transform 1 0 2868 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3263
timestamp 1713400504
transform 1 0 2764 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3264
timestamp 1713400504
transform 1 0 3012 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3265
timestamp 1713400504
transform 1 0 2812 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3266
timestamp 1713400504
transform 1 0 2788 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3267
timestamp 1713400504
transform 1 0 2716 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3268
timestamp 1713400504
transform 1 0 2724 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3269
timestamp 1713400504
transform 1 0 2636 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3270
timestamp 1713400504
transform 1 0 2948 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3271
timestamp 1713400504
transform 1 0 2932 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3272
timestamp 1713400504
transform 1 0 3012 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3273
timestamp 1713400504
transform 1 0 3004 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3274
timestamp 1713400504
transform 1 0 2940 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3275
timestamp 1713400504
transform 1 0 2652 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3276
timestamp 1713400504
transform 1 0 2604 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3277
timestamp 1713400504
transform 1 0 2732 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_3278
timestamp 1713400504
transform 1 0 2724 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3279
timestamp 1713400504
transform 1 0 2668 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3280
timestamp 1713400504
transform 1 0 2604 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3281
timestamp 1713400504
transform 1 0 2684 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3282
timestamp 1713400504
transform 1 0 2572 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3283
timestamp 1713400504
transform 1 0 2564 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3284
timestamp 1713400504
transform 1 0 2124 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3285
timestamp 1713400504
transform 1 0 2100 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_3286
timestamp 1713400504
transform 1 0 2100 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3287
timestamp 1713400504
transform 1 0 2068 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3288
timestamp 1713400504
transform 1 0 2020 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3289
timestamp 1713400504
transform 1 0 2404 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3290
timestamp 1713400504
transform 1 0 2324 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3291
timestamp 1713400504
transform 1 0 2180 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3292
timestamp 1713400504
transform 1 0 2140 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3293
timestamp 1713400504
transform 1 0 2060 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3294
timestamp 1713400504
transform 1 0 1940 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3295
timestamp 1713400504
transform 1 0 1940 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3296
timestamp 1713400504
transform 1 0 1844 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3297
timestamp 1713400504
transform 1 0 1844 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_3298
timestamp 1713400504
transform 1 0 1796 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3299
timestamp 1713400504
transform 1 0 1788 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_3300
timestamp 1713400504
transform 1 0 1788 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3301
timestamp 1713400504
transform 1 0 1724 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3302
timestamp 1713400504
transform 1 0 1724 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3303
timestamp 1713400504
transform 1 0 1660 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3304
timestamp 1713400504
transform 1 0 1556 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_3305
timestamp 1713400504
transform 1 0 1532 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3306
timestamp 1713400504
transform 1 0 1292 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3307
timestamp 1713400504
transform 1 0 1276 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3308
timestamp 1713400504
transform 1 0 1212 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3309
timestamp 1713400504
transform 1 0 1212 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3310
timestamp 1713400504
transform 1 0 1212 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3311
timestamp 1713400504
transform 1 0 1204 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3312
timestamp 1713400504
transform 1 0 1180 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3313
timestamp 1713400504
transform 1 0 1180 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3314
timestamp 1713400504
transform 1 0 1172 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3315
timestamp 1713400504
transform 1 0 1164 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3316
timestamp 1713400504
transform 1 0 1156 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3317
timestamp 1713400504
transform 1 0 1036 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3318
timestamp 1713400504
transform 1 0 948 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3319
timestamp 1713400504
transform 1 0 892 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3320
timestamp 1713400504
transform 1 0 884 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3321
timestamp 1713400504
transform 1 0 1956 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3322
timestamp 1713400504
transform 1 0 1892 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3323
timestamp 1713400504
transform 1 0 1860 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3324
timestamp 1713400504
transform 1 0 1860 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3325
timestamp 1713400504
transform 1 0 1828 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3326
timestamp 1713400504
transform 1 0 1732 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3327
timestamp 1713400504
transform 1 0 1620 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3328
timestamp 1713400504
transform 1 0 1620 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3329
timestamp 1713400504
transform 1 0 1572 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3330
timestamp 1713400504
transform 1 0 1308 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3331
timestamp 1713400504
transform 1 0 1292 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_3332
timestamp 1713400504
transform 1 0 1276 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3333
timestamp 1713400504
transform 1 0 1260 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3334
timestamp 1713400504
transform 1 0 1180 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3335
timestamp 1713400504
transform 1 0 1164 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3336
timestamp 1713400504
transform 1 0 1148 0 1 1955
box -2 -2 2 2
use M2_M1  M2_M1_3337
timestamp 1713400504
transform 1 0 1116 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3338
timestamp 1713400504
transform 1 0 1108 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3339
timestamp 1713400504
transform 1 0 1084 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3340
timestamp 1713400504
transform 1 0 1956 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3341
timestamp 1713400504
transform 1 0 1948 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_3342
timestamp 1713400504
transform 1 0 1940 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_3343
timestamp 1713400504
transform 1 0 1900 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3344
timestamp 1713400504
transform 1 0 1884 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3345
timestamp 1713400504
transform 1 0 1860 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3346
timestamp 1713400504
transform 1 0 1780 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3347
timestamp 1713400504
transform 1 0 1764 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3348
timestamp 1713400504
transform 1 0 1660 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3349
timestamp 1713400504
transform 1 0 1636 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3350
timestamp 1713400504
transform 1 0 1572 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3351
timestamp 1713400504
transform 1 0 1572 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3352
timestamp 1713400504
transform 1 0 1484 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3353
timestamp 1713400504
transform 1 0 1388 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3354
timestamp 1713400504
transform 1 0 1388 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3355
timestamp 1713400504
transform 1 0 1388 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3356
timestamp 1713400504
transform 1 0 1364 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3357
timestamp 1713400504
transform 1 0 1324 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3358
timestamp 1713400504
transform 1 0 1316 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3359
timestamp 1713400504
transform 1 0 1316 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3360
timestamp 1713400504
transform 1 0 1300 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3361
timestamp 1713400504
transform 1 0 2044 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_3362
timestamp 1713400504
transform 1 0 1996 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3363
timestamp 1713400504
transform 1 0 1972 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3364
timestamp 1713400504
transform 1 0 1932 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3365
timestamp 1713400504
transform 1 0 1860 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3366
timestamp 1713400504
transform 1 0 1844 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3367
timestamp 1713400504
transform 1 0 1828 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3368
timestamp 1713400504
transform 1 0 1580 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_3369
timestamp 1713400504
transform 1 0 1476 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3370
timestamp 1713400504
transform 1 0 1380 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_3371
timestamp 1713400504
transform 1 0 1372 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3372
timestamp 1713400504
transform 1 0 1372 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_3373
timestamp 1713400504
transform 1 0 1348 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_3374
timestamp 1713400504
transform 1 0 1348 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3375
timestamp 1713400504
transform 1 0 1284 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3376
timestamp 1713400504
transform 1 0 1284 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_3377
timestamp 1713400504
transform 1 0 1956 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3378
timestamp 1713400504
transform 1 0 1924 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3379
timestamp 1713400504
transform 1 0 1900 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_3380
timestamp 1713400504
transform 1 0 1884 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3381
timestamp 1713400504
transform 1 0 1868 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3382
timestamp 1713400504
transform 1 0 1844 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3383
timestamp 1713400504
transform 1 0 1836 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3384
timestamp 1713400504
transform 1 0 1796 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_3385
timestamp 1713400504
transform 1 0 1652 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3386
timestamp 1713400504
transform 1 0 1452 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3387
timestamp 1713400504
transform 1 0 1364 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3388
timestamp 1713400504
transform 1 0 1340 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3389
timestamp 1713400504
transform 1 0 2020 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3390
timestamp 1713400504
transform 1 0 1940 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3391
timestamp 1713400504
transform 1 0 1932 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_3392
timestamp 1713400504
transform 1 0 1348 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3393
timestamp 1713400504
transform 1 0 1332 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3394
timestamp 1713400504
transform 1 0 876 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3395
timestamp 1713400504
transform 1 0 812 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3396
timestamp 1713400504
transform 1 0 772 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3397
timestamp 1713400504
transform 1 0 332 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3398
timestamp 1713400504
transform 1 0 196 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3399
timestamp 1713400504
transform 1 0 1740 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3400
timestamp 1713400504
transform 1 0 1596 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3401
timestamp 1713400504
transform 1 0 1228 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3402
timestamp 1713400504
transform 1 0 844 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3403
timestamp 1713400504
transform 1 0 724 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3404
timestamp 1713400504
transform 1 0 676 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3405
timestamp 1713400504
transform 1 0 556 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3406
timestamp 1713400504
transform 1 0 556 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3407
timestamp 1713400504
transform 1 0 2844 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3408
timestamp 1713400504
transform 1 0 2708 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3409
timestamp 1713400504
transform 1 0 2620 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3410
timestamp 1713400504
transform 1 0 1564 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3411
timestamp 1713400504
transform 1 0 1340 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3412
timestamp 1713400504
transform 1 0 1116 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3413
timestamp 1713400504
transform 1 0 1092 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3414
timestamp 1713400504
transform 1 0 1084 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3415
timestamp 1713400504
transform 1 0 1076 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3416
timestamp 1713400504
transform 1 0 1052 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3417
timestamp 1713400504
transform 1 0 924 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3418
timestamp 1713400504
transform 1 0 788 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3419
timestamp 1713400504
transform 1 0 2492 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3420
timestamp 1713400504
transform 1 0 2492 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3421
timestamp 1713400504
transform 1 0 1700 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3422
timestamp 1713400504
transform 1 0 1252 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3423
timestamp 1713400504
transform 1 0 1148 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3424
timestamp 1713400504
transform 1 0 1060 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3425
timestamp 1713400504
transform 1 0 1044 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3426
timestamp 1713400504
transform 1 0 1012 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3427
timestamp 1713400504
transform 1 0 972 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3428
timestamp 1713400504
transform 1 0 2508 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3429
timestamp 1713400504
transform 1 0 2500 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3430
timestamp 1713400504
transform 1 0 2108 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3431
timestamp 1713400504
transform 1 0 1660 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3432
timestamp 1713400504
transform 1 0 1220 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3433
timestamp 1713400504
transform 1 0 788 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3434
timestamp 1713400504
transform 1 0 764 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3435
timestamp 1713400504
transform 1 0 748 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3436
timestamp 1713400504
transform 1 0 164 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3437
timestamp 1713400504
transform 1 0 164 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3438
timestamp 1713400504
transform 1 0 1428 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3439
timestamp 1713400504
transform 1 0 1404 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3440
timestamp 1713400504
transform 1 0 1180 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3441
timestamp 1713400504
transform 1 0 756 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3442
timestamp 1713400504
transform 1 0 716 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3443
timestamp 1713400504
transform 1 0 708 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3444
timestamp 1713400504
transform 1 0 692 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_3445
timestamp 1713400504
transform 1 0 228 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3446
timestamp 1713400504
transform 1 0 196 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3447
timestamp 1713400504
transform 1 0 2764 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3448
timestamp 1713400504
transform 1 0 2732 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3449
timestamp 1713400504
transform 1 0 1524 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3450
timestamp 1713400504
transform 1 0 1196 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3451
timestamp 1713400504
transform 1 0 1044 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3452
timestamp 1713400504
transform 1 0 988 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3453
timestamp 1713400504
transform 1 0 892 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3454
timestamp 1713400504
transform 1 0 852 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3455
timestamp 1713400504
transform 1 0 236 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3456
timestamp 1713400504
transform 1 0 204 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3457
timestamp 1713400504
transform 1 0 2860 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3458
timestamp 1713400504
transform 1 0 2820 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_3459
timestamp 1713400504
transform 1 0 2748 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3460
timestamp 1713400504
transform 1 0 1404 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3461
timestamp 1713400504
transform 1 0 1164 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3462
timestamp 1713400504
transform 1 0 956 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3463
timestamp 1713400504
transform 1 0 796 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3464
timestamp 1713400504
transform 1 0 796 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3465
timestamp 1713400504
transform 1 0 572 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3466
timestamp 1713400504
transform 1 0 516 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3467
timestamp 1713400504
transform 1 0 2172 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3468
timestamp 1713400504
transform 1 0 1412 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3469
timestamp 1713400504
transform 1 0 1276 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3470
timestamp 1713400504
transform 1 0 1276 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3471
timestamp 1713400504
transform 1 0 1172 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3472
timestamp 1713400504
transform 1 0 996 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3473
timestamp 1713400504
transform 1 0 972 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3474
timestamp 1713400504
transform 1 0 708 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3475
timestamp 1713400504
transform 1 0 684 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3476
timestamp 1713400504
transform 1 0 1500 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3477
timestamp 1713400504
transform 1 0 1340 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3478
timestamp 1713400504
transform 1 0 1244 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3479
timestamp 1713400504
transform 1 0 1108 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3480
timestamp 1713400504
transform 1 0 940 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3481
timestamp 1713400504
transform 1 0 932 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3482
timestamp 1713400504
transform 1 0 884 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3483
timestamp 1713400504
transform 1 0 652 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3484
timestamp 1713400504
transform 1 0 2556 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3485
timestamp 1713400504
transform 1 0 2516 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3486
timestamp 1713400504
transform 1 0 2388 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3487
timestamp 1713400504
transform 1 0 1452 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3488
timestamp 1713400504
transform 1 0 1428 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3489
timestamp 1713400504
transform 1 0 1428 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3490
timestamp 1713400504
transform 1 0 1388 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3491
timestamp 1713400504
transform 1 0 1260 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3492
timestamp 1713400504
transform 1 0 1260 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3493
timestamp 1713400504
transform 1 0 1220 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3494
timestamp 1713400504
transform 1 0 1172 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3495
timestamp 1713400504
transform 1 0 1156 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3496
timestamp 1713400504
transform 1 0 1140 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3497
timestamp 1713400504
transform 1 0 1076 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3498
timestamp 1713400504
transform 1 0 1060 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3499
timestamp 1713400504
transform 1 0 2556 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3500
timestamp 1713400504
transform 1 0 2452 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3501
timestamp 1713400504
transform 1 0 2148 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3502
timestamp 1713400504
transform 1 0 1492 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3503
timestamp 1713400504
transform 1 0 1148 0 1 385
box -2 -2 2 2
use M2_M1  M2_M1_3504
timestamp 1713400504
transform 1 0 1124 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3505
timestamp 1713400504
transform 1 0 1124 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3506
timestamp 1713400504
transform 1 0 1124 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3507
timestamp 1713400504
transform 1 0 1084 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3508
timestamp 1713400504
transform 1 0 996 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3509
timestamp 1713400504
transform 1 0 1892 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3510
timestamp 1713400504
transform 1 0 1860 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3511
timestamp 1713400504
transform 1 0 1660 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3512
timestamp 1713400504
transform 1 0 1516 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3513
timestamp 1713400504
transform 1 0 1308 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3514
timestamp 1713400504
transform 1 0 1116 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3515
timestamp 1713400504
transform 1 0 1076 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3516
timestamp 1713400504
transform 1 0 1076 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3517
timestamp 1713400504
transform 1 0 1036 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3518
timestamp 1713400504
transform 1 0 996 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3519
timestamp 1713400504
transform 1 0 1956 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3520
timestamp 1713400504
transform 1 0 1724 0 1 2755
box -2 -2 2 2
use M2_M1  M2_M1_3521
timestamp 1713400504
transform 1 0 1676 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3522
timestamp 1713400504
transform 1 0 1628 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3523
timestamp 1713400504
transform 1 0 1500 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3524
timestamp 1713400504
transform 1 0 1236 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3525
timestamp 1713400504
transform 1 0 1012 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3526
timestamp 1713400504
transform 1 0 988 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3527
timestamp 1713400504
transform 1 0 932 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3528
timestamp 1713400504
transform 1 0 924 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3529
timestamp 1713400504
transform 1 0 692 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3530
timestamp 1713400504
transform 1 0 580 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3531
timestamp 1713400504
transform 1 0 1836 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3532
timestamp 1713400504
transform 1 0 1836 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3533
timestamp 1713400504
transform 1 0 1604 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3534
timestamp 1713400504
transform 1 0 1244 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3535
timestamp 1713400504
transform 1 0 1140 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3536
timestamp 1713400504
transform 1 0 1140 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_3537
timestamp 1713400504
transform 1 0 1108 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3538
timestamp 1713400504
transform 1 0 1028 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_3539
timestamp 1713400504
transform 1 0 1020 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3540
timestamp 1713400504
transform 1 0 964 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3541
timestamp 1713400504
transform 1 0 860 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3542
timestamp 1713400504
transform 1 0 1476 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3543
timestamp 1713400504
transform 1 0 1356 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3544
timestamp 1713400504
transform 1 0 1156 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3545
timestamp 1713400504
transform 1 0 1100 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3546
timestamp 1713400504
transform 1 0 1092 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3547
timestamp 1713400504
transform 1 0 1068 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3548
timestamp 1713400504
transform 1 0 1068 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3549
timestamp 1713400504
transform 1 0 1004 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3550
timestamp 1713400504
transform 1 0 860 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3551
timestamp 1713400504
transform 1 0 604 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3552
timestamp 1713400504
transform 1 0 556 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3553
timestamp 1713400504
transform 1 0 532 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3554
timestamp 1713400504
transform 1 0 1492 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3555
timestamp 1713400504
transform 1 0 1436 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3556
timestamp 1713400504
transform 1 0 1388 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3557
timestamp 1713400504
transform 1 0 1212 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3558
timestamp 1713400504
transform 1 0 1068 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3559
timestamp 1713400504
transform 1 0 924 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3560
timestamp 1713400504
transform 1 0 884 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3561
timestamp 1713400504
transform 1 0 588 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3562
timestamp 1713400504
transform 1 0 580 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3563
timestamp 1713400504
transform 1 0 556 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3564
timestamp 1713400504
transform 1 0 1316 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3565
timestamp 1713400504
transform 1 0 1316 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3566
timestamp 1713400504
transform 1 0 1244 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3567
timestamp 1713400504
transform 1 0 1132 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3568
timestamp 1713400504
transform 1 0 852 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3569
timestamp 1713400504
transform 1 0 852 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3570
timestamp 1713400504
transform 1 0 500 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3571
timestamp 1713400504
transform 1 0 476 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3572
timestamp 1713400504
transform 1 0 460 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3573
timestamp 1713400504
transform 1 0 1476 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3574
timestamp 1713400504
transform 1 0 1476 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3575
timestamp 1713400504
transform 1 0 1364 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3576
timestamp 1713400504
transform 1 0 1332 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3577
timestamp 1713400504
transform 1 0 1332 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3578
timestamp 1713400504
transform 1 0 1292 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3579
timestamp 1713400504
transform 1 0 1172 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3580
timestamp 1713400504
transform 1 0 988 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3581
timestamp 1713400504
transform 1 0 916 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3582
timestamp 1713400504
transform 1 0 876 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3583
timestamp 1713400504
transform 1 0 876 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3584
timestamp 1713400504
transform 1 0 756 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3585
timestamp 1713400504
transform 1 0 1476 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3586
timestamp 1713400504
transform 1 0 1420 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3587
timestamp 1713400504
transform 1 0 1420 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3588
timestamp 1713400504
transform 1 0 1420 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3589
timestamp 1713400504
transform 1 0 1268 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3590
timestamp 1713400504
transform 1 0 1116 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3591
timestamp 1713400504
transform 1 0 940 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3592
timestamp 1713400504
transform 1 0 900 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3593
timestamp 1713400504
transform 1 0 836 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3594
timestamp 1713400504
transform 1 0 828 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3595
timestamp 1713400504
transform 1 0 1492 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3596
timestamp 1713400504
transform 1 0 1484 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3597
timestamp 1713400504
transform 1 0 1484 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3598
timestamp 1713400504
transform 1 0 1460 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3599
timestamp 1713400504
transform 1 0 1420 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3600
timestamp 1713400504
transform 1 0 972 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3601
timestamp 1713400504
transform 1 0 820 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3602
timestamp 1713400504
transform 1 0 804 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3603
timestamp 1713400504
transform 1 0 756 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3604
timestamp 1713400504
transform 1 0 668 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3605
timestamp 1713400504
transform 1 0 1668 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3606
timestamp 1713400504
transform 1 0 1588 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3607
timestamp 1713400504
transform 1 0 1388 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3608
timestamp 1713400504
transform 1 0 796 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3609
timestamp 1713400504
transform 1 0 788 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3610
timestamp 1713400504
transform 1 0 772 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3611
timestamp 1713400504
transform 1 0 740 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3612
timestamp 1713400504
transform 1 0 716 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3613
timestamp 1713400504
transform 1 0 716 0 1 1895
box -2 -2 2 2
use M2_M1  M2_M1_3614
timestamp 1713400504
transform 1 0 636 0 1 1895
box -2 -2 2 2
use M2_M1  M2_M1_3615
timestamp 1713400504
transform 1 0 636 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3616
timestamp 1713400504
transform 1 0 1748 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3617
timestamp 1713400504
transform 1 0 1604 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3618
timestamp 1713400504
transform 1 0 1580 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3619
timestamp 1713400504
transform 1 0 1580 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3620
timestamp 1713400504
transform 1 0 1196 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3621
timestamp 1713400504
transform 1 0 972 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3622
timestamp 1713400504
transform 1 0 916 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3623
timestamp 1713400504
transform 1 0 844 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3624
timestamp 1713400504
transform 1 0 580 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3625
timestamp 1713400504
transform 1 0 564 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3626
timestamp 1713400504
transform 1 0 1700 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_3627
timestamp 1713400504
transform 1 0 1700 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3628
timestamp 1713400504
transform 1 0 1644 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3629
timestamp 1713400504
transform 1 0 1644 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3630
timestamp 1713400504
transform 1 0 1132 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3631
timestamp 1713400504
transform 1 0 908 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3632
timestamp 1713400504
transform 1 0 828 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3633
timestamp 1713400504
transform 1 0 724 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3634
timestamp 1713400504
transform 1 0 724 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3635
timestamp 1713400504
transform 1 0 692 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3636
timestamp 1713400504
transform 1 0 1764 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3637
timestamp 1713400504
transform 1 0 1396 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3638
timestamp 1713400504
transform 1 0 220 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3639
timestamp 1713400504
transform 1 0 68 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3640
timestamp 1713400504
transform 1 0 2804 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_3641
timestamp 1713400504
transform 1 0 1804 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3642
timestamp 1713400504
transform 1 0 1652 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_3643
timestamp 1713400504
transform 1 0 2020 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3644
timestamp 1713400504
transform 1 0 1964 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3645
timestamp 1713400504
transform 1 0 1812 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3646
timestamp 1713400504
transform 1 0 1564 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3647
timestamp 1713400504
transform 1 0 1540 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3648
timestamp 1713400504
transform 1 0 1788 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3649
timestamp 1713400504
transform 1 0 1756 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3650
timestamp 1713400504
transform 1 0 1700 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3651
timestamp 1713400504
transform 1 0 1820 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3652
timestamp 1713400504
transform 1 0 1876 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3653
timestamp 1713400504
transform 1 0 2932 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3654
timestamp 1713400504
transform 1 0 2852 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3655
timestamp 1713400504
transform 1 0 2772 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_3656
timestamp 1713400504
transform 1 0 2852 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3657
timestamp 1713400504
transform 1 0 2956 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3658
timestamp 1713400504
transform 1 0 2820 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_3659
timestamp 1713400504
transform 1 0 2812 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3660
timestamp 1713400504
transform 1 0 2788 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3661
timestamp 1713400504
transform 1 0 2620 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3662
timestamp 1713400504
transform 1 0 2580 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3663
timestamp 1713400504
transform 1 0 2988 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3664
timestamp 1713400504
transform 1 0 2924 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3665
timestamp 1713400504
transform 1 0 2628 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3666
timestamp 1713400504
transform 1 0 2556 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3667
timestamp 1713400504
transform 1 0 2948 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3668
timestamp 1713400504
transform 1 0 2948 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_3669
timestamp 1713400504
transform 1 0 2900 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3670
timestamp 1713400504
transform 1 0 2804 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3671
timestamp 1713400504
transform 1 0 2708 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3672
timestamp 1713400504
transform 1 0 2612 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3673
timestamp 1713400504
transform 1 0 2556 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3674
timestamp 1713400504
transform 1 0 2964 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3675
timestamp 1713400504
transform 1 0 2892 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_3676
timestamp 1713400504
transform 1 0 2756 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3677
timestamp 1713400504
transform 1 0 2652 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3678
timestamp 1713400504
transform 1 0 2548 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_3679
timestamp 1713400504
transform 1 0 324 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3680
timestamp 1713400504
transform 1 0 252 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3681
timestamp 1713400504
transform 1 0 444 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3682
timestamp 1713400504
transform 1 0 276 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3683
timestamp 1713400504
transform 1 0 276 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3684
timestamp 1713400504
transform 1 0 212 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3685
timestamp 1713400504
transform 1 0 276 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3686
timestamp 1713400504
transform 1 0 308 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3687
timestamp 1713400504
transform 1 0 228 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3688
timestamp 1713400504
transform 1 0 292 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3689
timestamp 1713400504
transform 1 0 2988 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3690
timestamp 1713400504
transform 1 0 1604 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_3691
timestamp 1713400504
transform 1 0 2692 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3692
timestamp 1713400504
transform 1 0 2164 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3693
timestamp 1713400504
transform 1 0 732 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_0
timestamp 1713400504
transform 1 0 2948 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1
timestamp 1713400504
transform 1 0 2820 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2
timestamp 1713400504
transform 1 0 2908 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3
timestamp 1713400504
transform 1 0 2796 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_4
timestamp 1713400504
transform 1 0 300 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5
timestamp 1713400504
transform 1 0 260 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_6
timestamp 1713400504
transform 1 0 164 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_7
timestamp 1713400504
transform 1 0 164 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_8
timestamp 1713400504
transform 1 0 132 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_9
timestamp 1713400504
transform 1 0 132 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_10
timestamp 1713400504
transform 1 0 124 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_11
timestamp 1713400504
transform 1 0 164 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_12
timestamp 1713400504
transform 1 0 156 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_13
timestamp 1713400504
transform 1 0 84 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_14
timestamp 1713400504
transform 1 0 76 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_15
timestamp 1713400504
transform 1 0 452 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_16
timestamp 1713400504
transform 1 0 252 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_17
timestamp 1713400504
transform 1 0 956 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_18
timestamp 1713400504
transform 1 0 780 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_19
timestamp 1713400504
transform 1 0 620 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_20
timestamp 1713400504
transform 1 0 468 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_21
timestamp 1713400504
transform 1 0 980 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_22
timestamp 1713400504
transform 1 0 980 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_23
timestamp 1713400504
transform 1 0 916 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_24
timestamp 1713400504
transform 1 0 884 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_25
timestamp 1713400504
transform 1 0 756 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_26
timestamp 1713400504
transform 1 0 668 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_27
timestamp 1713400504
transform 1 0 620 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_28
timestamp 1713400504
transform 1 0 2620 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_29
timestamp 1713400504
transform 1 0 2556 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_30
timestamp 1713400504
transform 1 0 2484 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_31
timestamp 1713400504
transform 1 0 2204 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_32
timestamp 1713400504
transform 1 0 2508 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_33
timestamp 1713400504
transform 1 0 2476 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_34
timestamp 1713400504
transform 1 0 2420 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_35
timestamp 1713400504
transform 1 0 2332 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_36
timestamp 1713400504
transform 1 0 2564 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_37
timestamp 1713400504
transform 1 0 2500 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_38
timestamp 1713400504
transform 1 0 2396 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_39
timestamp 1713400504
transform 1 0 2260 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_40
timestamp 1713400504
transform 1 0 2836 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_41
timestamp 1713400504
transform 1 0 2596 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_42
timestamp 1713400504
transform 1 0 2444 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_43
timestamp 1713400504
transform 1 0 2396 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_44
timestamp 1713400504
transform 1 0 204 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_45
timestamp 1713400504
transform 1 0 100 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_46
timestamp 1713400504
transform 1 0 972 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_47
timestamp 1713400504
transform 1 0 892 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_48
timestamp 1713400504
transform 1 0 1052 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_49
timestamp 1713400504
transform 1 0 964 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_50
timestamp 1713400504
transform 1 0 940 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_51
timestamp 1713400504
transform 1 0 868 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_52
timestamp 1713400504
transform 1 0 820 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_53
timestamp 1713400504
transform 1 0 740 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_54
timestamp 1713400504
transform 1 0 700 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_55
timestamp 1713400504
transform 1 0 580 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_56
timestamp 1713400504
transform 1 0 812 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_57
timestamp 1713400504
transform 1 0 492 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_58
timestamp 1713400504
transform 1 0 652 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_59
timestamp 1713400504
transform 1 0 508 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_60
timestamp 1713400504
transform 1 0 516 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_61
timestamp 1713400504
transform 1 0 444 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_62
timestamp 1713400504
transform 1 0 492 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_63
timestamp 1713400504
transform 1 0 428 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_64
timestamp 1713400504
transform 1 0 340 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_65
timestamp 1713400504
transform 1 0 508 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_66
timestamp 1713400504
transform 1 0 420 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_67
timestamp 1713400504
transform 1 0 284 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_68
timestamp 1713400504
transform 1 0 196 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_69
timestamp 1713400504
transform 1 0 316 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_70
timestamp 1713400504
transform 1 0 244 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_71
timestamp 1713400504
transform 1 0 300 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_72
timestamp 1713400504
transform 1 0 228 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_73
timestamp 1713400504
transform 1 0 276 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_74
timestamp 1713400504
transform 1 0 204 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_75
timestamp 1713400504
transform 1 0 204 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_76
timestamp 1713400504
transform 1 0 92 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_77
timestamp 1713400504
transform 1 0 340 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_78
timestamp 1713400504
transform 1 0 244 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_79
timestamp 1713400504
transform 1 0 116 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_80
timestamp 1713400504
transform 1 0 68 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_81
timestamp 1713400504
transform 1 0 116 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_82
timestamp 1713400504
transform 1 0 116 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_83
timestamp 1713400504
transform 1 0 244 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_84
timestamp 1713400504
transform 1 0 244 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_85
timestamp 1713400504
transform 1 0 236 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_86
timestamp 1713400504
transform 1 0 172 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_87
timestamp 1713400504
transform 1 0 164 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_88
timestamp 1713400504
transform 1 0 100 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_89
timestamp 1713400504
transform 1 0 308 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_90
timestamp 1713400504
transform 1 0 156 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_91
timestamp 1713400504
transform 1 0 356 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_92
timestamp 1713400504
transform 1 0 324 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_93
timestamp 1713400504
transform 1 0 620 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_94
timestamp 1713400504
transform 1 0 548 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_95
timestamp 1713400504
transform 1 0 468 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_96
timestamp 1713400504
transform 1 0 436 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_97
timestamp 1713400504
transform 1 0 388 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_98
timestamp 1713400504
transform 1 0 388 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_99
timestamp 1713400504
transform 1 0 1124 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_100
timestamp 1713400504
transform 1 0 1084 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_101
timestamp 1713400504
transform 1 0 1948 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_102
timestamp 1713400504
transform 1 0 1916 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_103
timestamp 1713400504
transform 1 0 2340 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_104
timestamp 1713400504
transform 1 0 2260 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_105
timestamp 1713400504
transform 1 0 2196 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_106
timestamp 1713400504
transform 1 0 2092 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_107
timestamp 1713400504
transform 1 0 2092 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_108
timestamp 1713400504
transform 1 0 2028 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_109
timestamp 1713400504
transform 1 0 2004 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_110
timestamp 1713400504
transform 1 0 2228 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_111
timestamp 1713400504
transform 1 0 2124 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_112
timestamp 1713400504
transform 1 0 2356 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_113
timestamp 1713400504
transform 1 0 2268 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_114
timestamp 1713400504
transform 1 0 2268 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_115
timestamp 1713400504
transform 1 0 2236 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_116
timestamp 1713400504
transform 1 0 1996 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_117
timestamp 1713400504
transform 1 0 2340 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_118
timestamp 1713400504
transform 1 0 2252 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_119
timestamp 1713400504
transform 1 0 1964 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_120
timestamp 1713400504
transform 1 0 2260 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_121
timestamp 1713400504
transform 1 0 2148 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_122
timestamp 1713400504
transform 1 0 2004 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_123
timestamp 1713400504
transform 1 0 1956 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_124
timestamp 1713400504
transform 1 0 1932 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_125
timestamp 1713400504
transform 1 0 1892 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_126
timestamp 1713400504
transform 1 0 1892 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_127
timestamp 1713400504
transform 1 0 2212 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_128
timestamp 1713400504
transform 1 0 2140 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_129
timestamp 1713400504
transform 1 0 2076 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_130
timestamp 1713400504
transform 1 0 1980 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_131
timestamp 1713400504
transform 1 0 1900 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_132
timestamp 1713400504
transform 1 0 2060 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_133
timestamp 1713400504
transform 1 0 1980 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_134
timestamp 1713400504
transform 1 0 1924 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_135
timestamp 1713400504
transform 1 0 2180 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_136
timestamp 1713400504
transform 1 0 2124 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_137
timestamp 1713400504
transform 1 0 2108 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_138
timestamp 1713400504
transform 1 0 2068 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_139
timestamp 1713400504
transform 1 0 2044 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_140
timestamp 1713400504
transform 1 0 348 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_141
timestamp 1713400504
transform 1 0 316 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_142
timestamp 1713400504
transform 1 0 476 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_143
timestamp 1713400504
transform 1 0 348 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_144
timestamp 1713400504
transform 1 0 2564 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_145
timestamp 1713400504
transform 1 0 2508 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_146
timestamp 1713400504
transform 1 0 1500 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_147
timestamp 1713400504
transform 1 0 2980 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_148
timestamp 1713400504
transform 1 0 2804 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_149
timestamp 1713400504
transform 1 0 2500 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_150
timestamp 1713400504
transform 1 0 2124 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_151
timestamp 1713400504
transform 1 0 1820 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_152
timestamp 1713400504
transform 1 0 2868 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_153
timestamp 1713400504
transform 1 0 2708 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_154
timestamp 1713400504
transform 1 0 1404 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_155
timestamp 1713400504
transform 1 0 2916 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_156
timestamp 1713400504
transform 1 0 2828 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_157
timestamp 1713400504
transform 1 0 2772 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_158
timestamp 1713400504
transform 1 0 2772 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_159
timestamp 1713400504
transform 1 0 1812 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_160
timestamp 1713400504
transform 1 0 1948 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_161
timestamp 1713400504
transform 1 0 1844 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_162
timestamp 1713400504
transform 1 0 3012 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_163
timestamp 1713400504
transform 1 0 3012 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_164
timestamp 1713400504
transform 1 0 1748 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_165
timestamp 1713400504
transform 1 0 1676 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_166
timestamp 1713400504
transform 1 0 2788 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_167
timestamp 1713400504
transform 1 0 2644 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_168
timestamp 1713400504
transform 1 0 2220 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_169
timestamp 1713400504
transform 1 0 2652 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_170
timestamp 1713400504
transform 1 0 2460 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_171
timestamp 1713400504
transform 1 0 2452 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_172
timestamp 1713400504
transform 1 0 1772 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_173
timestamp 1713400504
transform 1 0 1756 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_174
timestamp 1713400504
transform 1 0 1516 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_175
timestamp 1713400504
transform 1 0 1652 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_176
timestamp 1713400504
transform 1 0 1548 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_177
timestamp 1713400504
transform 1 0 1644 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_178
timestamp 1713400504
transform 1 0 1556 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_179
timestamp 1713400504
transform 1 0 1500 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_180
timestamp 1713400504
transform 1 0 1492 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_181
timestamp 1713400504
transform 1 0 1460 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_182
timestamp 1713400504
transform 1 0 1612 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_183
timestamp 1713400504
transform 1 0 1396 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_184
timestamp 1713400504
transform 1 0 1340 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_185
timestamp 1713400504
transform 1 0 1268 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_186
timestamp 1713400504
transform 1 0 1548 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_187
timestamp 1713400504
transform 1 0 1468 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_188
timestamp 1713400504
transform 1 0 1436 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_189
timestamp 1713400504
transform 1 0 1412 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_190
timestamp 1713400504
transform 1 0 1412 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_191
timestamp 1713400504
transform 1 0 1348 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_192
timestamp 1713400504
transform 1 0 1284 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_193
timestamp 1713400504
transform 1 0 1236 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_194
timestamp 1713400504
transform 1 0 172 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_195
timestamp 1713400504
transform 1 0 100 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_196
timestamp 1713400504
transform 1 0 1212 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_197
timestamp 1713400504
transform 1 0 1188 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_198
timestamp 1713400504
transform 1 0 2428 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_199
timestamp 1713400504
transform 1 0 2220 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_200
timestamp 1713400504
transform 1 0 2188 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_201
timestamp 1713400504
transform 1 0 2188 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_202
timestamp 1713400504
transform 1 0 2180 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_203
timestamp 1713400504
transform 1 0 1692 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_204
timestamp 1713400504
transform 1 0 2628 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_205
timestamp 1713400504
transform 1 0 2596 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_206
timestamp 1713400504
transform 1 0 2604 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_207
timestamp 1713400504
transform 1 0 2564 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_208
timestamp 1713400504
transform 1 0 2028 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_209
timestamp 1713400504
transform 1 0 1964 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_210
timestamp 1713400504
transform 1 0 1868 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_211
timestamp 1713400504
transform 1 0 1756 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_212
timestamp 1713400504
transform 1 0 1732 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_213
timestamp 1713400504
transform 1 0 1604 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_214
timestamp 1713400504
transform 1 0 1548 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_215
timestamp 1713400504
transform 1 0 1500 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_216
timestamp 1713400504
transform 1 0 1700 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_217
timestamp 1713400504
transform 1 0 1692 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_218
timestamp 1713400504
transform 1 0 1532 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_219
timestamp 1713400504
transform 1 0 1444 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_220
timestamp 1713400504
transform 1 0 1436 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_221
timestamp 1713400504
transform 1 0 2012 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_222
timestamp 1713400504
transform 1 0 1932 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_223
timestamp 1713400504
transform 1 0 1908 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_224
timestamp 1713400504
transform 1 0 1804 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_225
timestamp 1713400504
transform 1 0 1804 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_226
timestamp 1713400504
transform 1 0 1668 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_227
timestamp 1713400504
transform 1 0 1508 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_228
timestamp 1713400504
transform 1 0 1508 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_229
timestamp 1713400504
transform 1 0 1412 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_230
timestamp 1713400504
transform 1 0 1316 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_231
timestamp 1713400504
transform 1 0 1260 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_232
timestamp 1713400504
transform 1 0 1260 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_233
timestamp 1713400504
transform 1 0 1228 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_234
timestamp 1713400504
transform 1 0 1972 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_235
timestamp 1713400504
transform 1 0 1972 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_236
timestamp 1713400504
transform 1 0 1932 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_237
timestamp 1713400504
transform 1 0 1876 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_238
timestamp 1713400504
transform 1 0 1772 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_239
timestamp 1713400504
transform 1 0 1652 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_240
timestamp 1713400504
transform 1 0 1204 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_241
timestamp 1713400504
transform 1 0 1140 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_242
timestamp 1713400504
transform 1 0 1132 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_243
timestamp 1713400504
transform 1 0 1036 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_244
timestamp 1713400504
transform 1 0 1164 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_245
timestamp 1713400504
transform 1 0 1076 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_246
timestamp 1713400504
transform 1 0 996 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_247
timestamp 1713400504
transform 1 0 1100 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_248
timestamp 1713400504
transform 1 0 964 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_249
timestamp 1713400504
transform 1 0 780 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_250
timestamp 1713400504
transform 1 0 2228 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_251
timestamp 1713400504
transform 1 0 2036 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_252
timestamp 1713400504
transform 1 0 1956 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_253
timestamp 1713400504
transform 1 0 1948 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_254
timestamp 1713400504
transform 1 0 1860 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_255
timestamp 1713400504
transform 1 0 2196 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_256
timestamp 1713400504
transform 1 0 2092 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_257
timestamp 1713400504
transform 1 0 2324 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_258
timestamp 1713400504
transform 1 0 2268 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_259
timestamp 1713400504
transform 1 0 1092 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_260
timestamp 1713400504
transform 1 0 948 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_261
timestamp 1713400504
transform 1 0 1076 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_262
timestamp 1713400504
transform 1 0 1036 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_263
timestamp 1713400504
transform 1 0 2284 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_264
timestamp 1713400504
transform 1 0 2228 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_265
timestamp 1713400504
transform 1 0 2156 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_266
timestamp 1713400504
transform 1 0 2100 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_267
timestamp 1713400504
transform 1 0 1932 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_268
timestamp 1713400504
transform 1 0 1916 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_269
timestamp 1713400504
transform 1 0 1884 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_270
timestamp 1713400504
transform 1 0 1876 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_271
timestamp 1713400504
transform 1 0 2060 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_272
timestamp 1713400504
transform 1 0 2036 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_273
timestamp 1713400504
transform 1 0 2180 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_274
timestamp 1713400504
transform 1 0 2124 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_275
timestamp 1713400504
transform 1 0 1996 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_276
timestamp 1713400504
transform 1 0 1948 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_277
timestamp 1713400504
transform 1 0 1684 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_278
timestamp 1713400504
transform 1 0 1908 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_279
timestamp 1713400504
transform 1 0 1764 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_280
timestamp 1713400504
transform 1 0 1540 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_281
timestamp 1713400504
transform 1 0 1804 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_282
timestamp 1713400504
transform 1 0 1620 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_283
timestamp 1713400504
transform 1 0 2116 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_284
timestamp 1713400504
transform 1 0 1604 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_285
timestamp 1713400504
transform 1 0 1604 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_286
timestamp 1713400504
transform 1 0 1500 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_287
timestamp 1713400504
transform 1 0 1556 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_288
timestamp 1713400504
transform 1 0 1388 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_289
timestamp 1713400504
transform 1 0 1316 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_290
timestamp 1713400504
transform 1 0 1268 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_291
timestamp 1713400504
transform 1 0 1548 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_292
timestamp 1713400504
transform 1 0 1460 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_293
timestamp 1713400504
transform 1 0 1396 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_294
timestamp 1713400504
transform 1 0 1252 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_295
timestamp 1713400504
transform 1 0 1236 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_296
timestamp 1713400504
transform 1 0 1444 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_297
timestamp 1713400504
transform 1 0 1364 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_298
timestamp 1713400504
transform 1 0 2444 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_299
timestamp 1713400504
transform 1 0 1644 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_300
timestamp 1713400504
transform 1 0 1644 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_301
timestamp 1713400504
transform 1 0 1460 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_302
timestamp 1713400504
transform 1 0 1252 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_303
timestamp 1713400504
transform 1 0 1188 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_304
timestamp 1713400504
transform 1 0 2092 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_305
timestamp 1713400504
transform 1 0 1988 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_306
timestamp 1713400504
transform 1 0 1924 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_307
timestamp 1713400504
transform 1 0 1820 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_308
timestamp 1713400504
transform 1 0 2132 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_309
timestamp 1713400504
transform 1 0 2084 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_310
timestamp 1713400504
transform 1 0 2020 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_311
timestamp 1713400504
transform 1 0 2180 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_312
timestamp 1713400504
transform 1 0 2140 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_313
timestamp 1713400504
transform 1 0 2468 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_314
timestamp 1713400504
transform 1 0 2372 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_315
timestamp 1713400504
transform 1 0 2308 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_316
timestamp 1713400504
transform 1 0 2148 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_317
timestamp 1713400504
transform 1 0 2780 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_318
timestamp 1713400504
transform 1 0 2508 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_319
timestamp 1713400504
transform 1 0 2508 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_320
timestamp 1713400504
transform 1 0 2396 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_321
timestamp 1713400504
transform 1 0 2356 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_322
timestamp 1713400504
transform 1 0 2740 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_323
timestamp 1713400504
transform 1 0 2644 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_324
timestamp 1713400504
transform 1 0 2420 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_325
timestamp 1713400504
transform 1 0 2300 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_326
timestamp 1713400504
transform 1 0 2932 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_327
timestamp 1713400504
transform 1 0 2844 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_328
timestamp 1713400504
transform 1 0 2764 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_329
timestamp 1713400504
transform 1 0 2700 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_330
timestamp 1713400504
transform 1 0 2700 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_331
timestamp 1713400504
transform 1 0 2628 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_332
timestamp 1713400504
transform 1 0 2988 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_333
timestamp 1713400504
transform 1 0 2892 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_334
timestamp 1713400504
transform 1 0 2692 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_335
timestamp 1713400504
transform 1 0 2660 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_336
timestamp 1713400504
transform 1 0 2580 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_337
timestamp 1713400504
transform 1 0 2444 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_338
timestamp 1713400504
transform 1 0 2972 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_339
timestamp 1713400504
transform 1 0 2876 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_340
timestamp 1713400504
transform 1 0 2676 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_341
timestamp 1713400504
transform 1 0 2668 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_342
timestamp 1713400504
transform 1 0 2540 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_343
timestamp 1713400504
transform 1 0 2692 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_344
timestamp 1713400504
transform 1 0 2628 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_345
timestamp 1713400504
transform 1 0 2628 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_346
timestamp 1713400504
transform 1 0 2436 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_347
timestamp 1713400504
transform 1 0 2356 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_348
timestamp 1713400504
transform 1 0 2340 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_349
timestamp 1713400504
transform 1 0 2820 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_350
timestamp 1713400504
transform 1 0 2668 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_351
timestamp 1713400504
transform 1 0 2644 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_352
timestamp 1713400504
transform 1 0 2516 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_353
timestamp 1713400504
transform 1 0 2956 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_354
timestamp 1713400504
transform 1 0 2732 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_355
timestamp 1713400504
transform 1 0 2956 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_356
timestamp 1713400504
transform 1 0 2900 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_357
timestamp 1713400504
transform 1 0 2780 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_358
timestamp 1713400504
transform 1 0 2724 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_359
timestamp 1713400504
transform 1 0 2692 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_360
timestamp 1713400504
transform 1 0 2412 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_361
timestamp 1713400504
transform 1 0 2828 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_362
timestamp 1713400504
transform 1 0 2684 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_363
timestamp 1713400504
transform 1 0 2300 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_364
timestamp 1713400504
transform 1 0 2028 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_365
timestamp 1713400504
transform 1 0 1852 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_366
timestamp 1713400504
transform 1 0 1380 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_367
timestamp 1713400504
transform 1 0 1500 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_368
timestamp 1713400504
transform 1 0 1452 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_369
timestamp 1713400504
transform 1 0 2516 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_370
timestamp 1713400504
transform 1 0 2436 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_371
timestamp 1713400504
transform 1 0 2964 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_372
timestamp 1713400504
transform 1 0 2836 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_373
timestamp 1713400504
transform 1 0 2860 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_374
timestamp 1713400504
transform 1 0 2804 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_375
timestamp 1713400504
transform 1 0 2620 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_376
timestamp 1713400504
transform 1 0 2980 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_377
timestamp 1713400504
transform 1 0 2876 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_378
timestamp 1713400504
transform 1 0 2844 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_379
timestamp 1713400504
transform 1 0 2860 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_380
timestamp 1713400504
transform 1 0 2740 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_381
timestamp 1713400504
transform 1 0 2676 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_382
timestamp 1713400504
transform 1 0 2972 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_383
timestamp 1713400504
transform 1 0 2820 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_384
timestamp 1713400504
transform 1 0 2404 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_385
timestamp 1713400504
transform 1 0 2300 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_386
timestamp 1713400504
transform 1 0 2124 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_387
timestamp 1713400504
transform 1 0 2220 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_388
timestamp 1713400504
transform 1 0 2068 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_389
timestamp 1713400504
transform 1 0 2404 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_390
timestamp 1713400504
transform 1 0 2316 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_391
timestamp 1713400504
transform 1 0 2724 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_392
timestamp 1713400504
transform 1 0 2636 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_393
timestamp 1713400504
transform 1 0 2876 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_394
timestamp 1713400504
transform 1 0 2828 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_395
timestamp 1713400504
transform 1 0 2748 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_396
timestamp 1713400504
transform 1 0 2204 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_397
timestamp 1713400504
transform 1 0 2108 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_398
timestamp 1713400504
transform 1 0 2076 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_399
timestamp 1713400504
transform 1 0 1980 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_400
timestamp 1713400504
transform 1 0 2164 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_401
timestamp 1713400504
transform 1 0 2116 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_402
timestamp 1713400504
transform 1 0 2284 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_403
timestamp 1713400504
transform 1 0 2052 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_404
timestamp 1713400504
transform 1 0 1916 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_405
timestamp 1713400504
transform 1 0 1820 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_406
timestamp 1713400504
transform 1 0 1444 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_407
timestamp 1713400504
transform 1 0 724 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_408
timestamp 1713400504
transform 1 0 684 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_409
timestamp 1713400504
transform 1 0 564 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_410
timestamp 1713400504
transform 1 0 364 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_411
timestamp 1713400504
transform 1 0 284 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_412
timestamp 1713400504
transform 1 0 772 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_413
timestamp 1713400504
transform 1 0 716 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_414
timestamp 1713400504
transform 1 0 620 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_415
timestamp 1713400504
transform 1 0 620 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_416
timestamp 1713400504
transform 1 0 508 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_417
timestamp 1713400504
transform 1 0 356 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_418
timestamp 1713400504
transform 1 0 348 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_419
timestamp 1713400504
transform 1 0 340 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_420
timestamp 1713400504
transform 1 0 652 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_421
timestamp 1713400504
transform 1 0 604 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_422
timestamp 1713400504
transform 1 0 884 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_423
timestamp 1713400504
transform 1 0 828 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_424
timestamp 1713400504
transform 1 0 764 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_425
timestamp 1713400504
transform 1 0 612 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_426
timestamp 1713400504
transform 1 0 572 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_427
timestamp 1713400504
transform 1 0 508 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_428
timestamp 1713400504
transform 1 0 500 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_429
timestamp 1713400504
transform 1 0 292 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_430
timestamp 1713400504
transform 1 0 420 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_431
timestamp 1713400504
transform 1 0 364 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_432
timestamp 1713400504
transform 1 0 284 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_433
timestamp 1713400504
transform 1 0 420 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_434
timestamp 1713400504
transform 1 0 324 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_435
timestamp 1713400504
transform 1 0 212 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_436
timestamp 1713400504
transform 1 0 124 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_437
timestamp 1713400504
transform 1 0 100 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_438
timestamp 1713400504
transform 1 0 100 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_439
timestamp 1713400504
transform 1 0 212 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_440
timestamp 1713400504
transform 1 0 140 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_441
timestamp 1713400504
transform 1 0 92 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_442
timestamp 1713400504
transform 1 0 188 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_443
timestamp 1713400504
transform 1 0 124 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_444
timestamp 1713400504
transform 1 0 84 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_445
timestamp 1713400504
transform 1 0 196 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_446
timestamp 1713400504
transform 1 0 156 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_447
timestamp 1713400504
transform 1 0 84 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_448
timestamp 1713400504
transform 1 0 276 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_449
timestamp 1713400504
transform 1 0 220 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_450
timestamp 1713400504
transform 1 0 228 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_451
timestamp 1713400504
transform 1 0 148 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_452
timestamp 1713400504
transform 1 0 564 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_453
timestamp 1713400504
transform 1 0 468 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_454
timestamp 1713400504
transform 1 0 404 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_455
timestamp 1713400504
transform 1 0 372 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_456
timestamp 1713400504
transform 1 0 348 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_457
timestamp 1713400504
transform 1 0 324 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_458
timestamp 1713400504
transform 1 0 2492 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_459
timestamp 1713400504
transform 1 0 2132 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_460
timestamp 1713400504
transform 1 0 2116 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_461
timestamp 1713400504
transform 1 0 1924 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_462
timestamp 1713400504
transform 1 0 1868 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_463
timestamp 1713400504
transform 1 0 1780 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_464
timestamp 1713400504
transform 1 0 1780 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_465
timestamp 1713400504
transform 1 0 1556 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_466
timestamp 1713400504
transform 1 0 1348 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_467
timestamp 1713400504
transform 1 0 1300 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_468
timestamp 1713400504
transform 1 0 2892 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_469
timestamp 1713400504
transform 1 0 2716 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_470
timestamp 1713400504
transform 1 0 2540 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_471
timestamp 1713400504
transform 1 0 2732 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_472
timestamp 1713400504
transform 1 0 2684 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_473
timestamp 1713400504
transform 1 0 2772 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_474
timestamp 1713400504
transform 1 0 2732 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_475
timestamp 1713400504
transform 1 0 2948 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_476
timestamp 1713400504
transform 1 0 2900 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_477
timestamp 1713400504
transform 1 0 476 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_478
timestamp 1713400504
transform 1 0 396 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_479
timestamp 1713400504
transform 1 0 572 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_480
timestamp 1713400504
transform 1 0 484 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_481
timestamp 1713400504
transform 1 0 204 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_482
timestamp 1713400504
transform 1 0 148 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_483
timestamp 1713400504
transform 1 0 700 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_484
timestamp 1713400504
transform 1 0 620 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_485
timestamp 1713400504
transform 1 0 748 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_486
timestamp 1713400504
transform 1 0 684 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_487
timestamp 1713400504
transform 1 0 620 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_488
timestamp 1713400504
transform 1 0 548 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_489
timestamp 1713400504
transform 1 0 620 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_490
timestamp 1713400504
transform 1 0 516 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_491
timestamp 1713400504
transform 1 0 620 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_492
timestamp 1713400504
transform 1 0 532 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_493
timestamp 1713400504
transform 1 0 276 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_494
timestamp 1713400504
transform 1 0 204 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_495
timestamp 1713400504
transform 1 0 1084 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_496
timestamp 1713400504
transform 1 0 972 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_497
timestamp 1713400504
transform 1 0 284 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_498
timestamp 1713400504
transform 1 0 196 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_499
timestamp 1713400504
transform 1 0 204 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_500
timestamp 1713400504
transform 1 0 116 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_501
timestamp 1713400504
transform 1 0 180 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_502
timestamp 1713400504
transform 1 0 140 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_503
timestamp 1713400504
transform 1 0 924 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_504
timestamp 1713400504
transform 1 0 884 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_505
timestamp 1713400504
transform 1 0 1148 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_506
timestamp 1713400504
transform 1 0 1036 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_507
timestamp 1713400504
transform 1 0 1092 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_508
timestamp 1713400504
transform 1 0 996 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_509
timestamp 1713400504
transform 1 0 1028 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_510
timestamp 1713400504
transform 1 0 932 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_511
timestamp 1713400504
transform 1 0 644 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_512
timestamp 1713400504
transform 1 0 804 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_513
timestamp 1713400504
transform 1 0 740 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_514
timestamp 1713400504
transform 1 0 2932 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_515
timestamp 1713400504
transform 1 0 2860 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_516
timestamp 1713400504
transform 1 0 2772 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_517
timestamp 1713400504
transform 1 0 2676 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_518
timestamp 1713400504
transform 1 0 2636 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_519
timestamp 1713400504
transform 1 0 2540 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_520
timestamp 1713400504
transform 1 0 2532 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_521
timestamp 1713400504
transform 1 0 2500 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_522
timestamp 1713400504
transform 1 0 2484 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_523
timestamp 1713400504
transform 1 0 2436 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_524
timestamp 1713400504
transform 1 0 2956 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_525
timestamp 1713400504
transform 1 0 2932 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_526
timestamp 1713400504
transform 1 0 2924 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_527
timestamp 1713400504
transform 1 0 2924 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_528
timestamp 1713400504
transform 1 0 2924 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_529
timestamp 1713400504
transform 1 0 2868 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_530
timestamp 1713400504
transform 1 0 2852 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_531
timestamp 1713400504
transform 1 0 2852 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_532
timestamp 1713400504
transform 1 0 2820 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_533
timestamp 1713400504
transform 1 0 2764 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_534
timestamp 1713400504
transform 1 0 2684 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_535
timestamp 1713400504
transform 1 0 2620 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_536
timestamp 1713400504
transform 1 0 2572 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_537
timestamp 1713400504
transform 1 0 2604 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_538
timestamp 1713400504
transform 1 0 2508 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_539
timestamp 1713400504
transform 1 0 2212 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_540
timestamp 1713400504
transform 1 0 2052 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_541
timestamp 1713400504
transform 1 0 1852 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_542
timestamp 1713400504
transform 1 0 1836 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_543
timestamp 1713400504
transform 1 0 1668 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_544
timestamp 1713400504
transform 1 0 1660 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_545
timestamp 1713400504
transform 1 0 1620 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_546
timestamp 1713400504
transform 1 0 1596 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_547
timestamp 1713400504
transform 1 0 1300 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_548
timestamp 1713400504
transform 1 0 1172 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_549
timestamp 1713400504
transform 1 0 1076 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_550
timestamp 1713400504
transform 1 0 1068 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_551
timestamp 1713400504
transform 1 0 980 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_552
timestamp 1713400504
transform 1 0 2788 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_553
timestamp 1713400504
transform 1 0 2780 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_554
timestamp 1713400504
transform 1 0 2764 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_555
timestamp 1713400504
transform 1 0 2732 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_556
timestamp 1713400504
transform 1 0 2556 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_557
timestamp 1713400504
transform 1 0 2460 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_558
timestamp 1713400504
transform 1 0 2460 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_559
timestamp 1713400504
transform 1 0 2460 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_560
timestamp 1713400504
transform 1 0 2412 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_561
timestamp 1713400504
transform 1 0 2412 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_562
timestamp 1713400504
transform 1 0 2220 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_563
timestamp 1713400504
transform 1 0 2220 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_564
timestamp 1713400504
transform 1 0 2220 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_565
timestamp 1713400504
transform 1 0 2212 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_566
timestamp 1713400504
transform 1 0 2164 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_567
timestamp 1713400504
transform 1 0 2324 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_568
timestamp 1713400504
transform 1 0 2228 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_569
timestamp 1713400504
transform 1 0 2156 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_570
timestamp 1713400504
transform 1 0 2084 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_571
timestamp 1713400504
transform 1 0 2036 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_572
timestamp 1713400504
transform 1 0 2036 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_573
timestamp 1713400504
transform 1 0 1996 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_574
timestamp 1713400504
transform 1 0 1812 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_575
timestamp 1713400504
transform 1 0 1812 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_576
timestamp 1713400504
transform 1 0 1716 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_577
timestamp 1713400504
transform 1 0 1708 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_578
timestamp 1713400504
transform 1 0 1564 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_579
timestamp 1713400504
transform 1 0 1516 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_580
timestamp 1713400504
transform 1 0 1516 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_581
timestamp 1713400504
transform 1 0 1476 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_582
timestamp 1713400504
transform 1 0 1468 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_583
timestamp 1713400504
transform 1 0 1444 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_584
timestamp 1713400504
transform 1 0 1988 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_585
timestamp 1713400504
transform 1 0 1876 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_586
timestamp 1713400504
transform 1 0 1852 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_587
timestamp 1713400504
transform 1 0 1708 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_588
timestamp 1713400504
transform 1 0 1652 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_589
timestamp 1713400504
transform 1 0 1652 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_590
timestamp 1713400504
transform 1 0 1644 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_591
timestamp 1713400504
transform 1 0 1580 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_592
timestamp 1713400504
transform 1 0 1140 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_593
timestamp 1713400504
transform 1 0 1060 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_594
timestamp 1713400504
transform 1 0 1044 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_595
timestamp 1713400504
transform 1 0 1036 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_596
timestamp 1713400504
transform 1 0 836 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_597
timestamp 1713400504
transform 1 0 796 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_598
timestamp 1713400504
transform 1 0 740 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_599
timestamp 1713400504
transform 1 0 436 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_600
timestamp 1713400504
transform 1 0 964 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_601
timestamp 1713400504
transform 1 0 940 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_602
timestamp 1713400504
transform 1 0 940 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_603
timestamp 1713400504
transform 1 0 908 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_604
timestamp 1713400504
transform 1 0 892 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_605
timestamp 1713400504
transform 1 0 804 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_606
timestamp 1713400504
transform 1 0 716 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_607
timestamp 1713400504
transform 1 0 652 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_608
timestamp 1713400504
transform 1 0 612 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_609
timestamp 1713400504
transform 1 0 580 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_610
timestamp 1713400504
transform 1 0 508 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_611
timestamp 1713400504
transform 1 0 476 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_612
timestamp 1713400504
transform 1 0 396 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_613
timestamp 1713400504
transform 1 0 140 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_614
timestamp 1713400504
transform 1 0 92 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_615
timestamp 1713400504
transform 1 0 596 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_616
timestamp 1713400504
transform 1 0 596 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_617
timestamp 1713400504
transform 1 0 596 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_618
timestamp 1713400504
transform 1 0 468 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_619
timestamp 1713400504
transform 1 0 420 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_620
timestamp 1713400504
transform 1 0 388 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_621
timestamp 1713400504
transform 1 0 252 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_622
timestamp 1713400504
transform 1 0 236 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_623
timestamp 1713400504
transform 1 0 92 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_624
timestamp 1713400504
transform 1 0 84 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_625
timestamp 1713400504
transform 1 0 84 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_626
timestamp 1713400504
transform 1 0 756 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_627
timestamp 1713400504
transform 1 0 708 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_628
timestamp 1713400504
transform 1 0 2412 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_629
timestamp 1713400504
transform 1 0 2412 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_630
timestamp 1713400504
transform 1 0 2380 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_631
timestamp 1713400504
transform 1 0 2316 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_632
timestamp 1713400504
transform 1 0 2308 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_633
timestamp 1713400504
transform 1 0 2268 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_634
timestamp 1713400504
transform 1 0 2180 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_635
timestamp 1713400504
transform 1 0 2084 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_636
timestamp 1713400504
transform 1 0 2076 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_637
timestamp 1713400504
transform 1 0 2036 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_638
timestamp 1713400504
transform 1 0 2004 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_639
timestamp 1713400504
transform 1 0 1924 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_640
timestamp 1713400504
transform 1 0 2692 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_641
timestamp 1713400504
transform 1 0 2684 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_642
timestamp 1713400504
transform 1 0 2668 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_643
timestamp 1713400504
transform 1 0 2668 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_644
timestamp 1713400504
transform 1 0 2508 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_645
timestamp 1713400504
transform 1 0 2436 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_646
timestamp 1713400504
transform 1 0 2372 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_647
timestamp 1713400504
transform 1 0 2364 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_648
timestamp 1713400504
transform 1 0 2364 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_649
timestamp 1713400504
transform 1 0 2364 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_650
timestamp 1713400504
transform 1 0 2316 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_651
timestamp 1713400504
transform 1 0 2316 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_652
timestamp 1713400504
transform 1 0 2308 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_653
timestamp 1713400504
transform 1 0 2236 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_654
timestamp 1713400504
transform 1 0 2116 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_655
timestamp 1713400504
transform 1 0 2084 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_656
timestamp 1713400504
transform 1 0 2052 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_657
timestamp 1713400504
transform 1 0 2044 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_658
timestamp 1713400504
transform 1 0 2036 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_659
timestamp 1713400504
transform 1 0 1908 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_660
timestamp 1713400504
transform 1 0 1908 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_661
timestamp 1713400504
transform 1 0 1828 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_662
timestamp 1713400504
transform 1 0 1828 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_663
timestamp 1713400504
transform 1 0 1788 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_664
timestamp 1713400504
transform 1 0 1652 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_665
timestamp 1713400504
transform 1 0 1636 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_666
timestamp 1713400504
transform 1 0 2156 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_667
timestamp 1713400504
transform 1 0 2140 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_668
timestamp 1713400504
transform 1 0 1988 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_669
timestamp 1713400504
transform 1 0 1788 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_670
timestamp 1713400504
transform 1 0 1724 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_671
timestamp 1713400504
transform 1 0 1716 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_672
timestamp 1713400504
transform 1 0 1604 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_673
timestamp 1713400504
transform 1 0 1580 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_674
timestamp 1713400504
transform 1 0 1452 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_675
timestamp 1713400504
transform 1 0 1396 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_676
timestamp 1713400504
transform 1 0 1316 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_677
timestamp 1713400504
transform 1 0 1268 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_678
timestamp 1713400504
transform 1 0 1220 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_679
timestamp 1713400504
transform 1 0 1220 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_680
timestamp 1713400504
transform 1 0 2884 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_681
timestamp 1713400504
transform 1 0 2868 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_682
timestamp 1713400504
transform 1 0 2860 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_683
timestamp 1713400504
transform 1 0 2844 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_684
timestamp 1713400504
transform 1 0 2812 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_685
timestamp 1713400504
transform 1 0 2740 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_686
timestamp 1713400504
transform 1 0 2716 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_687
timestamp 1713400504
transform 1 0 2708 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_688
timestamp 1713400504
transform 1 0 2660 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_689
timestamp 1713400504
transform 1 0 2604 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_690
timestamp 1713400504
transform 1 0 2492 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_691
timestamp 1713400504
transform 1 0 2444 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_692
timestamp 1713400504
transform 1 0 2540 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_693
timestamp 1713400504
transform 1 0 2516 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_694
timestamp 1713400504
transform 1 0 2532 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_695
timestamp 1713400504
transform 1 0 2532 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_696
timestamp 1713400504
transform 1 0 2436 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_697
timestamp 1713400504
transform 1 0 2428 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_698
timestamp 1713400504
transform 1 0 2908 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_699
timestamp 1713400504
transform 1 0 2820 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_700
timestamp 1713400504
transform 1 0 2772 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_701
timestamp 1713400504
transform 1 0 2772 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_702
timestamp 1713400504
transform 1 0 2772 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_703
timestamp 1713400504
transform 1 0 2740 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_704
timestamp 1713400504
transform 1 0 2484 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_705
timestamp 1713400504
transform 1 0 2460 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_706
timestamp 1713400504
transform 1 0 2460 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_707
timestamp 1713400504
transform 1 0 2180 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_708
timestamp 1713400504
transform 1 0 2172 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_709
timestamp 1713400504
transform 1 0 2124 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_710
timestamp 1713400504
transform 1 0 2108 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_711
timestamp 1713400504
transform 1 0 2100 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_712
timestamp 1713400504
transform 1 0 2012 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_713
timestamp 1713400504
transform 1 0 1812 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_714
timestamp 1713400504
transform 1 0 1812 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_715
timestamp 1713400504
transform 1 0 1756 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_716
timestamp 1713400504
transform 1 0 1676 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_717
timestamp 1713400504
transform 1 0 1676 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_718
timestamp 1713400504
transform 1 0 1476 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_719
timestamp 1713400504
transform 1 0 1436 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_720
timestamp 1713400504
transform 1 0 1436 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_721
timestamp 1713400504
transform 1 0 1364 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_722
timestamp 1713400504
transform 1 0 1356 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_723
timestamp 1713400504
transform 1 0 1308 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_724
timestamp 1713400504
transform 1 0 1244 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_725
timestamp 1713400504
transform 1 0 1244 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_726
timestamp 1713400504
transform 1 0 1780 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_727
timestamp 1713400504
transform 1 0 1732 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_728
timestamp 1713400504
transform 1 0 1716 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_729
timestamp 1713400504
transform 1 0 1612 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_730
timestamp 1713400504
transform 1 0 1612 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_731
timestamp 1713400504
transform 1 0 1604 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_732
timestamp 1713400504
transform 1 0 1268 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_733
timestamp 1713400504
transform 1 0 1196 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_734
timestamp 1713400504
transform 1 0 1196 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_735
timestamp 1713400504
transform 1 0 1108 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_736
timestamp 1713400504
transform 1 0 1092 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_737
timestamp 1713400504
transform 1 0 1052 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_738
timestamp 1713400504
transform 1 0 980 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_739
timestamp 1713400504
transform 1 0 356 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_740
timestamp 1713400504
transform 1 0 324 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_741
timestamp 1713400504
transform 1 0 180 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_742
timestamp 1713400504
transform 1 0 980 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_743
timestamp 1713400504
transform 1 0 964 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_744
timestamp 1713400504
transform 1 0 908 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_745
timestamp 1713400504
transform 1 0 884 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_746
timestamp 1713400504
transform 1 0 884 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_747
timestamp 1713400504
transform 1 0 828 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_748
timestamp 1713400504
transform 1 0 812 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_749
timestamp 1713400504
transform 1 0 788 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_750
timestamp 1713400504
transform 1 0 700 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_751
timestamp 1713400504
transform 1 0 652 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_752
timestamp 1713400504
transform 1 0 580 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_753
timestamp 1713400504
transform 1 0 580 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_754
timestamp 1713400504
transform 1 0 540 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_755
timestamp 1713400504
transform 1 0 540 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_756
timestamp 1713400504
transform 1 0 532 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_757
timestamp 1713400504
transform 1 0 508 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_758
timestamp 1713400504
transform 1 0 500 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_759
timestamp 1713400504
transform 1 0 500 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_760
timestamp 1713400504
transform 1 0 500 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_761
timestamp 1713400504
transform 1 0 396 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_762
timestamp 1713400504
transform 1 0 332 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_763
timestamp 1713400504
transform 1 0 300 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_764
timestamp 1713400504
transform 1 0 268 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_765
timestamp 1713400504
transform 1 0 236 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_766
timestamp 1713400504
transform 1 0 236 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_767
timestamp 1713400504
transform 1 0 228 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_768
timestamp 1713400504
transform 1 0 180 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_769
timestamp 1713400504
transform 1 0 1988 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_770
timestamp 1713400504
transform 1 0 1964 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_771
timestamp 1713400504
transform 1 0 1924 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_772
timestamp 1713400504
transform 1 0 1916 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_773
timestamp 1713400504
transform 1 0 1916 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_774
timestamp 1713400504
transform 1 0 1892 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_775
timestamp 1713400504
transform 1 0 1860 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_776
timestamp 1713400504
transform 1 0 1828 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_777
timestamp 1713400504
transform 1 0 1828 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_778
timestamp 1713400504
transform 1 0 1820 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_779
timestamp 1713400504
transform 1 0 1788 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_780
timestamp 1713400504
transform 1 0 1780 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_781
timestamp 1713400504
transform 1 0 3004 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_782
timestamp 1713400504
transform 1 0 2948 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_783
timestamp 1713400504
transform 1 0 2644 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_784
timestamp 1713400504
transform 1 0 2596 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_785
timestamp 1713400504
transform 1 0 2396 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_786
timestamp 1713400504
transform 1 0 2084 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_787
timestamp 1713400504
transform 1 0 1980 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_788
timestamp 1713400504
transform 1 0 2540 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_789
timestamp 1713400504
transform 1 0 2460 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_790
timestamp 1713400504
transform 1 0 2444 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_791
timestamp 1713400504
transform 1 0 2356 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_792
timestamp 1713400504
transform 1 0 2324 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_793
timestamp 1713400504
transform 1 0 2324 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_794
timestamp 1713400504
transform 1 0 1988 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_795
timestamp 1713400504
transform 1 0 1940 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_796
timestamp 1713400504
transform 1 0 1716 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_797
timestamp 1713400504
transform 1 0 1564 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_798
timestamp 1713400504
transform 1 0 1564 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_799
timestamp 1713400504
transform 1 0 1476 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_800
timestamp 1713400504
transform 1 0 1508 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_801
timestamp 1713400504
transform 1 0 1468 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_802
timestamp 1713400504
transform 1 0 1444 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_803
timestamp 1713400504
transform 1 0 1684 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_804
timestamp 1713400504
transform 1 0 1596 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_805
timestamp 1713400504
transform 1 0 1420 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_806
timestamp 1713400504
transform 1 0 1332 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_807
timestamp 1713400504
transform 1 0 740 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_808
timestamp 1713400504
transform 1 0 684 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_809
timestamp 1713400504
transform 1 0 1380 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_810
timestamp 1713400504
transform 1 0 1324 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_811
timestamp 1713400504
transform 1 0 1332 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_812
timestamp 1713400504
transform 1 0 1268 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_813
timestamp 1713400504
transform 1 0 908 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_814
timestamp 1713400504
transform 1 0 852 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_815
timestamp 1713400504
transform 1 0 1340 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_816
timestamp 1713400504
transform 1 0 820 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_817
timestamp 1713400504
transform 1 0 788 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_818
timestamp 1713400504
transform 1 0 732 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_819
timestamp 1713400504
transform 1 0 732 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_820
timestamp 1713400504
transform 1 0 708 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_821
timestamp 1713400504
transform 1 0 652 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_822
timestamp 1713400504
transform 1 0 620 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_823
timestamp 1713400504
transform 1 0 596 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_824
timestamp 1713400504
transform 1 0 596 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_825
timestamp 1713400504
transform 1 0 540 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_826
timestamp 1713400504
transform 1 0 524 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_827
timestamp 1713400504
transform 1 0 484 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_828
timestamp 1713400504
transform 1 0 444 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_829
timestamp 1713400504
transform 1 0 444 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_830
timestamp 1713400504
transform 1 0 396 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_831
timestamp 1713400504
transform 1 0 380 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_832
timestamp 1713400504
transform 1 0 324 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_833
timestamp 1713400504
transform 1 0 252 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_834
timestamp 1713400504
transform 1 0 1500 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_835
timestamp 1713400504
transform 1 0 1444 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_836
timestamp 1713400504
transform 1 0 1324 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_837
timestamp 1713400504
transform 1 0 1268 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_838
timestamp 1713400504
transform 1 0 796 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_839
timestamp 1713400504
transform 1 0 724 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_840
timestamp 1713400504
transform 1 0 628 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_841
timestamp 1713400504
transform 1 0 548 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_842
timestamp 1713400504
transform 1 0 452 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_843
timestamp 1713400504
transform 1 0 380 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_844
timestamp 1713400504
transform 1 0 740 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_845
timestamp 1713400504
transform 1 0 708 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_846
timestamp 1713400504
transform 1 0 788 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_847
timestamp 1713400504
transform 1 0 684 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_848
timestamp 1713400504
transform 1 0 820 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_849
timestamp 1713400504
transform 1 0 700 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_850
timestamp 1713400504
transform 1 0 804 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_851
timestamp 1713400504
transform 1 0 540 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_852
timestamp 1713400504
transform 1 0 644 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_853
timestamp 1713400504
transform 1 0 532 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_854
timestamp 1713400504
transform 1 0 628 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_855
timestamp 1713400504
transform 1 0 524 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_856
timestamp 1713400504
transform 1 0 1028 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_857
timestamp 1713400504
transform 1 0 1020 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_858
timestamp 1713400504
transform 1 0 516 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_859
timestamp 1713400504
transform 1 0 420 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_860
timestamp 1713400504
transform 1 0 460 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_861
timestamp 1713400504
transform 1 0 388 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_862
timestamp 1713400504
transform 1 0 460 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_863
timestamp 1713400504
transform 1 0 388 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_864
timestamp 1713400504
transform 1 0 292 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_865
timestamp 1713400504
transform 1 0 252 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_866
timestamp 1713400504
transform 1 0 212 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_867
timestamp 1713400504
transform 1 0 148 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_868
timestamp 1713400504
transform 1 0 212 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_869
timestamp 1713400504
transform 1 0 148 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_870
timestamp 1713400504
transform 1 0 380 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_871
timestamp 1713400504
transform 1 0 292 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_872
timestamp 1713400504
transform 1 0 412 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_873
timestamp 1713400504
transform 1 0 316 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_874
timestamp 1713400504
transform 1 0 388 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_875
timestamp 1713400504
transform 1 0 324 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_876
timestamp 1713400504
transform 1 0 596 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_877
timestamp 1713400504
transform 1 0 508 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_878
timestamp 1713400504
transform 1 0 748 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_879
timestamp 1713400504
transform 1 0 644 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_880
timestamp 1713400504
transform 1 0 908 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_881
timestamp 1713400504
transform 1 0 812 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_882
timestamp 1713400504
transform 1 0 820 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_883
timestamp 1713400504
transform 1 0 724 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_884
timestamp 1713400504
transform 1 0 420 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_885
timestamp 1713400504
transform 1 0 356 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_886
timestamp 1713400504
transform 1 0 1556 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_887
timestamp 1713400504
transform 1 0 1428 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_888
timestamp 1713400504
transform 1 0 356 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_889
timestamp 1713400504
transform 1 0 324 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_890
timestamp 1713400504
transform 1 0 252 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_891
timestamp 1713400504
transform 1 0 332 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_892
timestamp 1713400504
transform 1 0 220 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_893
timestamp 1713400504
transform 1 0 420 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_894
timestamp 1713400504
transform 1 0 324 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_895
timestamp 1713400504
transform 1 0 540 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_896
timestamp 1713400504
transform 1 0 460 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_897
timestamp 1713400504
transform 1 0 708 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_898
timestamp 1713400504
transform 1 0 628 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_899
timestamp 1713400504
transform 1 0 628 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_900
timestamp 1713400504
transform 1 0 596 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_901
timestamp 1713400504
transform 1 0 732 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_902
timestamp 1713400504
transform 1 0 676 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_903
timestamp 1713400504
transform 1 0 852 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_904
timestamp 1713400504
transform 1 0 852 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_905
timestamp 1713400504
transform 1 0 820 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_906
timestamp 1713400504
transform 1 0 820 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_907
timestamp 1713400504
transform 1 0 932 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_908
timestamp 1713400504
transform 1 0 900 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_909
timestamp 1713400504
transform 1 0 844 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_910
timestamp 1713400504
transform 1 0 820 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_911
timestamp 1713400504
transform 1 0 820 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_912
timestamp 1713400504
transform 1 0 788 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_913
timestamp 1713400504
transform 1 0 756 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_914
timestamp 1713400504
transform 1 0 620 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_915
timestamp 1713400504
transform 1 0 524 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_916
timestamp 1713400504
transform 1 0 476 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_917
timestamp 1713400504
transform 1 0 316 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_918
timestamp 1713400504
transform 1 0 492 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_919
timestamp 1713400504
transform 1 0 228 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_920
timestamp 1713400504
transform 1 0 340 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_921
timestamp 1713400504
transform 1 0 284 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_922
timestamp 1713400504
transform 1 0 1684 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_923
timestamp 1713400504
transform 1 0 1276 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_924
timestamp 1713400504
transform 1 0 932 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_925
timestamp 1713400504
transform 1 0 1476 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_926
timestamp 1713400504
transform 1 0 1044 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_927
timestamp 1713400504
transform 1 0 932 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_928
timestamp 1713400504
transform 1 0 740 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_929
timestamp 1713400504
transform 1 0 732 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_930
timestamp 1713400504
transform 1 0 524 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_931
timestamp 1713400504
transform 1 0 492 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_932
timestamp 1713400504
transform 1 0 492 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_933
timestamp 1713400504
transform 1 0 364 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_934
timestamp 1713400504
transform 1 0 276 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_935
timestamp 1713400504
transform 1 0 212 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_936
timestamp 1713400504
transform 1 0 172 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_937
timestamp 1713400504
transform 1 0 172 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_938
timestamp 1713400504
transform 1 0 124 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_939
timestamp 1713400504
transform 1 0 284 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_940
timestamp 1713400504
transform 1 0 220 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_941
timestamp 1713400504
transform 1 0 492 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_942
timestamp 1713400504
transform 1 0 420 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_943
timestamp 1713400504
transform 1 0 380 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_944
timestamp 1713400504
transform 1 0 268 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_945
timestamp 1713400504
transform 1 0 244 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_946
timestamp 1713400504
transform 1 0 660 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_947
timestamp 1713400504
transform 1 0 556 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_948
timestamp 1713400504
transform 1 0 460 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_949
timestamp 1713400504
transform 1 0 436 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_950
timestamp 1713400504
transform 1 0 436 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_951
timestamp 1713400504
transform 1 0 300 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_952
timestamp 1713400504
transform 1 0 692 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_953
timestamp 1713400504
transform 1 0 676 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_954
timestamp 1713400504
transform 1 0 500 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_955
timestamp 1713400504
transform 1 0 452 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_956
timestamp 1713400504
transform 1 0 844 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_957
timestamp 1713400504
transform 1 0 820 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_958
timestamp 1713400504
transform 1 0 740 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_959
timestamp 1713400504
transform 1 0 620 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_960
timestamp 1713400504
transform 1 0 596 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_961
timestamp 1713400504
transform 1 0 460 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_962
timestamp 1713400504
transform 1 0 372 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_963
timestamp 1713400504
transform 1 0 340 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_964
timestamp 1713400504
transform 1 0 812 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_965
timestamp 1713400504
transform 1 0 684 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_966
timestamp 1713400504
transform 1 0 628 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_967
timestamp 1713400504
transform 1 0 540 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_968
timestamp 1713400504
transform 1 0 348 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_969
timestamp 1713400504
transform 1 0 516 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_970
timestamp 1713400504
transform 1 0 460 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_971
timestamp 1713400504
transform 1 0 268 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_972
timestamp 1713400504
transform 1 0 172 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_973
timestamp 1713400504
transform 1 0 156 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_974
timestamp 1713400504
transform 1 0 844 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_975
timestamp 1713400504
transform 1 0 772 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_976
timestamp 1713400504
transform 1 0 444 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_977
timestamp 1713400504
transform 1 0 388 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_978
timestamp 1713400504
transform 1 0 708 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_979
timestamp 1713400504
transform 1 0 468 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_980
timestamp 1713400504
transform 1 0 812 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_981
timestamp 1713400504
transform 1 0 764 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_982
timestamp 1713400504
transform 1 0 748 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_983
timestamp 1713400504
transform 1 0 612 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_984
timestamp 1713400504
transform 1 0 628 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_985
timestamp 1713400504
transform 1 0 572 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_986
timestamp 1713400504
transform 1 0 932 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_987
timestamp 1713400504
transform 1 0 804 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_988
timestamp 1713400504
transform 1 0 556 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_989
timestamp 1713400504
transform 1 0 220 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_990
timestamp 1713400504
transform 1 0 1164 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_991
timestamp 1713400504
transform 1 0 804 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_992
timestamp 1713400504
transform 1 0 732 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_993
timestamp 1713400504
transform 1 0 660 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_994
timestamp 1713400504
transform 1 0 676 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_995
timestamp 1713400504
transform 1 0 580 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_996
timestamp 1713400504
transform 1 0 580 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_997
timestamp 1713400504
transform 1 0 412 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_998
timestamp 1713400504
transform 1 0 324 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_999
timestamp 1713400504
transform 1 0 228 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1000
timestamp 1713400504
transform 1 0 348 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1001
timestamp 1713400504
transform 1 0 268 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1002
timestamp 1713400504
transform 1 0 444 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1003
timestamp 1713400504
transform 1 0 316 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1004
timestamp 1713400504
transform 1 0 356 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_1005
timestamp 1713400504
transform 1 0 228 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_1006
timestamp 1713400504
transform 1 0 348 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1007
timestamp 1713400504
transform 1 0 204 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1008
timestamp 1713400504
transform 1 0 652 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1009
timestamp 1713400504
transform 1 0 452 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1010
timestamp 1713400504
transform 1 0 292 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1011
timestamp 1713400504
transform 1 0 268 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1012
timestamp 1713400504
transform 1 0 332 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1013
timestamp 1713400504
transform 1 0 244 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1014
timestamp 1713400504
transform 1 0 276 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1015
timestamp 1713400504
transform 1 0 204 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1016
timestamp 1713400504
transform 1 0 244 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1017
timestamp 1713400504
transform 1 0 172 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1018
timestamp 1713400504
transform 1 0 92 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1019
timestamp 1713400504
transform 1 0 1508 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_1020
timestamp 1713400504
transform 1 0 1404 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_1021
timestamp 1713400504
transform 1 0 1324 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_1022
timestamp 1713400504
transform 1 0 884 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_1023
timestamp 1713400504
transform 1 0 380 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_1024
timestamp 1713400504
transform 1 0 420 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_1025
timestamp 1713400504
transform 1 0 356 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_1026
timestamp 1713400504
transform 1 0 372 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1027
timestamp 1713400504
transform 1 0 276 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1028
timestamp 1713400504
transform 1 0 1740 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1029
timestamp 1713400504
transform 1 0 1692 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1030
timestamp 1713400504
transform 1 0 716 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1031
timestamp 1713400504
transform 1 0 628 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1032
timestamp 1713400504
transform 1 0 844 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1033
timestamp 1713400504
transform 1 0 764 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1034
timestamp 1713400504
transform 1 0 556 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1035
timestamp 1713400504
transform 1 0 460 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1036
timestamp 1713400504
transform 1 0 964 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1037
timestamp 1713400504
transform 1 0 924 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1038
timestamp 1713400504
transform 1 0 1164 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_1039
timestamp 1713400504
transform 1 0 1060 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_1040
timestamp 1713400504
transform 1 0 836 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1041
timestamp 1713400504
transform 1 0 772 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1042
timestamp 1713400504
transform 1 0 548 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1043
timestamp 1713400504
transform 1 0 468 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1044
timestamp 1713400504
transform 1 0 220 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_1045
timestamp 1713400504
transform 1 0 140 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_1046
timestamp 1713400504
transform 1 0 220 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1047
timestamp 1713400504
transform 1 0 132 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1048
timestamp 1713400504
transform 1 0 1092 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1049
timestamp 1713400504
transform 1 0 1004 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1050
timestamp 1713400504
transform 1 0 868 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1051
timestamp 1713400504
transform 1 0 780 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1052
timestamp 1713400504
transform 1 0 196 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1053
timestamp 1713400504
transform 1 0 132 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1054
timestamp 1713400504
transform 1 0 620 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1055
timestamp 1713400504
transform 1 0 548 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1056
timestamp 1713400504
transform 1 0 412 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1057
timestamp 1713400504
transform 1 0 372 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1058
timestamp 1713400504
transform 1 0 460 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_1059
timestamp 1713400504
transform 1 0 380 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_1060
timestamp 1713400504
transform 1 0 1500 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_1061
timestamp 1713400504
transform 1 0 1420 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_1062
timestamp 1713400504
transform 1 0 2364 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1063
timestamp 1713400504
transform 1 0 2292 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1064
timestamp 1713400504
transform 1 0 2340 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1065
timestamp 1713400504
transform 1 0 2292 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1066
timestamp 1713400504
transform 1 0 1972 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1067
timestamp 1713400504
transform 1 0 1844 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1068
timestamp 1713400504
transform 1 0 1948 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1069
timestamp 1713400504
transform 1 0 1876 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1070
timestamp 1713400504
transform 1 0 1972 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1071
timestamp 1713400504
transform 1 0 1924 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1072
timestamp 1713400504
transform 1 0 1244 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1073
timestamp 1713400504
transform 1 0 1076 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1074
timestamp 1713400504
transform 1 0 1076 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1075
timestamp 1713400504
transform 1 0 996 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1076
timestamp 1713400504
transform 1 0 1300 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1077
timestamp 1713400504
transform 1 0 1236 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1078
timestamp 1713400504
transform 1 0 1188 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1079
timestamp 1713400504
transform 1 0 1076 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1080
timestamp 1713400504
transform 1 0 1236 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1081
timestamp 1713400504
transform 1 0 1108 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1082
timestamp 1713400504
transform 1 0 1060 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1083
timestamp 1713400504
transform 1 0 1204 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1084
timestamp 1713400504
transform 1 0 868 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1085
timestamp 1713400504
transform 1 0 756 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1086
timestamp 1713400504
transform 1 0 1356 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1087
timestamp 1713400504
transform 1 0 1300 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1088
timestamp 1713400504
transform 1 0 1556 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1089
timestamp 1713400504
transform 1 0 1420 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1090
timestamp 1713400504
transform 1 0 1244 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1091
timestamp 1713400504
transform 1 0 1156 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1092
timestamp 1713400504
transform 1 0 1156 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1093
timestamp 1713400504
transform 1 0 932 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1094
timestamp 1713400504
transform 1 0 884 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1095
timestamp 1713400504
transform 1 0 1308 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1096
timestamp 1713400504
transform 1 0 1196 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1097
timestamp 1713400504
transform 1 0 2204 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1098
timestamp 1713400504
transform 1 0 2100 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1099
timestamp 1713400504
transform 1 0 1964 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1100
timestamp 1713400504
transform 1 0 2204 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_1101
timestamp 1713400504
transform 1 0 1892 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_1102
timestamp 1713400504
transform 1 0 2172 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_1103
timestamp 1713400504
transform 1 0 1924 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_1104
timestamp 1713400504
transform 1 0 2364 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1105
timestamp 1713400504
transform 1 0 2260 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1106
timestamp 1713400504
transform 1 0 2444 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_1107
timestamp 1713400504
transform 1 0 2340 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_1108
timestamp 1713400504
transform 1 0 2380 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1109
timestamp 1713400504
transform 1 0 2324 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1110
timestamp 1713400504
transform 1 0 2876 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1111
timestamp 1713400504
transform 1 0 2740 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1112
timestamp 1713400504
transform 1 0 2980 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_1113
timestamp 1713400504
transform 1 0 2836 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_1114
timestamp 1713400504
transform 1 0 2876 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_1115
timestamp 1713400504
transform 1 0 2740 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_1116
timestamp 1713400504
transform 1 0 2884 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1117
timestamp 1713400504
transform 1 0 2756 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1118
timestamp 1713400504
transform 1 0 2828 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1119
timestamp 1713400504
transform 1 0 2692 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1120
timestamp 1713400504
transform 1 0 2996 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1121
timestamp 1713400504
transform 1 0 2868 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1122
timestamp 1713400504
transform 1 0 2980 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1123
timestamp 1713400504
transform 1 0 2868 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1124
timestamp 1713400504
transform 1 0 2244 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1125
timestamp 1713400504
transform 1 0 2012 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1126
timestamp 1713400504
transform 1 0 2228 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_1127
timestamp 1713400504
transform 1 0 2116 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_1128
timestamp 1713400504
transform 1 0 2404 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1129
timestamp 1713400504
transform 1 0 2116 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1130
timestamp 1713400504
transform 1 0 2236 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1131
timestamp 1713400504
transform 1 0 2052 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1132
timestamp 1713400504
transform 1 0 2292 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_1133
timestamp 1713400504
transform 1 0 2180 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_1134
timestamp 1713400504
transform 1 0 2284 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1135
timestamp 1713400504
transform 1 0 1932 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1136
timestamp 1713400504
transform 1 0 2180 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1137
timestamp 1713400504
transform 1 0 2084 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1138
timestamp 1713400504
transform 1 0 2452 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1139
timestamp 1713400504
transform 1 0 2300 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1140
timestamp 1713400504
transform 1 0 2972 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1141
timestamp 1713400504
transform 1 0 2948 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1142
timestamp 1713400504
transform 1 0 2868 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1143
timestamp 1713400504
transform 1 0 2812 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1144
timestamp 1713400504
transform 1 0 2740 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1145
timestamp 1713400504
transform 1 0 2684 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1146
timestamp 1713400504
transform 1 0 2676 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1147
timestamp 1713400504
transform 1 0 2660 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1148
timestamp 1713400504
transform 1 0 2580 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_1149
timestamp 1713400504
transform 1 0 2548 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_1150
timestamp 1713400504
transform 1 0 2540 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1151
timestamp 1713400504
transform 1 0 2500 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1152
timestamp 1713400504
transform 1 0 2500 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1153
timestamp 1713400504
transform 1 0 2468 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_1154
timestamp 1713400504
transform 1 0 2420 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_1155
timestamp 1713400504
transform 1 0 2420 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_1156
timestamp 1713400504
transform 1 0 2212 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_1157
timestamp 1713400504
transform 1 0 2204 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1158
timestamp 1713400504
transform 1 0 2076 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1159
timestamp 1713400504
transform 1 0 2540 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1160
timestamp 1713400504
transform 1 0 2452 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1161
timestamp 1713400504
transform 1 0 2604 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1162
timestamp 1713400504
transform 1 0 2508 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1163
timestamp 1713400504
transform 1 0 2636 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1164
timestamp 1713400504
transform 1 0 2460 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1165
timestamp 1713400504
transform 1 0 2396 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1166
timestamp 1713400504
transform 1 0 2348 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1167
timestamp 1713400504
transform 1 0 2444 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1168
timestamp 1713400504
transform 1 0 2356 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1169
timestamp 1713400504
transform 1 0 2508 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1170
timestamp 1713400504
transform 1 0 2332 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1171
timestamp 1713400504
transform 1 0 2428 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1172
timestamp 1713400504
transform 1 0 2340 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1173
timestamp 1713400504
transform 1 0 2452 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1174
timestamp 1713400504
transform 1 0 2316 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1175
timestamp 1713400504
transform 1 0 2428 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1176
timestamp 1713400504
transform 1 0 2284 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1177
timestamp 1713400504
transform 1 0 2340 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1178
timestamp 1713400504
transform 1 0 2132 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1179
timestamp 1713400504
transform 1 0 2300 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_1180
timestamp 1713400504
transform 1 0 2212 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_1181
timestamp 1713400504
transform 1 0 2684 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1182
timestamp 1713400504
transform 1 0 2348 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1183
timestamp 1713400504
transform 1 0 2364 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1184
timestamp 1713400504
transform 1 0 2020 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1185
timestamp 1713400504
transform 1 0 2148 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1186
timestamp 1713400504
transform 1 0 1516 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1187
timestamp 1713400504
transform 1 0 2796 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1188
timestamp 1713400504
transform 1 0 2748 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_1189
timestamp 1713400504
transform 1 0 2716 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1190
timestamp 1713400504
transform 1 0 2716 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_1191
timestamp 1713400504
transform 1 0 2884 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1192
timestamp 1713400504
transform 1 0 2820 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1193
timestamp 1713400504
transform 1 0 2772 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1194
timestamp 1713400504
transform 1 0 2724 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1195
timestamp 1713400504
transform 1 0 2884 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1196
timestamp 1713400504
transform 1 0 2748 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1197
timestamp 1713400504
transform 1 0 2852 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1198
timestamp 1713400504
transform 1 0 2788 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1199
timestamp 1713400504
transform 1 0 2884 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1200
timestamp 1713400504
transform 1 0 2764 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1201
timestamp 1713400504
transform 1 0 2876 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1202
timestamp 1713400504
transform 1 0 2788 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1203
timestamp 1713400504
transform 1 0 2620 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1204
timestamp 1713400504
transform 1 0 2588 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1205
timestamp 1713400504
transform 1 0 2492 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1206
timestamp 1713400504
transform 1 0 2388 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1207
timestamp 1713400504
transform 1 0 2620 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1208
timestamp 1713400504
transform 1 0 2572 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1209
timestamp 1713400504
transform 1 0 2540 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_1210
timestamp 1713400504
transform 1 0 2524 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_1211
timestamp 1713400504
transform 1 0 2564 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1212
timestamp 1713400504
transform 1 0 2516 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1213
timestamp 1713400504
transform 1 0 2484 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1214
timestamp 1713400504
transform 1 0 2420 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1215
timestamp 1713400504
transform 1 0 2492 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1216
timestamp 1713400504
transform 1 0 2436 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1217
timestamp 1713400504
transform 1 0 2324 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1218
timestamp 1713400504
transform 1 0 2324 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1219
timestamp 1713400504
transform 1 0 1860 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1220
timestamp 1713400504
transform 1 0 2732 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_1221
timestamp 1713400504
transform 1 0 2524 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_1222
timestamp 1713400504
transform 1 0 2516 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1223
timestamp 1713400504
transform 1 0 1996 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1224
timestamp 1713400504
transform 1 0 2556 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_1225
timestamp 1713400504
transform 1 0 2500 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_1226
timestamp 1713400504
transform 1 0 2492 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_1227
timestamp 1713400504
transform 1 0 1452 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_1228
timestamp 1713400504
transform 1 0 2524 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1229
timestamp 1713400504
transform 1 0 2476 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1230
timestamp 1713400504
transform 1 0 1652 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1231
timestamp 1713400504
transform 1 0 2268 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1232
timestamp 1713400504
transform 1 0 1540 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1233
timestamp 1713400504
transform 1 0 2268 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_1234
timestamp 1713400504
transform 1 0 1828 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1235
timestamp 1713400504
transform 1 0 2604 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1236
timestamp 1713400504
transform 1 0 2308 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1237
timestamp 1713400504
transform 1 0 2748 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1238
timestamp 1713400504
transform 1 0 2612 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1239
timestamp 1713400504
transform 1 0 2572 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1240
timestamp 1713400504
transform 1 0 2468 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1241
timestamp 1713400504
transform 1 0 1836 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1242
timestamp 1713400504
transform 1 0 1740 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1243
timestamp 1713400504
transform 1 0 2668 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1244
timestamp 1713400504
transform 1 0 2620 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1245
timestamp 1713400504
transform 1 0 2740 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1246
timestamp 1713400504
transform 1 0 2724 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1247
timestamp 1713400504
transform 1 0 2492 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1248
timestamp 1713400504
transform 1 0 2396 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1249
timestamp 1713400504
transform 1 0 1628 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1250
timestamp 1713400504
transform 1 0 1372 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1251
timestamp 1713400504
transform 1 0 2588 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1252
timestamp 1713400504
transform 1 0 2500 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1253
timestamp 1713400504
transform 1 0 2908 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1254
timestamp 1713400504
transform 1 0 2764 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1255
timestamp 1713400504
transform 1 0 2844 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_1256
timestamp 1713400504
transform 1 0 2652 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_1257
timestamp 1713400504
transform 1 0 1996 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_1258
timestamp 1713400504
transform 1 0 1940 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_1259
timestamp 1713400504
transform 1 0 2812 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_1260
timestamp 1713400504
transform 1 0 2628 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_1261
timestamp 1713400504
transform 1 0 2676 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1262
timestamp 1713400504
transform 1 0 2548 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1263
timestamp 1713400504
transform 1 0 2660 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_1264
timestamp 1713400504
transform 1 0 2572 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_1265
timestamp 1713400504
transform 1 0 2580 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1266
timestamp 1713400504
transform 1 0 2500 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1267
timestamp 1713400504
transform 1 0 2636 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1268
timestamp 1713400504
transform 1 0 2540 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1269
timestamp 1713400504
transform 1 0 2700 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1270
timestamp 1713400504
transform 1 0 2620 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1271
timestamp 1713400504
transform 1 0 2892 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1272
timestamp 1713400504
transform 1 0 2812 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1273
timestamp 1713400504
transform 1 0 1764 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_1274
timestamp 1713400504
transform 1 0 1396 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_1275
timestamp 1713400504
transform 1 0 1852 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_1276
timestamp 1713400504
transform 1 0 1740 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_1277
timestamp 1713400504
transform 1 0 1700 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1278
timestamp 1713400504
transform 1 0 1652 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1279
timestamp 1713400504
transform 1 0 1628 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1280
timestamp 1713400504
transform 1 0 1596 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1281
timestamp 1713400504
transform 1 0 1692 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1282
timestamp 1713400504
transform 1 0 1364 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1283
timestamp 1713400504
transform 1 0 1372 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1284
timestamp 1713400504
transform 1 0 1108 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1285
timestamp 1713400504
transform 1 0 1324 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_1286
timestamp 1713400504
transform 1 0 1244 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_1287
timestamp 1713400504
transform 1 0 1284 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1288
timestamp 1713400504
transform 1 0 1268 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1289
timestamp 1713400504
transform 1 0 1292 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_1290
timestamp 1713400504
transform 1 0 1260 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_1291
timestamp 1713400504
transform 1 0 1852 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1292
timestamp 1713400504
transform 1 0 1676 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1293
timestamp 1713400504
transform 1 0 1556 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1294
timestamp 1713400504
transform 1 0 1484 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1295
timestamp 1713400504
transform 1 0 1484 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1296
timestamp 1713400504
transform 1 0 1452 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1297
timestamp 1713400504
transform 1 0 2556 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1298
timestamp 1713400504
transform 1 0 2380 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1299
timestamp 1713400504
transform 1 0 2380 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1300
timestamp 1713400504
transform 1 0 1540 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1301
timestamp 1713400504
transform 1 0 2684 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1302
timestamp 1713400504
transform 1 0 2572 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1303
timestamp 1713400504
transform 1 0 1508 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1304
timestamp 1713400504
transform 1 0 1452 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1305
timestamp 1713400504
transform 1 0 1636 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1306
timestamp 1713400504
transform 1 0 1524 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1307
timestamp 1713400504
transform 1 0 1476 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1308
timestamp 1713400504
transform 1 0 1444 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1309
timestamp 1713400504
transform 1 0 1836 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1310
timestamp 1713400504
transform 1 0 1508 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1311
timestamp 1713400504
transform 1 0 2444 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1312
timestamp 1713400504
transform 1 0 2084 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1313
timestamp 1713400504
transform 1 0 2180 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1314
timestamp 1713400504
transform 1 0 2172 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_1315
timestamp 1713400504
transform 1 0 2124 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1316
timestamp 1713400504
transform 1 0 2116 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1317
timestamp 1713400504
transform 1 0 2116 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_1318
timestamp 1713400504
transform 1 0 2100 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1319
timestamp 1713400504
transform 1 0 2084 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1320
timestamp 1713400504
transform 1 0 2188 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1321
timestamp 1713400504
transform 1 0 2188 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_1322
timestamp 1713400504
transform 1 0 2172 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1323
timestamp 1713400504
transform 1 0 2116 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1324
timestamp 1713400504
transform 1 0 2108 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1325
timestamp 1713400504
transform 1 0 2084 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_1326
timestamp 1713400504
transform 1 0 2740 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1327
timestamp 1713400504
transform 1 0 2428 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1328
timestamp 1713400504
transform 1 0 2756 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1329
timestamp 1713400504
transform 1 0 2420 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1330
timestamp 1713400504
transform 1 0 2540 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1331
timestamp 1713400504
transform 1 0 2396 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1332
timestamp 1713400504
transform 1 0 2716 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1333
timestamp 1713400504
transform 1 0 2428 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1334
timestamp 1713400504
transform 1 0 2684 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1335
timestamp 1713400504
transform 1 0 2412 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1336
timestamp 1713400504
transform 1 0 2724 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1337
timestamp 1713400504
transform 1 0 2420 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1338
timestamp 1713400504
transform 1 0 1852 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1339
timestamp 1713400504
transform 1 0 1668 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1340
timestamp 1713400504
transform 1 0 1860 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_1341
timestamp 1713400504
transform 1 0 1572 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_1342
timestamp 1713400504
transform 1 0 1900 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_1343
timestamp 1713400504
transform 1 0 1620 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_1344
timestamp 1713400504
transform 1 0 1812 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1345
timestamp 1713400504
transform 1 0 1604 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1346
timestamp 1713400504
transform 1 0 1868 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1347
timestamp 1713400504
transform 1 0 1660 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1348
timestamp 1713400504
transform 1 0 2132 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1349
timestamp 1713400504
transform 1 0 2076 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1350
timestamp 1713400504
transform 1 0 1940 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1351
timestamp 1713400504
transform 1 0 1852 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1352
timestamp 1713400504
transform 1 0 2316 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_1353
timestamp 1713400504
transform 1 0 2212 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1354
timestamp 1713400504
transform 1 0 2108 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_1355
timestamp 1713400504
transform 1 0 2028 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1356
timestamp 1713400504
transform 1 0 1988 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1357
timestamp 1713400504
transform 1 0 2052 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1358
timestamp 1713400504
transform 1 0 1948 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1359
timestamp 1713400504
transform 1 0 1868 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1360
timestamp 1713400504
transform 1 0 1404 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1361
timestamp 1713400504
transform 1 0 2908 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_1362
timestamp 1713400504
transform 1 0 2908 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1363
timestamp 1713400504
transform 1 0 2164 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1364
timestamp 1713400504
transform 1 0 2060 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1365
timestamp 1713400504
transform 1 0 2020 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1366
timestamp 1713400504
transform 1 0 1388 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1367
timestamp 1713400504
transform 1 0 2132 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1368
timestamp 1713400504
transform 1 0 2044 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_1369
timestamp 1713400504
transform 1 0 2044 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1370
timestamp 1713400504
transform 1 0 2020 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1371
timestamp 1713400504
transform 1 0 1956 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1372
timestamp 1713400504
transform 1 0 1948 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_1373
timestamp 1713400504
transform 1 0 1524 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1374
timestamp 1713400504
transform 1 0 2060 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1375
timestamp 1713400504
transform 1 0 2004 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1376
timestamp 1713400504
transform 1 0 1964 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1377
timestamp 1713400504
transform 1 0 1940 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1378
timestamp 1713400504
transform 1 0 1612 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1379
timestamp 1713400504
transform 1 0 2124 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1380
timestamp 1713400504
transform 1 0 2028 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1381
timestamp 1713400504
transform 1 0 2324 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1382
timestamp 1713400504
transform 1 0 2284 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1383
timestamp 1713400504
transform 1 0 2260 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1384
timestamp 1713400504
transform 1 0 2220 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1385
timestamp 1713400504
transform 1 0 2340 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1386
timestamp 1713400504
transform 1 0 2164 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_1387
timestamp 1713400504
transform 1 0 2196 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1388
timestamp 1713400504
transform 1 0 2148 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1389
timestamp 1713400504
transform 1 0 2100 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1390
timestamp 1713400504
transform 1 0 1980 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1391
timestamp 1713400504
transform 1 0 1916 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1392
timestamp 1713400504
transform 1 0 1836 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1393
timestamp 1713400504
transform 1 0 1636 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1394
timestamp 1713400504
transform 1 0 1636 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1395
timestamp 1713400504
transform 1 0 1572 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1396
timestamp 1713400504
transform 1 0 1716 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1397
timestamp 1713400504
transform 1 0 1612 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1398
timestamp 1713400504
transform 1 0 1628 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1399
timestamp 1713400504
transform 1 0 1588 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1400
timestamp 1713400504
transform 1 0 1804 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1401
timestamp 1713400504
transform 1 0 1740 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1402
timestamp 1713400504
transform 1 0 1708 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1403
timestamp 1713400504
transform 1 0 1820 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1404
timestamp 1713400504
transform 1 0 1724 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1405
timestamp 1713400504
transform 1 0 1852 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1406
timestamp 1713400504
transform 1 0 1724 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1407
timestamp 1713400504
transform 1 0 1908 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_1408
timestamp 1713400504
transform 1 0 1724 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_1409
timestamp 1713400504
transform 1 0 1716 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_1410
timestamp 1713400504
transform 1 0 1556 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_1411
timestamp 1713400504
transform 1 0 1724 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_1412
timestamp 1713400504
transform 1 0 1500 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_1413
timestamp 1713400504
transform 1 0 1812 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1414
timestamp 1713400504
transform 1 0 1724 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1415
timestamp 1713400504
transform 1 0 1684 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1416
timestamp 1713400504
transform 1 0 1604 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1417
timestamp 1713400504
transform 1 0 1804 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1418
timestamp 1713400504
transform 1 0 1772 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1419
timestamp 1713400504
transform 1 0 1812 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1420
timestamp 1713400504
transform 1 0 1716 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1421
timestamp 1713400504
transform 1 0 1804 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1422
timestamp 1713400504
transform 1 0 1620 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1423
timestamp 1713400504
transform 1 0 1508 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1424
timestamp 1713400504
transform 1 0 1700 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1425
timestamp 1713400504
transform 1 0 1612 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1426
timestamp 1713400504
transform 1 0 1692 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1427
timestamp 1713400504
transform 1 0 1588 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1428
timestamp 1713400504
transform 1 0 1716 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1429
timestamp 1713400504
transform 1 0 1468 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1430
timestamp 1713400504
transform 1 0 1716 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1431
timestamp 1713400504
transform 1 0 1620 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1432
timestamp 1713400504
transform 1 0 1708 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1433
timestamp 1713400504
transform 1 0 1580 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1434
timestamp 1713400504
transform 1 0 1620 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_1435
timestamp 1713400504
transform 1 0 1524 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_1436
timestamp 1713400504
transform 1 0 1676 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1437
timestamp 1713400504
transform 1 0 1532 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1438
timestamp 1713400504
transform 1 0 1468 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1439
timestamp 1713400504
transform 1 0 1636 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1440
timestamp 1713400504
transform 1 0 1572 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1441
timestamp 1713400504
transform 1 0 1436 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1442
timestamp 1713400504
transform 1 0 1580 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1443
timestamp 1713400504
transform 1 0 1404 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1444
timestamp 1713400504
transform 1 0 1308 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1445
timestamp 1713400504
transform 1 0 1508 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_1446
timestamp 1713400504
transform 1 0 1420 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_1447
timestamp 1713400504
transform 1 0 1484 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_1448
timestamp 1713400504
transform 1 0 1420 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_1449
timestamp 1713400504
transform 1 0 1436 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1450
timestamp 1713400504
transform 1 0 1324 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1451
timestamp 1713400504
transform 1 0 1676 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_1452
timestamp 1713400504
transform 1 0 1628 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_1453
timestamp 1713400504
transform 1 0 1692 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_1454
timestamp 1713400504
transform 1 0 1588 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_1455
timestamp 1713400504
transform 1 0 1580 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1456
timestamp 1713400504
transform 1 0 1476 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1457
timestamp 1713400504
transform 1 0 1532 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1458
timestamp 1713400504
transform 1 0 1484 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1459
timestamp 1713400504
transform 1 0 1588 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1460
timestamp 1713400504
transform 1 0 1468 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1461
timestamp 1713400504
transform 1 0 1356 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1462
timestamp 1713400504
transform 1 0 1324 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1463
timestamp 1713400504
transform 1 0 1148 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1464
timestamp 1713400504
transform 1 0 884 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1465
timestamp 1713400504
transform 1 0 996 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1466
timestamp 1713400504
transform 1 0 860 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1467
timestamp 1713400504
transform 1 0 1044 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_1468
timestamp 1713400504
transform 1 0 1036 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1469
timestamp 1713400504
transform 1 0 964 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1470
timestamp 1713400504
transform 1 0 964 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_1471
timestamp 1713400504
transform 1 0 1148 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1472
timestamp 1713400504
transform 1 0 1116 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1473
timestamp 1713400504
transform 1 0 1084 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1474
timestamp 1713400504
transform 1 0 1020 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1475
timestamp 1713400504
transform 1 0 980 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1476
timestamp 1713400504
transform 1 0 980 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1477
timestamp 1713400504
transform 1 0 1004 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1478
timestamp 1713400504
transform 1 0 964 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1479
timestamp 1713400504
transform 1 0 924 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1480
timestamp 1713400504
transform 1 0 924 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1481
timestamp 1713400504
transform 1 0 772 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1482
timestamp 1713400504
transform 1 0 724 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1483
timestamp 1713400504
transform 1 0 1036 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_1484
timestamp 1713400504
transform 1 0 972 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1485
timestamp 1713400504
transform 1 0 900 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_1486
timestamp 1713400504
transform 1 0 900 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1487
timestamp 1713400504
transform 1 0 876 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_1488
timestamp 1713400504
transform 1 0 868 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1489
timestamp 1713400504
transform 1 0 756 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1490
timestamp 1713400504
transform 1 0 868 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1491
timestamp 1713400504
transform 1 0 748 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1492
timestamp 1713400504
transform 1 0 972 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1493
timestamp 1713400504
transform 1 0 876 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1494
timestamp 1713400504
transform 1 0 1124 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1495
timestamp 1713400504
transform 1 0 1028 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1496
timestamp 1713400504
transform 1 0 1268 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1497
timestamp 1713400504
transform 1 0 868 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1498
timestamp 1713400504
transform 1 0 972 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1499
timestamp 1713400504
transform 1 0 868 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1500
timestamp 1713400504
transform 1 0 764 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1501
timestamp 1713400504
transform 1 0 740 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1502
timestamp 1713400504
transform 1 0 948 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1503
timestamp 1713400504
transform 1 0 844 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1504
timestamp 1713400504
transform 1 0 1620 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1505
timestamp 1713400504
transform 1 0 1564 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1506
timestamp 1713400504
transform 1 0 1468 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1507
timestamp 1713400504
transform 1 0 1420 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1508
timestamp 1713400504
transform 1 0 1292 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1509
timestamp 1713400504
transform 1 0 1252 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1510
timestamp 1713400504
transform 1 0 1188 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1511
timestamp 1713400504
transform 1 0 1188 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1512
timestamp 1713400504
transform 1 0 1116 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1513
timestamp 1713400504
transform 1 0 1356 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1514
timestamp 1713400504
transform 1 0 1284 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1515
timestamp 1713400504
transform 1 0 1404 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1516
timestamp 1713400504
transform 1 0 1292 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1517
timestamp 1713400504
transform 1 0 1268 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1518
timestamp 1713400504
transform 1 0 1220 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1519
timestamp 1713400504
transform 1 0 1188 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1520
timestamp 1713400504
transform 1 0 1252 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1521
timestamp 1713400504
transform 1 0 1204 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1522
timestamp 1713400504
transform 1 0 1324 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1523
timestamp 1713400504
transform 1 0 1260 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1524
timestamp 1713400504
transform 1 0 1324 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1525
timestamp 1713400504
transform 1 0 1204 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1526
timestamp 1713400504
transform 1 0 1540 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1527
timestamp 1713400504
transform 1 0 1436 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1528
timestamp 1713400504
transform 1 0 1388 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1529
timestamp 1713400504
transform 1 0 1180 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1530
timestamp 1713400504
transform 1 0 1460 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1531
timestamp 1713400504
transform 1 0 1276 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1532
timestamp 1713400504
transform 1 0 1300 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1533
timestamp 1713400504
transform 1 0 1236 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1534
timestamp 1713400504
transform 1 0 1156 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1535
timestamp 1713400504
transform 1 0 932 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1536
timestamp 1713400504
transform 1 0 1076 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1537
timestamp 1713400504
transform 1 0 1036 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1538
timestamp 1713400504
transform 1 0 860 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1539
timestamp 1713400504
transform 1 0 724 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1540
timestamp 1713400504
transform 1 0 1052 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1541
timestamp 1713400504
transform 1 0 948 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1542
timestamp 1713400504
transform 1 0 1020 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1543
timestamp 1713400504
transform 1 0 836 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1544
timestamp 1713400504
transform 1 0 1148 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1545
timestamp 1713400504
transform 1 0 1092 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1546
timestamp 1713400504
transform 1 0 1092 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1547
timestamp 1713400504
transform 1 0 852 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1548
timestamp 1713400504
transform 1 0 988 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1549
timestamp 1713400504
transform 1 0 948 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1550
timestamp 1713400504
transform 1 0 724 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1551
timestamp 1713400504
transform 1 0 964 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1552
timestamp 1713400504
transform 1 0 740 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1553
timestamp 1713400504
transform 1 0 724 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1554
timestamp 1713400504
transform 1 0 660 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1555
timestamp 1713400504
transform 1 0 556 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1556
timestamp 1713400504
transform 1 0 820 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1557
timestamp 1713400504
transform 1 0 732 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1558
timestamp 1713400504
transform 1 0 1156 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1559
timestamp 1713400504
transform 1 0 1092 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1560
timestamp 1713400504
transform 1 0 1132 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1561
timestamp 1713400504
transform 1 0 1028 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1562
timestamp 1713400504
transform 1 0 1124 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1563
timestamp 1713400504
transform 1 0 964 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1564
timestamp 1713400504
transform 1 0 1132 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1565
timestamp 1713400504
transform 1 0 1084 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1566
timestamp 1713400504
transform 1 0 1244 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1567
timestamp 1713400504
transform 1 0 828 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_1568
timestamp 1713400504
transform 1 0 676 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1569
timestamp 1713400504
transform 1 0 548 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1570
timestamp 1713400504
transform 1 0 844 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1571
timestamp 1713400504
transform 1 0 740 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1572
timestamp 1713400504
transform 1 0 844 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1573
timestamp 1713400504
transform 1 0 652 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1574
timestamp 1713400504
transform 1 0 1380 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1575
timestamp 1713400504
transform 1 0 1228 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1576
timestamp 1713400504
transform 1 0 1268 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1577
timestamp 1713400504
transform 1 0 1148 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1578
timestamp 1713400504
transform 1 0 1252 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1579
timestamp 1713400504
transform 1 0 1092 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1580
timestamp 1713400504
transform 1 0 1100 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_1581
timestamp 1713400504
transform 1 0 1044 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_1582
timestamp 1713400504
transform 1 0 1044 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1583
timestamp 1713400504
transform 1 0 764 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1584
timestamp 1713400504
transform 1 0 1100 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1585
timestamp 1713400504
transform 1 0 1020 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_1586
timestamp 1713400504
transform 1 0 940 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1587
timestamp 1713400504
transform 1 0 900 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_1588
timestamp 1713400504
transform 1 0 844 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_1589
timestamp 1713400504
transform 1 0 1292 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1590
timestamp 1713400504
transform 1 0 1292 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1591
timestamp 1713400504
transform 1 0 1108 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1592
timestamp 1713400504
transform 1 0 996 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1593
timestamp 1713400504
transform 1 0 956 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1594
timestamp 1713400504
transform 1 0 884 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1595
timestamp 1713400504
transform 1 0 884 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1596
timestamp 1713400504
transform 1 0 884 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1597
timestamp 1713400504
transform 1 0 1148 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1598
timestamp 1713400504
transform 1 0 972 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1599
timestamp 1713400504
transform 1 0 796 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1600
timestamp 1713400504
transform 1 0 772 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1601
timestamp 1713400504
transform 1 0 756 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1602
timestamp 1713400504
transform 1 0 1156 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1603
timestamp 1713400504
transform 1 0 1100 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1604
timestamp 1713400504
transform 1 0 1012 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1605
timestamp 1713400504
transform 1 0 876 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_1606
timestamp 1713400504
transform 1 0 812 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1607
timestamp 1713400504
transform 1 0 780 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1608
timestamp 1713400504
transform 1 0 772 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_1609
timestamp 1713400504
transform 1 0 900 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1610
timestamp 1713400504
transform 1 0 772 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1611
timestamp 1713400504
transform 1 0 1180 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1612
timestamp 1713400504
transform 1 0 1132 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1613
timestamp 1713400504
transform 1 0 1172 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_1614
timestamp 1713400504
transform 1 0 964 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_1615
timestamp 1713400504
transform 1 0 2556 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_1616
timestamp 1713400504
transform 1 0 2508 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_1617
timestamp 1713400504
transform 1 0 2564 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1618
timestamp 1713400504
transform 1 0 2524 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1619
timestamp 1713400504
transform 1 0 2524 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1620
timestamp 1713400504
transform 1 0 2452 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1621
timestamp 1713400504
transform 1 0 2596 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1622
timestamp 1713400504
transform 1 0 2540 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1623
timestamp 1713400504
transform 1 0 2196 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1624
timestamp 1713400504
transform 1 0 2100 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1625
timestamp 1713400504
transform 1 0 2244 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1626
timestamp 1713400504
transform 1 0 2164 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1627
timestamp 1713400504
transform 1 0 1468 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1628
timestamp 1713400504
transform 1 0 1420 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1629
timestamp 1713400504
transform 1 0 1740 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1630
timestamp 1713400504
transform 1 0 1644 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1631
timestamp 1713400504
transform 1 0 1428 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1632
timestamp 1713400504
transform 1 0 1348 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_1633
timestamp 1713400504
transform 1 0 1292 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_1634
timestamp 1713400504
transform 1 0 1220 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_1635
timestamp 1713400504
transform 1 0 1236 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_1636
timestamp 1713400504
transform 1 0 1108 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_1637
timestamp 1713400504
transform 1 0 1348 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_1638
timestamp 1713400504
transform 1 0 1028 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_1639
timestamp 1713400504
transform 1 0 1236 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_1640
timestamp 1713400504
transform 1 0 1124 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_1641
timestamp 1713400504
transform 1 0 1804 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_1642
timestamp 1713400504
transform 1 0 1708 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_1643
timestamp 1713400504
transform 1 0 2004 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_1644
timestamp 1713400504
transform 1 0 1900 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_1645
timestamp 1713400504
transform 1 0 2172 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1646
timestamp 1713400504
transform 1 0 2100 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1647
timestamp 1713400504
transform 1 0 2532 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_1648
timestamp 1713400504
transform 1 0 2452 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_1649
timestamp 1713400504
transform 1 0 2764 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_1650
timestamp 1713400504
transform 1 0 2652 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_1651
timestamp 1713400504
transform 1 0 2844 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1652
timestamp 1713400504
transform 1 0 2724 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1653
timestamp 1713400504
transform 1 0 2956 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1654
timestamp 1713400504
transform 1 0 2860 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1655
timestamp 1713400504
transform 1 0 2796 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1656
timestamp 1713400504
transform 1 0 2676 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1657
timestamp 1713400504
transform 1 0 2948 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1658
timestamp 1713400504
transform 1 0 2804 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1659
timestamp 1713400504
transform 1 0 2900 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_1660
timestamp 1713400504
transform 1 0 2812 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_1661
timestamp 1713400504
transform 1 0 2804 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1662
timestamp 1713400504
transform 1 0 2740 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1663
timestamp 1713400504
transform 1 0 2756 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1664
timestamp 1713400504
transform 1 0 2716 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1665
timestamp 1713400504
transform 1 0 2332 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1666
timestamp 1713400504
transform 1 0 2236 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1667
timestamp 1713400504
transform 1 0 2132 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1668
timestamp 1713400504
transform 1 0 2044 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1669
timestamp 1713400504
transform 1 0 1668 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_1670
timestamp 1713400504
transform 1 0 1596 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_1671
timestamp 1713400504
transform 1 0 1596 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1672
timestamp 1713400504
transform 1 0 1516 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1673
timestamp 1713400504
transform 1 0 1644 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_1674
timestamp 1713400504
transform 1 0 1564 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_1675
timestamp 1713400504
transform 1 0 1836 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1676
timestamp 1713400504
transform 1 0 1756 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1677
timestamp 1713400504
transform 1 0 1948 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1678
timestamp 1713400504
transform 1 0 1860 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1679
timestamp 1713400504
transform 1 0 1804 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1680
timestamp 1713400504
transform 1 0 1764 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1681
timestamp 1713400504
transform 1 0 1772 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1682
timestamp 1713400504
transform 1 0 1700 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1683
timestamp 1713400504
transform 1 0 1716 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1684
timestamp 1713400504
transform 1 0 1604 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1685
timestamp 1713400504
transform 1 0 1900 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1686
timestamp 1713400504
transform 1 0 1844 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1687
timestamp 1713400504
transform 1 0 2620 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1688
timestamp 1713400504
transform 1 0 2484 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1689
timestamp 1713400504
transform 1 0 2580 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_1690
timestamp 1713400504
transform 1 0 2532 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_1691
timestamp 1713400504
transform 1 0 2948 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1692
timestamp 1713400504
transform 1 0 2820 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1693
timestamp 1713400504
transform 1 0 2348 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_1694
timestamp 1713400504
transform 1 0 2252 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_1695
timestamp 1713400504
transform 1 0 2492 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_1696
timestamp 1713400504
transform 1 0 2324 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_1697
timestamp 1713400504
transform 1 0 2412 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1698
timestamp 1713400504
transform 1 0 2132 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1699
timestamp 1713400504
transform 1 0 2092 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1700
timestamp 1713400504
transform 1 0 2052 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1701
timestamp 1713400504
transform 1 0 2020 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_1702
timestamp 1713400504
transform 1 0 1932 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_1703
timestamp 1713400504
transform 1 0 2196 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1704
timestamp 1713400504
transform 1 0 2092 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1705
timestamp 1713400504
transform 1 0 2028 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1706
timestamp 1713400504
transform 1 0 2108 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_1707
timestamp 1713400504
transform 1 0 2076 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_1708
timestamp 1713400504
transform 1 0 2316 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1709
timestamp 1713400504
transform 1 0 2156 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1710
timestamp 1713400504
transform 1 0 2260 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1711
timestamp 1713400504
transform 1 0 2212 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1712
timestamp 1713400504
transform 1 0 2188 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_1713
timestamp 1713400504
transform 1 0 2140 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_1714
timestamp 1713400504
transform 1 0 2164 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_1715
timestamp 1713400504
transform 1 0 2084 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_1716
timestamp 1713400504
transform 1 0 2180 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1717
timestamp 1713400504
transform 1 0 2076 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1718
timestamp 1713400504
transform 1 0 2276 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_1719
timestamp 1713400504
transform 1 0 2148 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_1720
timestamp 1713400504
transform 1 0 2132 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1721
timestamp 1713400504
transform 1 0 2068 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1722
timestamp 1713400504
transform 1 0 2972 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1723
timestamp 1713400504
transform 1 0 2900 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1724
timestamp 1713400504
transform 1 0 2860 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1725
timestamp 1713400504
transform 1 0 2780 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1726
timestamp 1713400504
transform 1 0 2756 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1727
timestamp 1713400504
transform 1 0 2716 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1728
timestamp 1713400504
transform 1 0 2764 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1729
timestamp 1713400504
transform 1 0 2692 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1730
timestamp 1713400504
transform 1 0 2732 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1731
timestamp 1713400504
transform 1 0 2700 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1732
timestamp 1713400504
transform 1 0 2828 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_1733
timestamp 1713400504
transform 1 0 2756 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_1734
timestamp 1713400504
transform 1 0 2868 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1735
timestamp 1713400504
transform 1 0 2836 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1736
timestamp 1713400504
transform 1 0 2788 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1737
timestamp 1713400504
transform 1 0 2660 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1738
timestamp 1713400504
transform 1 0 2580 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1739
timestamp 1713400504
transform 1 0 2804 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1740
timestamp 1713400504
transform 1 0 2572 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1741
timestamp 1713400504
transform 1 0 2876 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_1742
timestamp 1713400504
transform 1 0 2700 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_1743
timestamp 1713400504
transform 1 0 2812 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_1744
timestamp 1713400504
transform 1 0 2708 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_1745
timestamp 1713400504
transform 1 0 2108 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1746
timestamp 1713400504
transform 1 0 1964 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_1747
timestamp 1713400504
transform 1 0 268 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1748
timestamp 1713400504
transform 1 0 164 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1749
timestamp 1713400504
transform 1 0 108 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1750
timestamp 1713400504
transform 1 0 76 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1751
timestamp 1713400504
transform 1 0 516 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1752
timestamp 1713400504
transform 1 0 388 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1753
timestamp 1713400504
transform 1 0 676 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1754
timestamp 1713400504
transform 1 0 476 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1755
timestamp 1713400504
transform 1 0 476 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1756
timestamp 1713400504
transform 1 0 396 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1757
timestamp 1713400504
transform 1 0 468 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1758
timestamp 1713400504
transform 1 0 428 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1759
timestamp 1713400504
transform 1 0 228 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1760
timestamp 1713400504
transform 1 0 460 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1761
timestamp 1713400504
transform 1 0 220 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1762
timestamp 1713400504
transform 1 0 172 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1763
timestamp 1713400504
transform 1 0 172 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1764
timestamp 1713400504
transform 1 0 444 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_1765
timestamp 1713400504
transform 1 0 316 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_1766
timestamp 1713400504
transform 1 0 508 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1767
timestamp 1713400504
transform 1 0 68 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1768
timestamp 1713400504
transform 1 0 2964 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1769
timestamp 1713400504
transform 1 0 2812 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1770
timestamp 1713400504
transform 1 0 2436 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1771
timestamp 1713400504
transform 1 0 2356 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1772
timestamp 1713400504
transform 1 0 2292 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1773
timestamp 1713400504
transform 1 0 2956 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_1774
timestamp 1713400504
transform 1 0 2876 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1775
timestamp 1713400504
transform 1 0 2988 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1776
timestamp 1713400504
transform 1 0 2996 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1777
timestamp 1713400504
transform 1 0 2612 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1778
timestamp 1713400504
transform 1 0 3004 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1779
timestamp 1713400504
transform 1 0 2876 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1780
timestamp 1713400504
transform 1 0 2852 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1781
timestamp 1713400504
transform 1 0 2732 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1782
timestamp 1713400504
transform 1 0 2708 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1783
timestamp 1713400504
transform 1 0 2580 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1784
timestamp 1713400504
transform 1 0 3020 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_1785
timestamp 1713400504
transform 1 0 2908 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1786
timestamp 1713400504
transform 1 0 3020 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_1787
timestamp 1713400504
transform 1 0 2892 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1788
timestamp 1713400504
transform 1 0 3004 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1789
timestamp 1713400504
transform 1 0 2980 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1790
timestamp 1713400504
transform 1 0 2892 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1791
timestamp 1713400504
transform 1 0 2852 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1792
timestamp 1713400504
transform 1 0 2788 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1793
timestamp 1713400504
transform 1 0 2684 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1794
timestamp 1713400504
transform 1 0 2628 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1795
timestamp 1713400504
transform 1 0 2628 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1796
timestamp 1713400504
transform 1 0 2532 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1797
timestamp 1713400504
transform 1 0 2092 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_1798
timestamp 1713400504
transform 1 0 1972 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_1799
timestamp 1713400504
transform 1 0 1884 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_1800
timestamp 1713400504
transform 1 0 1932 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1801
timestamp 1713400504
transform 1 0 1876 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1802
timestamp 1713400504
transform 1 0 1788 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1803
timestamp 1713400504
transform 1 0 1788 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1804
timestamp 1713400504
transform 1 0 1748 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1805
timestamp 1713400504
transform 1 0 1828 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1806
timestamp 1713400504
transform 1 0 1780 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_1807
timestamp 1713400504
transform 1 0 1756 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_1808
timestamp 1713400504
transform 1 0 1260 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_1809
timestamp 1713400504
transform 1 0 1132 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_1810
timestamp 1713400504
transform 1 0 1060 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_1811
timestamp 1713400504
transform 1 0 1484 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1812
timestamp 1713400504
transform 1 0 1332 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1813
timestamp 1713400504
transform 1 0 1252 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1814
timestamp 1713400504
transform 1 0 1196 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1815
timestamp 1713400504
transform 1 0 1700 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_1816
timestamp 1713400504
transform 1 0 1668 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_1817
timestamp 1713400504
transform 1 0 1588 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_1818
timestamp 1713400504
transform 1 0 1556 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_1819
timestamp 1713400504
transform 1 0 1540 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1820
timestamp 1713400504
transform 1 0 1468 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_1821
timestamp 1713400504
transform 1 0 1452 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1822
timestamp 1713400504
transform 1 0 1404 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_1823
timestamp 1713400504
transform 1 0 1404 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1824
timestamp 1713400504
transform 1 0 1404 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1825
timestamp 1713400504
transform 1 0 1692 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_1826
timestamp 1713400504
transform 1 0 1692 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1827
timestamp 1713400504
transform 1 0 1636 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_1828
timestamp 1713400504
transform 1 0 1564 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1829
timestamp 1713400504
transform 1 0 2300 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1830
timestamp 1713400504
transform 1 0 2092 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_1831
timestamp 1713400504
transform 1 0 2092 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1832
timestamp 1713400504
transform 1 0 2028 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_1833
timestamp 1713400504
transform 1 0 2028 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_1834
timestamp 1713400504
transform 1 0 1948 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_1835
timestamp 1713400504
transform 1 0 1756 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1836
timestamp 1713400504
transform 1 0 2972 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1837
timestamp 1713400504
transform 1 0 2972 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1838
timestamp 1713400504
transform 1 0 2244 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1839
timestamp 1713400504
transform 1 0 1876 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1840
timestamp 1713400504
transform 1 0 2292 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1841
timestamp 1713400504
transform 1 0 2964 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1842
timestamp 1713400504
transform 1 0 2876 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1843
timestamp 1713400504
transform 1 0 2980 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1844
timestamp 1713400504
transform 1 0 2860 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1845
timestamp 1713400504
transform 1 0 2860 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1846
timestamp 1713400504
transform 1 0 2716 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1847
timestamp 1713400504
transform 1 0 2652 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1848
timestamp 1713400504
transform 1 0 2636 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1849
timestamp 1713400504
transform 1 0 2484 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1850
timestamp 1713400504
transform 1 0 2516 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1851
timestamp 1713400504
transform 1 0 2476 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1852
timestamp 1713400504
transform 1 0 2396 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1853
timestamp 1713400504
transform 1 0 2540 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1854
timestamp 1713400504
transform 1 0 2500 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1855
timestamp 1713400504
transform 1 0 2412 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1856
timestamp 1713400504
transform 1 0 2844 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1857
timestamp 1713400504
transform 1 0 2700 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1858
timestamp 1713400504
transform 1 0 2812 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_1859
timestamp 1713400504
transform 1 0 2812 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1860
timestamp 1713400504
transform 1 0 2740 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_1861
timestamp 1713400504
transform 1 0 2836 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1862
timestamp 1713400504
transform 1 0 2292 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1863
timestamp 1713400504
transform 1 0 2172 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1864
timestamp 1713400504
transform 1 0 2460 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1865
timestamp 1713400504
transform 1 0 2380 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1866
timestamp 1713400504
transform 1 0 2308 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_1867
timestamp 1713400504
transform 1 0 2196 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_1868
timestamp 1713400504
transform 1 0 2076 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_1869
timestamp 1713400504
transform 1 0 1868 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_1870
timestamp 1713400504
transform 1 0 2060 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1871
timestamp 1713400504
transform 1 0 1948 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1872
timestamp 1713400504
transform 1 0 1916 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1873
timestamp 1713400504
transform 1 0 1764 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_1874
timestamp 1713400504
transform 1 0 2068 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1875
timestamp 1713400504
transform 1 0 1964 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1876
timestamp 1713400504
transform 1 0 1892 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1877
timestamp 1713400504
transform 1 0 1820 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1878
timestamp 1713400504
transform 1 0 1628 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1879
timestamp 1713400504
transform 1 0 1508 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1880
timestamp 1713400504
transform 1 0 1452 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1881
timestamp 1713400504
transform 1 0 1412 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1882
timestamp 1713400504
transform 1 0 1524 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1883
timestamp 1713400504
transform 1 0 1444 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1884
timestamp 1713400504
transform 1 0 1644 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1885
timestamp 1713400504
transform 1 0 1580 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1886
timestamp 1713400504
transform 1 0 1548 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1887
timestamp 1713400504
transform 1 0 1436 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_1888
timestamp 1713400504
transform 1 0 1412 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1889
timestamp 1713400504
transform 1 0 1396 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_1890
timestamp 1713400504
transform 1 0 1340 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1891
timestamp 1713400504
transform 1 0 1596 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_1892
timestamp 1713400504
transform 1 0 1452 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_1893
timestamp 1713400504
transform 1 0 2444 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1894
timestamp 1713400504
transform 1 0 1884 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1895
timestamp 1713400504
transform 1 0 1788 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1896
timestamp 1713400504
transform 1 0 1660 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1897
timestamp 1713400504
transform 1 0 1548 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1898
timestamp 1713400504
transform 1 0 1892 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_1899
timestamp 1713400504
transform 1 0 1772 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_1900
timestamp 1713400504
transform 1 0 1724 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_1901
timestamp 1713400504
transform 1 0 1804 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1902
timestamp 1713400504
transform 1 0 1780 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1903
timestamp 1713400504
transform 1 0 1764 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1904
timestamp 1713400504
transform 1 0 1740 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1905
timestamp 1713400504
transform 1 0 1740 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1906
timestamp 1713400504
transform 1 0 2164 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_1907
timestamp 1713400504
transform 1 0 2148 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1908
timestamp 1713400504
transform 1 0 2116 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1909
timestamp 1713400504
transform 1 0 1932 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_1910
timestamp 1713400504
transform 1 0 1716 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1911
timestamp 1713400504
transform 1 0 2420 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1912
timestamp 1713400504
transform 1 0 2404 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1913
timestamp 1713400504
transform 1 0 2244 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1914
timestamp 1713400504
transform 1 0 2068 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1915
timestamp 1713400504
transform 1 0 1828 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1916
timestamp 1713400504
transform 1 0 2620 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_1917
timestamp 1713400504
transform 1 0 2580 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1918
timestamp 1713400504
transform 1 0 2444 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1919
timestamp 1713400504
transform 1 0 3004 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1920
timestamp 1713400504
transform 1 0 2820 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1921
timestamp 1713400504
transform 1 0 3012 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1922
timestamp 1713400504
transform 1 0 2812 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1923
timestamp 1713400504
transform 1 0 2868 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1924
timestamp 1713400504
transform 1 0 2764 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1925
timestamp 1713400504
transform 1 0 3004 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_1926
timestamp 1713400504
transform 1 0 2812 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1927
timestamp 1713400504
transform 1 0 2796 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1928
timestamp 1713400504
transform 1 0 2788 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_1929
timestamp 1713400504
transform 1 0 2716 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_1930
timestamp 1713400504
transform 1 0 2724 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1931
timestamp 1713400504
transform 1 0 2636 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1932
timestamp 1713400504
transform 1 0 2932 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1933
timestamp 1713400504
transform 1 0 3004 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1934
timestamp 1713400504
transform 1 0 2940 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1935
timestamp 1713400504
transform 1 0 2636 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1936
timestamp 1713400504
transform 1 0 2732 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1937
timestamp 1713400504
transform 1 0 2700 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_1938
timestamp 1713400504
transform 1 0 2668 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_1939
timestamp 1713400504
transform 1 0 2604 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_1940
timestamp 1713400504
transform 1 0 2684 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1941
timestamp 1713400504
transform 1 0 2564 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1942
timestamp 1713400504
transform 1 0 2404 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1943
timestamp 1713400504
transform 1 0 2324 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1944
timestamp 1713400504
transform 1 0 2228 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_1945
timestamp 1713400504
transform 1 0 2180 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1946
timestamp 1713400504
transform 1 0 2140 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1947
timestamp 1713400504
transform 1 0 2060 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1948
timestamp 1713400504
transform 1 0 1940 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1949
timestamp 1713400504
transform 1 0 1844 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1950
timestamp 1713400504
transform 1 0 1788 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1951
timestamp 1713400504
transform 1 0 1788 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1952
timestamp 1713400504
transform 1 0 1724 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1953
timestamp 1713400504
transform 1 0 1724 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1954
timestamp 1713400504
transform 1 0 1660 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1955
timestamp 1713400504
transform 1 0 1660 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1956
timestamp 1713400504
transform 1 0 1660 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1957
timestamp 1713400504
transform 1 0 1556 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1958
timestamp 1713400504
transform 1 0 1532 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1959
timestamp 1713400504
transform 1 0 1532 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1960
timestamp 1713400504
transform 1 0 1292 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1961
timestamp 1713400504
transform 1 0 1276 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1962
timestamp 1713400504
transform 1 0 1212 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1963
timestamp 1713400504
transform 1 0 1204 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1964
timestamp 1713400504
transform 1 0 1180 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1965
timestamp 1713400504
transform 1 0 1156 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1966
timestamp 1713400504
transform 1 0 1156 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1967
timestamp 1713400504
transform 1 0 1036 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1968
timestamp 1713400504
transform 1 0 948 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1969
timestamp 1713400504
transform 1 0 884 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1970
timestamp 1713400504
transform 1 0 1964 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1971
timestamp 1713400504
transform 1 0 1892 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1972
timestamp 1713400504
transform 1 0 1860 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1973
timestamp 1713400504
transform 1 0 1860 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1974
timestamp 1713400504
transform 1 0 1860 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1975
timestamp 1713400504
transform 1 0 1860 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1976
timestamp 1713400504
transform 1 0 1828 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_1977
timestamp 1713400504
transform 1 0 1788 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1978
timestamp 1713400504
transform 1 0 1780 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_1979
timestamp 1713400504
transform 1 0 1732 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1980
timestamp 1713400504
transform 1 0 1572 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_1981
timestamp 1713400504
transform 1 0 1516 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_1982
timestamp 1713400504
transform 1 0 1516 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1983
timestamp 1713400504
transform 1 0 1428 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_1984
timestamp 1713400504
transform 1 0 1396 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1985
timestamp 1713400504
transform 1 0 1316 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1986
timestamp 1713400504
transform 1 0 1292 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1987
timestamp 1713400504
transform 1 0 1276 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1988
timestamp 1713400504
transform 1 0 1260 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1989
timestamp 1713400504
transform 1 0 1244 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1990
timestamp 1713400504
transform 1 0 1180 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1991
timestamp 1713400504
transform 1 0 1180 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1992
timestamp 1713400504
transform 1 0 1148 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1993
timestamp 1713400504
transform 1 0 1116 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1994
timestamp 1713400504
transform 1 0 1108 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1995
timestamp 1713400504
transform 1 0 1084 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1996
timestamp 1713400504
transform 1 0 1956 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1997
timestamp 1713400504
transform 1 0 1940 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1998
timestamp 1713400504
transform 1 0 1900 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1999
timestamp 1713400504
transform 1 0 1900 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2000
timestamp 1713400504
transform 1 0 1884 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2001
timestamp 1713400504
transform 1 0 1860 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2002
timestamp 1713400504
transform 1 0 1852 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2003
timestamp 1713400504
transform 1 0 1852 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2004
timestamp 1713400504
transform 1 0 1772 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2005
timestamp 1713400504
transform 1 0 1756 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2006
timestamp 1713400504
transform 1 0 1660 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2007
timestamp 1713400504
transform 1 0 1644 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2008
timestamp 1713400504
transform 1 0 1572 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2009
timestamp 1713400504
transform 1 0 1484 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2010
timestamp 1713400504
transform 1 0 1388 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2011
timestamp 1713400504
transform 1 0 1388 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2012
timestamp 1713400504
transform 1 0 1364 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2013
timestamp 1713400504
transform 1 0 1324 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2014
timestamp 1713400504
transform 1 0 2044 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2015
timestamp 1713400504
transform 1 0 1996 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2016
timestamp 1713400504
transform 1 0 1972 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2017
timestamp 1713400504
transform 1 0 1924 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2018
timestamp 1713400504
transform 1 0 1860 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2019
timestamp 1713400504
transform 1 0 1836 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2020
timestamp 1713400504
transform 1 0 1828 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2021
timestamp 1713400504
transform 1 0 1676 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2022
timestamp 1713400504
transform 1 0 1580 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2023
timestamp 1713400504
transform 1 0 1476 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2024
timestamp 1713400504
transform 1 0 1476 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2025
timestamp 1713400504
transform 1 0 1372 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2026
timestamp 1713400504
transform 1 0 1356 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_2027
timestamp 1713400504
transform 1 0 1348 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2028
timestamp 1713400504
transform 1 0 1284 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_2029
timestamp 1713400504
transform 1 0 1948 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2030
timestamp 1713400504
transform 1 0 1924 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_2031
timestamp 1713400504
transform 1 0 1908 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_2032
timestamp 1713400504
transform 1 0 1876 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2033
timestamp 1713400504
transform 1 0 1836 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2034
timestamp 1713400504
transform 1 0 1796 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_2035
timestamp 1713400504
transform 1 0 1740 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2036
timestamp 1713400504
transform 1 0 1652 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2037
timestamp 1713400504
transform 1 0 1452 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2038
timestamp 1713400504
transform 1 0 1396 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2039
timestamp 1713400504
transform 1 0 1364 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_2040
timestamp 1713400504
transform 1 0 1340 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2041
timestamp 1713400504
transform 1 0 1340 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2042
timestamp 1713400504
transform 1 0 2020 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_2043
timestamp 1713400504
transform 1 0 1932 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_2044
timestamp 1713400504
transform 1 0 1348 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_2045
timestamp 1713400504
transform 1 0 1332 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2046
timestamp 1713400504
transform 1 0 876 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_2047
timestamp 1713400504
transform 1 0 876 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_2048
timestamp 1713400504
transform 1 0 812 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2049
timestamp 1713400504
transform 1 0 812 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2050
timestamp 1713400504
transform 1 0 772 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_2051
timestamp 1713400504
transform 1 0 756 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_2052
timestamp 1713400504
transform 1 0 716 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_2053
timestamp 1713400504
transform 1 0 716 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2054
timestamp 1713400504
transform 1 0 332 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2055
timestamp 1713400504
transform 1 0 204 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2056
timestamp 1713400504
transform 1 0 196 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2057
timestamp 1713400504
transform 1 0 1740 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_2058
timestamp 1713400504
transform 1 0 1596 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2059
timestamp 1713400504
transform 1 0 1228 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2060
timestamp 1713400504
transform 1 0 844 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_2061
timestamp 1713400504
transform 1 0 724 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2062
timestamp 1713400504
transform 1 0 724 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2063
timestamp 1713400504
transform 1 0 692 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_2064
timestamp 1713400504
transform 1 0 676 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2065
timestamp 1713400504
transform 1 0 588 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2066
timestamp 1713400504
transform 1 0 2844 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2067
timestamp 1713400504
transform 1 0 2708 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_2068
timestamp 1713400504
transform 1 0 2708 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2069
timestamp 1713400504
transform 1 0 2620 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_2070
timestamp 1713400504
transform 1 0 1596 0 1 65
box -3 -3 3 3
use M3_M2  M3_M2_2071
timestamp 1713400504
transform 1 0 1572 0 1 65
box -3 -3 3 3
use M3_M2  M3_M2_2072
timestamp 1713400504
transform 1 0 1564 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_2073
timestamp 1713400504
transform 1 0 1340 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_2074
timestamp 1713400504
transform 1 0 1092 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2075
timestamp 1713400504
transform 1 0 1052 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_2076
timestamp 1713400504
transform 1 0 924 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_2077
timestamp 1713400504
transform 1 0 924 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2078
timestamp 1713400504
transform 1 0 788 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2079
timestamp 1713400504
transform 1 0 2492 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_2080
timestamp 1713400504
transform 1 0 1700 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_2081
timestamp 1713400504
transform 1 0 1460 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2082
timestamp 1713400504
transform 1 0 1252 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2083
timestamp 1713400504
transform 1 0 1148 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2084
timestamp 1713400504
transform 1 0 1044 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_2085
timestamp 1713400504
transform 1 0 1044 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2086
timestamp 1713400504
transform 1 0 1036 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_2087
timestamp 1713400504
transform 1 0 1036 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2088
timestamp 1713400504
transform 1 0 1020 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2089
timestamp 1713400504
transform 1 0 972 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2090
timestamp 1713400504
transform 1 0 2500 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2091
timestamp 1713400504
transform 1 0 2108 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2092
timestamp 1713400504
transform 1 0 2108 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2093
timestamp 1713400504
transform 1 0 1660 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2094
timestamp 1713400504
transform 1 0 1660 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_2095
timestamp 1713400504
transform 1 0 1228 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2096
timestamp 1713400504
transform 1 0 1228 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_2097
timestamp 1713400504
transform 1 0 1212 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2098
timestamp 1713400504
transform 1 0 788 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2099
timestamp 1713400504
transform 1 0 748 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2100
timestamp 1713400504
transform 1 0 748 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2101
timestamp 1713400504
transform 1 0 644 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2102
timestamp 1713400504
transform 1 0 644 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2103
timestamp 1713400504
transform 1 0 644 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2104
timestamp 1713400504
transform 1 0 164 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2105
timestamp 1713400504
transform 1 0 1428 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_2106
timestamp 1713400504
transform 1 0 1404 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2107
timestamp 1713400504
transform 1 0 1180 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_2108
timestamp 1713400504
transform 1 0 756 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2109
timestamp 1713400504
transform 1 0 756 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2110
timestamp 1713400504
transform 1 0 708 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2111
timestamp 1713400504
transform 1 0 692 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2112
timestamp 1713400504
transform 1 0 228 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_2113
timestamp 1713400504
transform 1 0 212 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2114
timestamp 1713400504
transform 1 0 2764 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2115
timestamp 1713400504
transform 1 0 2732 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2116
timestamp 1713400504
transform 1 0 1524 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2117
timestamp 1713400504
transform 1 0 1196 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2118
timestamp 1713400504
transform 1 0 1196 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2119
timestamp 1713400504
transform 1 0 1044 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_2120
timestamp 1713400504
transform 1 0 988 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_2121
timestamp 1713400504
transform 1 0 892 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2122
timestamp 1713400504
transform 1 0 892 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2123
timestamp 1713400504
transform 1 0 860 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_2124
timestamp 1713400504
transform 1 0 844 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2125
timestamp 1713400504
transform 1 0 236 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2126
timestamp 1713400504
transform 1 0 204 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2127
timestamp 1713400504
transform 1 0 2852 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_2128
timestamp 1713400504
transform 1 0 2820 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_2129
timestamp 1713400504
transform 1 0 2820 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_2130
timestamp 1713400504
transform 1 0 2804 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_2131
timestamp 1713400504
transform 1 0 2804 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_2132
timestamp 1713400504
transform 1 0 2740 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_2133
timestamp 1713400504
transform 1 0 1484 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_2134
timestamp 1713400504
transform 1 0 1404 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2135
timestamp 1713400504
transform 1 0 1204 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_2136
timestamp 1713400504
transform 1 0 1204 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_2137
timestamp 1713400504
transform 1 0 1164 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2138
timestamp 1713400504
transform 1 0 1004 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2139
timestamp 1713400504
transform 1 0 988 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2140
timestamp 1713400504
transform 1 0 956 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_2141
timestamp 1713400504
transform 1 0 956 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2142
timestamp 1713400504
transform 1 0 796 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2143
timestamp 1713400504
transform 1 0 796 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2144
timestamp 1713400504
transform 1 0 572 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2145
timestamp 1713400504
transform 1 0 516 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2146
timestamp 1713400504
transform 1 0 2172 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2147
timestamp 1713400504
transform 1 0 2052 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_2148
timestamp 1713400504
transform 1 0 2052 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_2149
timestamp 1713400504
transform 1 0 1412 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2150
timestamp 1713400504
transform 1 0 1284 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2151
timestamp 1713400504
transform 1 0 1172 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2152
timestamp 1713400504
transform 1 0 996 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_2153
timestamp 1713400504
transform 1 0 996 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_2154
timestamp 1713400504
transform 1 0 972 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2155
timestamp 1713400504
transform 1 0 964 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_2156
timestamp 1713400504
transform 1 0 956 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2157
timestamp 1713400504
transform 1 0 708 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2158
timestamp 1713400504
transform 1 0 700 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2159
timestamp 1713400504
transform 1 0 700 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_2160
timestamp 1713400504
transform 1 0 1500 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2161
timestamp 1713400504
transform 1 0 1340 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2162
timestamp 1713400504
transform 1 0 1244 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2163
timestamp 1713400504
transform 1 0 1244 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2164
timestamp 1713400504
transform 1 0 1108 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2165
timestamp 1713400504
transform 1 0 1108 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2166
timestamp 1713400504
transform 1 0 932 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2167
timestamp 1713400504
transform 1 0 932 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2168
timestamp 1713400504
transform 1 0 868 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2169
timestamp 1713400504
transform 1 0 668 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2170
timestamp 1713400504
transform 1 0 668 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2171
timestamp 1713400504
transform 1 0 2564 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_2172
timestamp 1713400504
transform 1 0 2556 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_2173
timestamp 1713400504
transform 1 0 2516 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_2174
timestamp 1713400504
transform 1 0 2388 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_2175
timestamp 1713400504
transform 1 0 1564 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_2176
timestamp 1713400504
transform 1 0 1428 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2177
timestamp 1713400504
transform 1 0 1388 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2178
timestamp 1713400504
transform 1 0 1260 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_2179
timestamp 1713400504
transform 1 0 1220 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2180
timestamp 1713400504
transform 1 0 1188 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2181
timestamp 1713400504
transform 1 0 1188 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2182
timestamp 1713400504
transform 1 0 1188 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2183
timestamp 1713400504
transform 1 0 1172 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2184
timestamp 1713400504
transform 1 0 1156 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2185
timestamp 1713400504
transform 1 0 1140 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_2186
timestamp 1713400504
transform 1 0 1076 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2187
timestamp 1713400504
transform 1 0 1060 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_2188
timestamp 1713400504
transform 1 0 1060 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2189
timestamp 1713400504
transform 1 0 2556 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_2190
timestamp 1713400504
transform 1 0 2452 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_2191
timestamp 1713400504
transform 1 0 2156 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_2192
timestamp 1713400504
transform 1 0 2148 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_2193
timestamp 1713400504
transform 1 0 1524 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_2194
timestamp 1713400504
transform 1 0 1492 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2195
timestamp 1713400504
transform 1 0 1164 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_2196
timestamp 1713400504
transform 1 0 1164 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_2197
timestamp 1713400504
transform 1 0 1156 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2198
timestamp 1713400504
transform 1 0 1124 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2199
timestamp 1713400504
transform 1 0 1124 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_2200
timestamp 1713400504
transform 1 0 1124 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2201
timestamp 1713400504
transform 1 0 1124 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_2202
timestamp 1713400504
transform 1 0 1084 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_2203
timestamp 1713400504
transform 1 0 996 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_2204
timestamp 1713400504
transform 1 0 1892 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_2205
timestamp 1713400504
transform 1 0 1868 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_2206
timestamp 1713400504
transform 1 0 1860 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_2207
timestamp 1713400504
transform 1 0 1676 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2208
timestamp 1713400504
transform 1 0 1644 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_2209
timestamp 1713400504
transform 1 0 1636 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2210
timestamp 1713400504
transform 1 0 1516 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2211
timestamp 1713400504
transform 1 0 1308 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2212
timestamp 1713400504
transform 1 0 1116 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_2213
timestamp 1713400504
transform 1 0 1116 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_2214
timestamp 1713400504
transform 1 0 1076 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2215
timestamp 1713400504
transform 1 0 1036 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2216
timestamp 1713400504
transform 1 0 1020 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_2217
timestamp 1713400504
transform 1 0 1012 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2218
timestamp 1713400504
transform 1 0 1012 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2219
timestamp 1713400504
transform 1 0 996 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2220
timestamp 1713400504
transform 1 0 1956 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_2221
timestamp 1713400504
transform 1 0 1724 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_2222
timestamp 1713400504
transform 1 0 1676 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_2223
timestamp 1713400504
transform 1 0 1628 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2224
timestamp 1713400504
transform 1 0 1500 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2225
timestamp 1713400504
transform 1 0 1500 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_2226
timestamp 1713400504
transform 1 0 1276 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_2227
timestamp 1713400504
transform 1 0 1276 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_2228
timestamp 1713400504
transform 1 0 1228 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2229
timestamp 1713400504
transform 1 0 1012 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_2230
timestamp 1713400504
transform 1 0 1012 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_2231
timestamp 1713400504
transform 1 0 988 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2232
timestamp 1713400504
transform 1 0 940 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_2233
timestamp 1713400504
transform 1 0 924 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_2234
timestamp 1713400504
transform 1 0 692 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2235
timestamp 1713400504
transform 1 0 692 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2236
timestamp 1713400504
transform 1 0 580 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2237
timestamp 1713400504
transform 1 0 1836 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_2238
timestamp 1713400504
transform 1 0 1604 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2239
timestamp 1713400504
transform 1 0 1244 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_2240
timestamp 1713400504
transform 1 0 1140 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_2241
timestamp 1713400504
transform 1 0 1108 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2242
timestamp 1713400504
transform 1 0 1100 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_2243
timestamp 1713400504
transform 1 0 1092 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2244
timestamp 1713400504
transform 1 0 1028 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2245
timestamp 1713400504
transform 1 0 1020 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_2246
timestamp 1713400504
transform 1 0 964 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2247
timestamp 1713400504
transform 1 0 860 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_2248
timestamp 1713400504
transform 1 0 1468 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2249
timestamp 1713400504
transform 1 0 1460 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_2250
timestamp 1713400504
transform 1 0 1356 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_2251
timestamp 1713400504
transform 1 0 1156 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_2252
timestamp 1713400504
transform 1 0 1100 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_2253
timestamp 1713400504
transform 1 0 1004 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2254
timestamp 1713400504
transform 1 0 868 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2255
timestamp 1713400504
transform 1 0 860 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2256
timestamp 1713400504
transform 1 0 604 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_2257
timestamp 1713400504
transform 1 0 1492 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2258
timestamp 1713400504
transform 1 0 1436 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_2259
timestamp 1713400504
transform 1 0 1388 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2260
timestamp 1713400504
transform 1 0 1212 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_2261
timestamp 1713400504
transform 1 0 1068 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_2262
timestamp 1713400504
transform 1 0 956 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_2263
timestamp 1713400504
transform 1 0 908 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2264
timestamp 1713400504
transform 1 0 884 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2265
timestamp 1713400504
transform 1 0 596 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2266
timestamp 1713400504
transform 1 0 596 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2267
timestamp 1713400504
transform 1 0 580 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_2268
timestamp 1713400504
transform 1 0 572 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2269
timestamp 1713400504
transform 1 0 556 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2270
timestamp 1713400504
transform 1 0 68 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_2271
timestamp 1713400504
transform 1 0 4 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_2272
timestamp 1713400504
transform 1 0 1316 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_2273
timestamp 1713400504
transform 1 0 1244 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2274
timestamp 1713400504
transform 1 0 1132 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2275
timestamp 1713400504
transform 1 0 852 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2276
timestamp 1713400504
transform 1 0 852 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_2277
timestamp 1713400504
transform 1 0 836 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2278
timestamp 1713400504
transform 1 0 620 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2279
timestamp 1713400504
transform 1 0 620 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2280
timestamp 1713400504
transform 1 0 500 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2281
timestamp 1713400504
transform 1 0 460 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_2282
timestamp 1713400504
transform 1 0 1476 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2283
timestamp 1713400504
transform 1 0 1476 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2284
timestamp 1713400504
transform 1 0 1364 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2285
timestamp 1713400504
transform 1 0 1332 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2286
timestamp 1713400504
transform 1 0 1332 0 1 65
box -3 -3 3 3
use M3_M2  M3_M2_2287
timestamp 1713400504
transform 1 0 1292 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_2288
timestamp 1713400504
transform 1 0 1204 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_2289
timestamp 1713400504
transform 1 0 1204 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2290
timestamp 1713400504
transform 1 0 1172 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_2291
timestamp 1713400504
transform 1 0 1172 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2292
timestamp 1713400504
transform 1 0 1172 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2293
timestamp 1713400504
transform 1 0 988 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_2294
timestamp 1713400504
transform 1 0 916 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2295
timestamp 1713400504
transform 1 0 916 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2296
timestamp 1713400504
transform 1 0 908 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2297
timestamp 1713400504
transform 1 0 876 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2298
timestamp 1713400504
transform 1 0 876 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2299
timestamp 1713400504
transform 1 0 876 0 1 65
box -3 -3 3 3
use M3_M2  M3_M2_2300
timestamp 1713400504
transform 1 0 756 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2301
timestamp 1713400504
transform 1 0 1476 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2302
timestamp 1713400504
transform 1 0 1420 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2303
timestamp 1713400504
transform 1 0 1420 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_2304
timestamp 1713400504
transform 1 0 1268 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2305
timestamp 1713400504
transform 1 0 1116 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2306
timestamp 1713400504
transform 1 0 1108 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2307
timestamp 1713400504
transform 1 0 940 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2308
timestamp 1713400504
transform 1 0 940 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_2309
timestamp 1713400504
transform 1 0 908 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2310
timestamp 1713400504
transform 1 0 908 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2311
timestamp 1713400504
transform 1 0 900 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_2312
timestamp 1713400504
transform 1 0 836 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2313
timestamp 1713400504
transform 1 0 836 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2314
timestamp 1713400504
transform 1 0 828 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_2315
timestamp 1713400504
transform 1 0 116 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2316
timestamp 1713400504
transform 1 0 116 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2317
timestamp 1713400504
transform 1 0 1484 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2318
timestamp 1713400504
transform 1 0 1420 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2319
timestamp 1713400504
transform 1 0 1020 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2320
timestamp 1713400504
transform 1 0 1020 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2321
timestamp 1713400504
transform 1 0 1020 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2322
timestamp 1713400504
transform 1 0 956 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2323
timestamp 1713400504
transform 1 0 820 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2324
timestamp 1713400504
transform 1 0 804 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2325
timestamp 1713400504
transform 1 0 756 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_2326
timestamp 1713400504
transform 1 0 668 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_2327
timestamp 1713400504
transform 1 0 668 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2328
timestamp 1713400504
transform 1 0 668 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2329
timestamp 1713400504
transform 1 0 1668 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_2330
timestamp 1713400504
transform 1 0 1588 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_2331
timestamp 1713400504
transform 1 0 1388 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2332
timestamp 1713400504
transform 1 0 804 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2333
timestamp 1713400504
transform 1 0 796 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2334
timestamp 1713400504
transform 1 0 796 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2335
timestamp 1713400504
transform 1 0 788 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2336
timestamp 1713400504
transform 1 0 764 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2337
timestamp 1713400504
transform 1 0 740 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2338
timestamp 1713400504
transform 1 0 716 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_2339
timestamp 1713400504
transform 1 0 636 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2340
timestamp 1713400504
transform 1 0 1748 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2341
timestamp 1713400504
transform 1 0 1580 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2342
timestamp 1713400504
transform 1 0 1580 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2343
timestamp 1713400504
transform 1 0 1196 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2344
timestamp 1713400504
transform 1 0 1012 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2345
timestamp 1713400504
transform 1 0 1012 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2346
timestamp 1713400504
transform 1 0 964 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2347
timestamp 1713400504
transform 1 0 916 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2348
timestamp 1713400504
transform 1 0 868 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2349
timestamp 1713400504
transform 1 0 868 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2350
timestamp 1713400504
transform 1 0 844 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2351
timestamp 1713400504
transform 1 0 580 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2352
timestamp 1713400504
transform 1 0 500 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2353
timestamp 1713400504
transform 1 0 468 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2354
timestamp 1713400504
transform 1 0 1644 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_2355
timestamp 1713400504
transform 1 0 1132 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2356
timestamp 1713400504
transform 1 0 908 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_2357
timestamp 1713400504
transform 1 0 908 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2358
timestamp 1713400504
transform 1 0 908 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_2359
timestamp 1713400504
transform 1 0 828 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2360
timestamp 1713400504
transform 1 0 828 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_2361
timestamp 1713400504
transform 1 0 828 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2362
timestamp 1713400504
transform 1 0 724 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_2363
timestamp 1713400504
transform 1 0 724 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2364
timestamp 1713400504
transform 1 0 1764 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_2365
timestamp 1713400504
transform 1 0 1388 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_2366
timestamp 1713400504
transform 1 0 300 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_2367
timestamp 1713400504
transform 1 0 300 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2368
timestamp 1713400504
transform 1 0 220 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2369
timestamp 1713400504
transform 1 0 68 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2370
timestamp 1713400504
transform 1 0 68 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2371
timestamp 1713400504
transform 1 0 2796 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2372
timestamp 1713400504
transform 1 0 2084 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2373
timestamp 1713400504
transform 1 0 1804 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2374
timestamp 1713400504
transform 1 0 1660 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2375
timestamp 1713400504
transform 1 0 2020 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2376
timestamp 1713400504
transform 1 0 1964 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2377
timestamp 1713400504
transform 1 0 1812 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2378
timestamp 1713400504
transform 1 0 1564 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2379
timestamp 1713400504
transform 1 0 1716 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2380
timestamp 1713400504
transform 1 0 1700 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_2381
timestamp 1713400504
transform 1 0 2932 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2382
timestamp 1713400504
transform 1 0 2852 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2383
timestamp 1713400504
transform 1 0 2844 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_2384
timestamp 1713400504
transform 1 0 2772 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_2385
timestamp 1713400504
transform 1 0 2956 0 1 75
box -3 -3 3 3
use M3_M2  M3_M2_2386
timestamp 1713400504
transform 1 0 2836 0 1 75
box -3 -3 3 3
use M3_M2  M3_M2_2387
timestamp 1713400504
transform 1 0 2788 0 1 75
box -3 -3 3 3
use M3_M2  M3_M2_2388
timestamp 1713400504
transform 1 0 2620 0 1 75
box -3 -3 3 3
use M3_M2  M3_M2_2389
timestamp 1713400504
transform 1 0 2988 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_2390
timestamp 1713400504
transform 1 0 2924 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_2391
timestamp 1713400504
transform 1 0 2772 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_2392
timestamp 1713400504
transform 1 0 2628 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2393
timestamp 1713400504
transform 1 0 2556 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2394
timestamp 1713400504
transform 1 0 2900 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2395
timestamp 1713400504
transform 1 0 2804 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2396
timestamp 1713400504
transform 1 0 2708 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2397
timestamp 1713400504
transform 1 0 2612 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2398
timestamp 1713400504
transform 1 0 2612 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2399
timestamp 1713400504
transform 1 0 2556 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2400
timestamp 1713400504
transform 1 0 2964 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2401
timestamp 1713400504
transform 1 0 2892 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2402
timestamp 1713400504
transform 1 0 2756 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2403
timestamp 1713400504
transform 1 0 2756 0 1 45
box -3 -3 3 3
use M3_M2  M3_M2_2404
timestamp 1713400504
transform 1 0 2652 0 1 45
box -3 -3 3 3
use M3_M2  M3_M2_2405
timestamp 1713400504
transform 1 0 2548 0 1 45
box -3 -3 3 3
use M3_M2  M3_M2_2406
timestamp 1713400504
transform 1 0 276 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_2407
timestamp 1713400504
transform 1 0 212 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2408
timestamp 1713400504
transform 1 0 276 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_2409
timestamp 1713400504
transform 1 0 300 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_2410
timestamp 1713400504
transform 1 0 228 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2411
timestamp 1713400504
transform 1 0 292 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2412
timestamp 1713400504
transform 1 0 2996 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2413
timestamp 1713400504
transform 1 0 2692 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2414
timestamp 1713400504
transform 1 0 2164 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_2415
timestamp 1713400504
transform 1 0 732 0 1 1465
box -3 -3 3 3
use MUX2X1  MUX2X1_0
timestamp 1713400504
transform 1 0 1000 0 -1 2770
box -5 -3 53 105
use MUX2X1  MUX2X1_1
timestamp 1713400504
transform 1 0 904 0 1 2770
box -5 -3 53 105
use MUX2X1  MUX2X1_2
timestamp 1713400504
transform 1 0 784 0 1 2770
box -5 -3 53 105
use MUX2X1  MUX2X1_3
timestamp 1713400504
transform 1 0 664 0 1 2770
box -5 -3 53 105
use MUX2X1  MUX2X1_4
timestamp 1713400504
transform 1 0 616 0 1 2570
box -5 -3 53 105
use MUX2X1  MUX2X1_5
timestamp 1713400504
transform 1 0 776 0 -1 2970
box -5 -3 53 105
use MUX2X1  MUX2X1_6
timestamp 1713400504
transform 1 0 616 0 -1 2970
box -5 -3 53 105
use MUX2X1  MUX2X1_7
timestamp 1713400504
transform 1 0 480 0 1 2770
box -5 -3 53 105
use MUX2X1  MUX2X1_8
timestamp 1713400504
transform 1 0 464 0 -1 2770
box -5 -3 53 105
use MUX2X1  MUX2X1_9
timestamp 1713400504
transform 1 0 472 0 1 2570
box -5 -3 53 105
use MUX2X1  MUX2X1_10
timestamp 1713400504
transform 1 0 248 0 -1 2970
box -5 -3 53 105
use MUX2X1  MUX2X1_11
timestamp 1713400504
transform 1 0 280 0 1 2770
box -5 -3 53 105
use MUX2X1  MUX2X1_12
timestamp 1713400504
transform 1 0 264 0 -1 2770
box -5 -3 53 105
use MUX2X1  MUX2X1_13
timestamp 1713400504
transform 1 0 240 0 1 2570
box -5 -3 53 105
use MUX2X1  MUX2X1_14
timestamp 1713400504
transform 1 0 304 0 -1 2570
box -5 -3 53 105
use MUX2X1  MUX2X1_15
timestamp 1713400504
transform 1 0 80 0 1 2770
box -5 -3 53 105
use MUX2X1  MUX2X1_16
timestamp 1713400504
transform 1 0 80 0 -1 2770
box -5 -3 53 105
use MUX2X1  MUX2X1_17
timestamp 1713400504
transform 1 0 96 0 -1 2570
box -5 -3 53 105
use MUX2X1  MUX2X1_18
timestamp 1713400504
transform 1 0 136 0 1 2370
box -5 -3 53 105
use MUX2X1  MUX2X1_19
timestamp 1713400504
transform 1 0 176 0 -1 2370
box -5 -3 53 105
use MUX2X1  MUX2X1_20
timestamp 1713400504
transform 1 0 176 0 -1 2170
box -5 -3 53 105
use MUX2X1  MUX2X1_21
timestamp 1713400504
transform 1 0 184 0 1 1970
box -5 -3 53 105
use MUX2X1  MUX2X1_22
timestamp 1713400504
transform 1 0 120 0 1 1770
box -5 -3 53 105
use MUX2X1  MUX2X1_23
timestamp 1713400504
transform 1 0 256 0 1 1770
box -5 -3 53 105
use MUX2X1  MUX2X1_24
timestamp 1713400504
transform 1 0 344 0 1 1770
box -5 -3 53 105
use NAND2X1  NAND2X1_0
timestamp 1713400504
transform 1 0 96 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_1
timestamp 1713400504
transform 1 0 184 0 1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_2
timestamp 1713400504
transform 1 0 408 0 -1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_3
timestamp 1713400504
transform 1 0 568 0 -1 2970
box -8 -3 32 105
use NAND2X1  NAND2X1_4
timestamp 1713400504
transform 1 0 856 0 -1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_5
timestamp 1713400504
transform 1 0 952 0 -1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_6
timestamp 1713400504
transform 1 0 1240 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_7
timestamp 1713400504
transform 1 0 1952 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_8
timestamp 1713400504
transform 1 0 1904 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_9
timestamp 1713400504
transform 1 0 1952 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_10
timestamp 1713400504
transform 1 0 1920 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_11
timestamp 1713400504
transform 1 0 912 0 -1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_12
timestamp 1713400504
transform 1 0 1656 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_13
timestamp 1713400504
transform 1 0 88 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_14
timestamp 1713400504
transform 1 0 728 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_15
timestamp 1713400504
transform 1 0 600 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_16
timestamp 1713400504
transform 1 0 736 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_17
timestamp 1713400504
transform 1 0 800 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_18
timestamp 1713400504
transform 1 0 896 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_19
timestamp 1713400504
transform 1 0 496 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_20
timestamp 1713400504
transform 1 0 752 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_21
timestamp 1713400504
transform 1 0 448 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_22
timestamp 1713400504
transform 1 0 456 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_23
timestamp 1713400504
transform 1 0 552 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_24
timestamp 1713400504
transform 1 0 600 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_25
timestamp 1713400504
transform 1 0 888 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_26
timestamp 1713400504
transform 1 0 584 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_27
timestamp 1713400504
transform 1 0 1072 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_28
timestamp 1713400504
transform 1 0 1120 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_29
timestamp 1713400504
transform 1 0 544 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_30
timestamp 1713400504
transform 1 0 1072 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_31
timestamp 1713400504
transform 1 0 600 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_32
timestamp 1713400504
transform 1 0 648 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_33
timestamp 1713400504
transform 1 0 680 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_34
timestamp 1713400504
transform 1 0 600 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_35
timestamp 1713400504
transform 1 0 256 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_36
timestamp 1713400504
transform 1 0 328 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_37
timestamp 1713400504
transform 1 0 256 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_38
timestamp 1713400504
transform 1 0 184 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_39
timestamp 1713400504
transform 1 0 264 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_40
timestamp 1713400504
transform 1 0 1008 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_41
timestamp 1713400504
transform 1 0 400 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_42
timestamp 1713400504
transform 1 0 784 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_43
timestamp 1713400504
transform 1 0 344 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_44
timestamp 1713400504
transform 1 0 552 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_45
timestamp 1713400504
transform 1 0 200 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_46
timestamp 1713400504
transform 1 0 208 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_47
timestamp 1713400504
transform 1 0 328 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_48
timestamp 1713400504
transform 1 0 488 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_49
timestamp 1713400504
transform 1 0 344 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_50
timestamp 1713400504
transform 1 0 248 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_51
timestamp 1713400504
transform 1 0 1536 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_52
timestamp 1713400504
transform 1 0 1280 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_53
timestamp 1713400504
transform 1 0 2432 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_54
timestamp 1713400504
transform 1 0 2280 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_55
timestamp 1713400504
transform 1 0 2208 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_56
timestamp 1713400504
transform 1 0 2616 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_57
timestamp 1713400504
transform 1 0 2440 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_58
timestamp 1713400504
transform 1 0 2280 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_59
timestamp 1713400504
transform 1 0 2600 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_60
timestamp 1713400504
transform 1 0 1816 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_61
timestamp 1713400504
transform 1 0 2864 0 -1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_62
timestamp 1713400504
transform 1 0 2936 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_63
timestamp 1713400504
transform 1 0 1576 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_64
timestamp 1713400504
transform 1 0 1336 0 1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_65
timestamp 1713400504
transform 1 0 2584 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_66
timestamp 1713400504
transform 1 0 2152 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_67
timestamp 1713400504
transform 1 0 2392 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_68
timestamp 1713400504
transform 1 0 2344 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_69
timestamp 1713400504
transform 1 0 2328 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_70
timestamp 1713400504
transform 1 0 2296 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_71
timestamp 1713400504
transform 1 0 2392 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_72
timestamp 1713400504
transform 1 0 2376 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_73
timestamp 1713400504
transform 1 0 2360 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_74
timestamp 1713400504
transform 1 0 2368 0 -1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_75
timestamp 1713400504
transform 1 0 2248 0 1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_76
timestamp 1713400504
transform 1 0 2320 0 -1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_77
timestamp 1713400504
transform 1 0 2296 0 1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_78
timestamp 1713400504
transform 1 0 2192 0 1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_79
timestamp 1713400504
transform 1 0 2104 0 1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_80
timestamp 1713400504
transform 1 0 2056 0 -1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_81
timestamp 1713400504
transform 1 0 1840 0 -1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_82
timestamp 1713400504
transform 1 0 1872 0 1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_83
timestamp 1713400504
transform 1 0 1920 0 1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_84
timestamp 1713400504
transform 1 0 1816 0 -1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_85
timestamp 1713400504
transform 1 0 1904 0 -1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_86
timestamp 1713400504
transform 1 0 1840 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_87
timestamp 1713400504
transform 1 0 1984 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_88
timestamp 1713400504
transform 1 0 1856 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_89
timestamp 1713400504
transform 1 0 2016 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_90
timestamp 1713400504
transform 1 0 2024 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_91
timestamp 1713400504
transform 1 0 2112 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_92
timestamp 1713400504
transform 1 0 2056 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_93
timestamp 1713400504
transform 1 0 1792 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_94
timestamp 1713400504
transform 1 0 1752 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_95
timestamp 1713400504
transform 1 0 1720 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_96
timestamp 1713400504
transform 1 0 1824 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_97
timestamp 1713400504
transform 1 0 1872 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_98
timestamp 1713400504
transform 1 0 1816 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_99
timestamp 1713400504
transform 1 0 2272 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_100
timestamp 1713400504
transform 1 0 1672 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_101
timestamp 1713400504
transform 1 0 1528 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_102
timestamp 1713400504
transform 1 0 1488 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_103
timestamp 1713400504
transform 1 0 1416 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_104
timestamp 1713400504
transform 1 0 1824 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_105
timestamp 1713400504
transform 1 0 1784 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_106
timestamp 1713400504
transform 1 0 1832 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_107
timestamp 1713400504
transform 1 0 848 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_108
timestamp 1713400504
transform 1 0 1136 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_109
timestamp 1713400504
transform 1 0 1032 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_110
timestamp 1713400504
transform 1 0 944 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_111
timestamp 1713400504
transform 1 0 1016 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_112
timestamp 1713400504
transform 1 0 1520 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_113
timestamp 1713400504
transform 1 0 1080 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_114
timestamp 1713400504
transform 1 0 1160 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_115
timestamp 1713400504
transform 1 0 1112 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_116
timestamp 1713400504
transform 1 0 1192 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_117
timestamp 1713400504
transform 1 0 736 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_118
timestamp 1713400504
transform 1 0 1152 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_119
timestamp 1713400504
transform 1 0 1088 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_120
timestamp 1713400504
transform 1 0 920 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_121
timestamp 1713400504
transform 1 0 984 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_122
timestamp 1713400504
transform 1 0 952 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_123
timestamp 1713400504
transform 1 0 1032 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_124
timestamp 1713400504
transform 1 0 1136 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_125
timestamp 1713400504
transform 1 0 1088 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_126
timestamp 1713400504
transform 1 0 1160 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_127
timestamp 1713400504
transform 1 0 2016 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_128
timestamp 1713400504
transform 1 0 2080 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_129
timestamp 1713400504
transform 1 0 2696 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_130
timestamp 1713400504
transform 1 0 2048 0 -1 370
box -8 -3 32 105
use NAND3X1  NAND3X1_0
timestamp 1713400504
transform 1 0 1952 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_1
timestamp 1713400504
transform 1 0 1880 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_2
timestamp 1713400504
transform 1 0 1816 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_3
timestamp 1713400504
transform 1 0 1992 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_4
timestamp 1713400504
transform 1 0 2024 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_5
timestamp 1713400504
transform 1 0 2016 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_6
timestamp 1713400504
transform 1 0 1632 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_7
timestamp 1713400504
transform 1 0 320 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_8
timestamp 1713400504
transform 1 0 336 0 -1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_9
timestamp 1713400504
transform 1 0 352 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_10
timestamp 1713400504
transform 1 0 272 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_11
timestamp 1713400504
transform 1 0 160 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_12
timestamp 1713400504
transform 1 0 352 0 -1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_13
timestamp 1713400504
transform 1 0 1432 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_14
timestamp 1713400504
transform 1 0 2232 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_15
timestamp 1713400504
transform 1 0 2512 0 -1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_16
timestamp 1713400504
transform 1 0 2400 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_17
timestamp 1713400504
transform 1 0 2328 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_18
timestamp 1713400504
transform 1 0 2424 0 -1 2570
box -8 -3 40 105
use NAND3X1  NAND3X1_19
timestamp 1713400504
transform 1 0 2400 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_20
timestamp 1713400504
transform 1 0 2104 0 1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_21
timestamp 1713400504
transform 1 0 2704 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_22
timestamp 1713400504
transform 1 0 1968 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_23
timestamp 1713400504
transform 1 0 2656 0 1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_24
timestamp 1713400504
transform 1 0 2128 0 1 2770
box -8 -3 40 105
use NAND3X1  NAND3X1_25
timestamp 1713400504
transform 1 0 1456 0 -1 2770
box -8 -3 40 105
use NAND3X1  NAND3X1_26
timestamp 1713400504
transform 1 0 2568 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_27
timestamp 1713400504
transform 1 0 2520 0 1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_28
timestamp 1713400504
transform 1 0 2304 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_29
timestamp 1713400504
transform 1 0 2592 0 1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_30
timestamp 1713400504
transform 1 0 2432 0 -1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_31
timestamp 1713400504
transform 1 0 2520 0 -1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_32
timestamp 1713400504
transform 1 0 2752 0 1 2570
box -8 -3 40 105
use NAND3X1  NAND3X1_33
timestamp 1713400504
transform 1 0 2960 0 1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_34
timestamp 1713400504
transform 1 0 2624 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_35
timestamp 1713400504
transform 1 0 2568 0 1 2770
box -8 -3 40 105
use NAND3X1  NAND3X1_36
timestamp 1713400504
transform 1 0 2424 0 1 2770
box -8 -3 40 105
use NAND3X1  NAND3X1_37
timestamp 1713400504
transform 1 0 2632 0 1 2770
box -8 -3 40 105
use NAND3X1  NAND3X1_38
timestamp 1713400504
transform 1 0 2672 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_39
timestamp 1713400504
transform 1 0 2896 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_40
timestamp 1713400504
transform 1 0 1728 0 1 2570
box -8 -3 40 105
use NAND3X1  NAND3X1_41
timestamp 1713400504
transform 1 0 1536 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_42
timestamp 1713400504
transform 1 0 1360 0 -1 2770
box -8 -3 40 105
use NAND3X1  NAND3X1_43
timestamp 1713400504
transform 1 0 1240 0 -1 2770
box -8 -3 40 105
use NAND3X1  NAND3X1_44
timestamp 1713400504
transform 1 0 1176 0 1 2770
box -8 -3 40 105
use NAND3X1  NAND3X1_45
timestamp 1713400504
transform 1 0 1528 0 -1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_46
timestamp 1713400504
transform 1 0 2656 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_47
timestamp 1713400504
transform 1 0 1520 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_48
timestamp 1713400504
transform 1 0 1256 0 1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_49
timestamp 1713400504
transform 1 0 2136 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_50
timestamp 1713400504
transform 1 0 1912 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_51
timestamp 1713400504
transform 1 0 2464 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_52
timestamp 1713400504
transform 1 0 2160 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_53
timestamp 1713400504
transform 1 0 2288 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_54
timestamp 1713400504
transform 1 0 2248 0 -1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_55
timestamp 1713400504
transform 1 0 2104 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_56
timestamp 1713400504
transform 1 0 2840 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_57
timestamp 1713400504
transform 1 0 2960 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_58
timestamp 1713400504
transform 1 0 2712 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_59
timestamp 1713400504
transform 1 0 2784 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_60
timestamp 1713400504
transform 1 0 2616 0 -1 170
box -8 -3 40 105
use NOR2X1  NOR2X1_0
timestamp 1713400504
transform 1 0 232 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_1
timestamp 1713400504
transform 1 0 192 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_2
timestamp 1713400504
transform 1 0 384 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_3
timestamp 1713400504
transform 1 0 584 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_4
timestamp 1713400504
transform 1 0 712 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_5
timestamp 1713400504
transform 1 0 920 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_6
timestamp 1713400504
transform 1 0 376 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_7
timestamp 1713400504
transform 1 0 448 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_8
timestamp 1713400504
transform 1 0 504 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_9
timestamp 1713400504
transform 1 0 576 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_10
timestamp 1713400504
transform 1 0 640 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_11
timestamp 1713400504
transform 1 0 368 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_12
timestamp 1713400504
transform 1 0 344 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_13
timestamp 1713400504
transform 1 0 544 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_14
timestamp 1713400504
transform 1 0 664 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_15
timestamp 1713400504
transform 1 0 680 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_16
timestamp 1713400504
transform 1 0 312 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_17
timestamp 1713400504
transform 1 0 488 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_18
timestamp 1713400504
transform 1 0 600 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_19
timestamp 1713400504
transform 1 0 752 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_20
timestamp 1713400504
transform 1 0 664 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_21
timestamp 1713400504
transform 1 0 1312 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_22
timestamp 1713400504
transform 1 0 1184 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_23
timestamp 1713400504
transform 1 0 2216 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_24
timestamp 1713400504
transform 1 0 2264 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_25
timestamp 1713400504
transform 1 0 2232 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_26
timestamp 1713400504
transform 1 0 2240 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_27
timestamp 1713400504
transform 1 0 2336 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_28
timestamp 1713400504
transform 1 0 2248 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_29
timestamp 1713400504
transform 1 0 2280 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_30
timestamp 1713400504
transform 1 0 2200 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_31
timestamp 1713400504
transform 1 0 1960 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_32
timestamp 1713400504
transform 1 0 1960 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_33
timestamp 1713400504
transform 1 0 1904 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_34
timestamp 1713400504
transform 1 0 2040 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_35
timestamp 1713400504
transform 1 0 1888 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_36
timestamp 1713400504
transform 1 0 2280 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_37
timestamp 1713400504
transform 1 0 1936 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_38
timestamp 1713400504
transform 1 0 1880 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_39
timestamp 1713400504
transform 1 0 2000 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_40
timestamp 1713400504
transform 1 0 1944 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_41
timestamp 1713400504
transform 1 0 1992 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_42
timestamp 1713400504
transform 1 0 2048 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_43
timestamp 1713400504
transform 1 0 2104 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_44
timestamp 1713400504
transform 1 0 2160 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_45
timestamp 1713400504
transform 1 0 2296 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_46
timestamp 1713400504
transform 1 0 2240 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_47
timestamp 1713400504
transform 1 0 2120 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_48
timestamp 1713400504
transform 1 0 1840 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_49
timestamp 1713400504
transform 1 0 120 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_50
timestamp 1713400504
transform 1 0 200 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_51
timestamp 1713400504
transform 1 0 408 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_52
timestamp 1713400504
transform 1 0 128 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_53
timestamp 1713400504
transform 1 0 376 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_54
timestamp 1713400504
transform 1 0 320 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_55
timestamp 1713400504
transform 1 0 216 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_56
timestamp 1713400504
transform 1 0 2296 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_57
timestamp 1713400504
transform 1 0 2336 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_58
timestamp 1713400504
transform 1 0 2432 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_59
timestamp 1713400504
transform 1 0 2320 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_60
timestamp 1713400504
transform 1 0 2424 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_61
timestamp 1713400504
transform 1 0 2392 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_62
timestamp 1713400504
transform 1 0 2184 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_63
timestamp 1713400504
transform 1 0 2344 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_64
timestamp 1713400504
transform 1 0 2152 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_65
timestamp 1713400504
transform 1 0 2736 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_66
timestamp 1713400504
transform 1 0 2520 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_67
timestamp 1713400504
transform 1 0 2472 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_68
timestamp 1713400504
transform 1 0 2536 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_69
timestamp 1713400504
transform 1 0 2632 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_70
timestamp 1713400504
transform 1 0 2552 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_71
timestamp 1713400504
transform 1 0 2496 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_72
timestamp 1713400504
transform 1 0 2760 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_73
timestamp 1713400504
transform 1 0 2600 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_74
timestamp 1713400504
transform 1 0 2616 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_75
timestamp 1713400504
transform 1 0 2528 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_76
timestamp 1713400504
transform 1 0 2624 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_77
timestamp 1713400504
transform 1 0 2800 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_78
timestamp 1713400504
transform 1 0 1784 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_79
timestamp 1713400504
transform 1 0 1736 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_80
timestamp 1713400504
transform 1 0 1816 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_81
timestamp 1713400504
transform 1 0 1304 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_82
timestamp 1713400504
transform 1 0 1760 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_83
timestamp 1713400504
transform 1 0 1864 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_84
timestamp 1713400504
transform 1 0 1488 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_85
timestamp 1713400504
transform 1 0 2544 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_86
timestamp 1713400504
transform 1 0 1536 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_87
timestamp 1713400504
transform 1 0 1352 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_88
timestamp 1713400504
transform 1 0 1824 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_89
timestamp 1713400504
transform 1 0 2432 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_90
timestamp 1713400504
transform 1 0 2384 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_91
timestamp 1713400504
transform 1 0 2040 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_92
timestamp 1713400504
transform 1 0 1640 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_93
timestamp 1713400504
transform 1 0 1552 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_94
timestamp 1713400504
transform 1 0 1824 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_95
timestamp 1713400504
transform 1 0 1600 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_96
timestamp 1713400504
transform 1 0 1552 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_97
timestamp 1713400504
transform 1 0 1688 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_98
timestamp 1713400504
transform 1 0 1776 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_99
timestamp 1713400504
transform 1 0 2192 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_100
timestamp 1713400504
transform 1 0 2296 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_101
timestamp 1713400504
transform 1 0 2888 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_102
timestamp 1713400504
transform 1 0 2600 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_103
timestamp 1713400504
transform 1 0 2640 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_104
timestamp 1713400504
transform 1 0 2968 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_105
timestamp 1713400504
transform 1 0 2880 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_106
timestamp 1713400504
transform 1 0 2552 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_107
timestamp 1713400504
transform 1 0 2656 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_108
timestamp 1713400504
transform 1 0 1984 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_109
timestamp 1713400504
transform 1 0 2424 0 -1 370
box -8 -3 32 105
use NOR3X1  NOR3X1_0
timestamp 1713400504
transform 1 0 1968 0 1 370
box -7 -3 68 105
use OAI21X1  OAI21X1_0
timestamp 1713400504
transform 1 0 1216 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_1
timestamp 1713400504
transform 1 0 1920 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_2
timestamp 1713400504
transform 1 0 1832 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_3
timestamp 1713400504
transform 1 0 152 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_4
timestamp 1713400504
transform 1 0 256 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_5
timestamp 1713400504
transform 1 0 688 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_6
timestamp 1713400504
transform 1 0 544 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_7
timestamp 1713400504
transform 1 0 544 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_8
timestamp 1713400504
transform 1 0 432 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_9
timestamp 1713400504
transform 1 0 816 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_10
timestamp 1713400504
transform 1 0 592 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_11
timestamp 1713400504
transform 1 0 872 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_12
timestamp 1713400504
transform 1 0 680 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_13
timestamp 1713400504
transform 1 0 952 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_14
timestamp 1713400504
transform 1 0 624 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_15
timestamp 1713400504
transform 1 0 816 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_16
timestamp 1713400504
transform 1 0 688 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_17
timestamp 1713400504
transform 1 0 392 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_18
timestamp 1713400504
transform 1 0 344 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_19
timestamp 1713400504
transform 1 0 528 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_20
timestamp 1713400504
transform 1 0 416 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_21
timestamp 1713400504
transform 1 0 528 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_22
timestamp 1713400504
transform 1 0 456 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_23
timestamp 1713400504
transform 1 0 872 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_24
timestamp 1713400504
transform 1 0 672 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_25
timestamp 1713400504
transform 1 0 640 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_26
timestamp 1713400504
transform 1 0 512 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_27
timestamp 1713400504
transform 1 0 968 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_28
timestamp 1713400504
transform 1 0 792 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_29
timestamp 1713400504
transform 1 0 1032 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_30
timestamp 1713400504
transform 1 0 768 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_31
timestamp 1713400504
transform 1 0 992 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_32
timestamp 1713400504
transform 1 0 760 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_33
timestamp 1713400504
transform 1 0 728 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_34
timestamp 1713400504
transform 1 0 488 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_35
timestamp 1713400504
transform 1 0 616 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_36
timestamp 1713400504
transform 1 0 496 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_37
timestamp 1713400504
transform 1 0 528 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_38
timestamp 1713400504
transform 1 0 704 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_39
timestamp 1713400504
transform 1 0 200 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_40
timestamp 1713400504
transform 1 0 296 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_41
timestamp 1713400504
transform 1 0 192 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_42
timestamp 1713400504
transform 1 0 416 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_43
timestamp 1713400504
transform 1 0 112 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_44
timestamp 1713400504
transform 1 0 336 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_45
timestamp 1713400504
transform 1 0 952 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_46
timestamp 1713400504
transform 1 0 568 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_47
timestamp 1713400504
transform 1 0 720 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_48
timestamp 1713400504
transform 1 0 368 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_49
timestamp 1713400504
transform 1 0 480 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_50
timestamp 1713400504
transform 1 0 408 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_51
timestamp 1713400504
transform 1 0 264 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_52
timestamp 1713400504
transform 1 0 304 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_53
timestamp 1713400504
transform 1 0 176 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_54
timestamp 1713400504
transform 1 0 256 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_55
timestamp 1713400504
transform 1 0 528 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_56
timestamp 1713400504
transform 1 0 336 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_57
timestamp 1713400504
transform 1 0 352 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_58
timestamp 1713400504
transform 1 0 88 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_59
timestamp 1713400504
transform 1 0 144 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_60
timestamp 1713400504
transform 1 0 1368 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_61
timestamp 1713400504
transform 1 0 2528 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_62
timestamp 1713400504
transform 1 0 2344 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_63
timestamp 1713400504
transform 1 0 2480 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_64
timestamp 1713400504
transform 1 0 2424 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_65
timestamp 1713400504
transform 1 0 2464 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_66
timestamp 1713400504
transform 1 0 2504 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_67
timestamp 1713400504
transform 1 0 2640 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_68
timestamp 1713400504
transform 1 0 2456 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_69
timestamp 1713400504
transform 1 0 1600 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_70
timestamp 1713400504
transform 1 0 1400 0 1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_71
timestamp 1713400504
transform 1 0 2560 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_72
timestamp 1713400504
transform 1 0 2824 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_73
timestamp 1713400504
transform 1 0 2880 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_74
timestamp 1713400504
transform 1 0 1968 0 1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_75
timestamp 1713400504
transform 1 0 2648 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_76
timestamp 1713400504
transform 1 0 2568 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_77
timestamp 1713400504
transform 1 0 2864 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_78
timestamp 1713400504
transform 1 0 1600 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_79
timestamp 1713400504
transform 1 0 1176 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_80
timestamp 1713400504
transform 1 0 1264 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_81
timestamp 1713400504
transform 1 0 2512 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_82
timestamp 1713400504
transform 1 0 1368 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_83
timestamp 1713400504
transform 1 0 2144 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_84
timestamp 1713400504
transform 1 0 2720 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_85
timestamp 1713400504
transform 1 0 2736 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_86
timestamp 1713400504
transform 1 0 2512 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_87
timestamp 1713400504
transform 1 0 2352 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_88
timestamp 1713400504
transform 1 0 2424 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_89
timestamp 1713400504
transform 1 0 2688 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_90
timestamp 1713400504
transform 1 0 2656 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_91
timestamp 1713400504
transform 1 0 2696 0 1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_92
timestamp 1713400504
transform 1 0 2304 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_93
timestamp 1713400504
transform 1 0 2352 0 1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_94
timestamp 1713400504
transform 1 0 2328 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_95
timestamp 1713400504
transform 1 0 2224 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_96
timestamp 1713400504
transform 1 0 2104 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_97
timestamp 1713400504
transform 1 0 2048 0 1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_98
timestamp 1713400504
transform 1 0 1640 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_99
timestamp 1713400504
transform 1 0 1512 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_100
timestamp 1713400504
transform 1 0 1576 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_101
timestamp 1713400504
transform 1 0 1568 0 1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_102
timestamp 1713400504
transform 1 0 1624 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_103
timestamp 1713400504
transform 1 0 1816 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_104
timestamp 1713400504
transform 1 0 1920 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_105
timestamp 1713400504
transform 1 0 1776 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_106
timestamp 1713400504
transform 1 0 2048 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_107
timestamp 1713400504
transform 1 0 2032 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_108
timestamp 1713400504
transform 1 0 1728 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_109
timestamp 1713400504
transform 1 0 1744 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_110
timestamp 1713400504
transform 1 0 1688 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_111
timestamp 1713400504
transform 1 0 1776 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_112
timestamp 1713400504
transform 1 0 1808 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_113
timestamp 1713400504
transform 1 0 1552 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_114
timestamp 1713400504
transform 1 0 1776 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_115
timestamp 1713400504
transform 1 0 1704 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_116
timestamp 1713400504
transform 1 0 1784 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_117
timestamp 1713400504
transform 1 0 1752 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_118
timestamp 1713400504
transform 1 0 1896 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_119
timestamp 1713400504
transform 1 0 1824 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_120
timestamp 1713400504
transform 1 0 1664 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_121
timestamp 1713400504
transform 1 0 1560 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_122
timestamp 1713400504
transform 1 0 1504 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_123
timestamp 1713400504
transform 1 0 1552 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_124
timestamp 1713400504
transform 1 0 1328 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_125
timestamp 1713400504
transform 1 0 1240 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_126
timestamp 1713400504
transform 1 0 1072 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_127
timestamp 1713400504
transform 1 0 864 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_128
timestamp 1713400504
transform 1 0 1064 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_129
timestamp 1713400504
transform 1 0 1120 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_130
timestamp 1713400504
transform 1 0 856 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_131
timestamp 1713400504
transform 1 0 832 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_132
timestamp 1713400504
transform 1 0 1584 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_133
timestamp 1713400504
transform 1 0 1504 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_134
timestamp 1713400504
transform 1 0 1264 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_135
timestamp 1713400504
transform 1 0 1256 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_136
timestamp 1713400504
transform 1 0 1336 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_137
timestamp 1713400504
transform 1 0 1384 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_138
timestamp 1713400504
transform 1 0 1360 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_139
timestamp 1713400504
transform 1 0 1440 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_140
timestamp 1713400504
transform 1 0 1456 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_141
timestamp 1713400504
transform 1 0 1360 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_142
timestamp 1713400504
transform 1 0 936 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_143
timestamp 1713400504
transform 1 0 840 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_144
timestamp 1713400504
transform 1 0 1032 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_145
timestamp 1713400504
transform 1 0 1176 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_146
timestamp 1713400504
transform 1 0 728 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_147
timestamp 1713400504
transform 1 0 640 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_148
timestamp 1713400504
transform 1 0 1376 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_149
timestamp 1713400504
transform 1 0 1304 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_150
timestamp 1713400504
transform 1 0 1040 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_151
timestamp 1713400504
transform 1 0 936 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_152
timestamp 1713400504
transform 1 0 1136 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_153
timestamp 1713400504
transform 1 0 1040 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_154
timestamp 1713400504
transform 1 0 944 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_155
timestamp 1713400504
transform 1 0 888 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_156
timestamp 1713400504
transform 1 0 2240 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_157
timestamp 1713400504
transform 1 0 2328 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_158
timestamp 1713400504
transform 1 0 1928 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_159
timestamp 1713400504
transform 1 0 2248 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_160
timestamp 1713400504
transform 1 0 2064 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_161
timestamp 1713400504
transform 1 0 2152 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_162
timestamp 1713400504
transform 1 0 2792 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_163
timestamp 1713400504
transform 1 0 2848 0 -1 170
box -8 -3 34 105
use OAI22X1  OAI22X1_0
timestamp 1713400504
transform 1 0 152 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_1
timestamp 1713400504
transform 1 0 2744 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_2
timestamp 1713400504
transform 1 0 2824 0 1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_3
timestamp 1713400504
transform 1 0 2568 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_4
timestamp 1713400504
transform 1 0 2832 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_5
timestamp 1713400504
transform 1 0 2080 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_6
timestamp 1713400504
transform 1 0 2144 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_7
timestamp 1713400504
transform 1 0 1648 0 1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_8
timestamp 1713400504
transform 1 0 1448 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_9
timestamp 1713400504
transform 1 0 1728 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_10
timestamp 1713400504
transform 1 0 1408 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_11
timestamp 1713400504
transform 1 0 1280 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_12
timestamp 1713400504
transform 1 0 1216 0 1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_13
timestamp 1713400504
transform 1 0 1328 0 -1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_14
timestamp 1713400504
transform 1 0 1216 0 -1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_15
timestamp 1713400504
transform 1 0 1784 0 -1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_16
timestamp 1713400504
transform 1 0 1984 0 -1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_17
timestamp 1713400504
transform 1 0 2152 0 -1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_18
timestamp 1713400504
transform 1 0 2432 0 -1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_19
timestamp 1713400504
transform 1 0 2744 0 -1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_20
timestamp 1713400504
transform 1 0 2704 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_21
timestamp 1713400504
transform 1 0 2880 0 -1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_22
timestamp 1713400504
transform 1 0 2944 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_23
timestamp 1713400504
transform 1 0 2840 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_24
timestamp 1713400504
transform 1 0 2632 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_25
timestamp 1713400504
transform 1 0 2656 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_26
timestamp 1713400504
transform 1 0 2784 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_27
timestamp 1713400504
transform 1 0 2896 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_28
timestamp 1713400504
transform 1 0 2920 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_29
timestamp 1713400504
transform 1 0 2792 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_30
timestamp 1713400504
transform 1 0 1992 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_31
timestamp 1713400504
transform 1 0 2096 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_32
timestamp 1713400504
transform 1 0 2272 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_33
timestamp 1713400504
transform 1 0 1912 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_34
timestamp 1713400504
transform 1 0 2032 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_35
timestamp 1713400504
transform 1 0 1904 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_36
timestamp 1713400504
transform 1 0 1696 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_37
timestamp 1713400504
transform 1 0 1864 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_38
timestamp 1713400504
transform 1 0 1920 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_39
timestamp 1713400504
transform 1 0 1584 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_40
timestamp 1713400504
transform 1 0 1792 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_41
timestamp 1713400504
transform 1 0 1688 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_42
timestamp 1713400504
transform 1 0 1056 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_43
timestamp 1713400504
transform 1 0 840 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_44
timestamp 1713400504
transform 1 0 952 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_45
timestamp 1713400504
transform 1 0 728 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_46
timestamp 1713400504
transform 1 0 992 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_47
timestamp 1713400504
transform 1 0 944 0 1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_48
timestamp 1713400504
transform 1 0 1088 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_49
timestamp 1713400504
transform 1 0 1008 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_50
timestamp 1713400504
transform 1 0 952 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_51
timestamp 1713400504
transform 1 0 848 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_52
timestamp 1713400504
transform 1 0 936 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_53
timestamp 1713400504
transform 1 0 720 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_54
timestamp 1713400504
transform 1 0 1280 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_55
timestamp 1713400504
transform 1 0 1296 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_56
timestamp 1713400504
transform 1 0 1160 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_57
timestamp 1713400504
transform 1 0 1184 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_58
timestamp 1713400504
transform 1 0 1224 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_59
timestamp 1713400504
transform 1 0 1240 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_60
timestamp 1713400504
transform 1 0 1184 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_61
timestamp 1713400504
transform 1 0 1272 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_62
timestamp 1713400504
transform 1 0 1264 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_63
timestamp 1713400504
transform 1 0 1352 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_64
timestamp 1713400504
transform 1 0 1160 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_65
timestamp 1713400504
transform 1 0 1384 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_66
timestamp 1713400504
transform 1 0 1040 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_67
timestamp 1713400504
transform 1 0 704 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_68
timestamp 1713400504
transform 1 0 816 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_69
timestamp 1713400504
transform 1 0 712 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_70
timestamp 1713400504
transform 1 0 1120 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_71
timestamp 1713400504
transform 1 0 936 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_72
timestamp 1713400504
transform 1 0 1064 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_73
timestamp 1713400504
transform 1 0 944 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_74
timestamp 1713400504
transform 1 0 824 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_75
timestamp 1713400504
transform 1 0 528 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_76
timestamp 1713400504
transform 1 0 824 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_77
timestamp 1713400504
transform 1 0 632 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_78
timestamp 1713400504
transform 1 0 968 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_79
timestamp 1713400504
transform 1 0 744 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_80
timestamp 1713400504
transform 1 0 856 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_81
timestamp 1713400504
transform 1 0 752 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_82
timestamp 1713400504
transform 1 0 1080 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_83
timestamp 1713400504
transform 1 0 1136 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_84
timestamp 1713400504
transform 1 0 928 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_85
timestamp 1713400504
transform 1 0 984 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_86
timestamp 1713400504
transform 1 0 856 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_87
timestamp 1713400504
transform 1 0 848 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_88
timestamp 1713400504
transform 1 0 808 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_89
timestamp 1713400504
transform 1 0 784 0 1 1370
box -8 -3 46 105
use OR2X1  OR2X1_0
timestamp 1713400504
transform 1 0 88 0 1 2170
box -8 -3 40 105
use OR2X1  OR2X1_1
timestamp 1713400504
transform 1 0 144 0 -1 2970
box -8 -3 40 105
use OR2X1  OR2X1_2
timestamp 1713400504
transform 1 0 424 0 -1 2970
box -8 -3 40 105
use OR2X1  OR2X1_3
timestamp 1713400504
transform 1 0 928 0 -1 2970
box -8 -3 40 105
use OR2X1  OR2X1_4
timestamp 1713400504
transform 1 0 1880 0 1 1970
box -8 -3 40 105
use OR2X1  OR2X1_5
timestamp 1713400504
transform 1 0 1640 0 -1 570
box -8 -3 40 105
use OR2X1  OR2X1_6
timestamp 1713400504
transform 1 0 1400 0 1 1570
box -8 -3 40 105
use OR2X1  OR2X1_7
timestamp 1713400504
transform 1 0 1312 0 1 1770
box -8 -3 40 105
use OR2X1  OR2X1_8
timestamp 1713400504
transform 1 0 1368 0 1 1370
box -8 -3 40 105
use OR2X1  OR2X1_9
timestamp 1713400504
transform 1 0 232 0 1 1170
box -8 -3 40 105
use OR2X1  OR2X1_10
timestamp 1713400504
transform 1 0 912 0 -1 170
box -8 -3 40 105
use OR2X1  OR2X1_11
timestamp 1713400504
transform 1 0 2152 0 1 370
box -8 -3 40 105
use OR2X1  OR2X1_12
timestamp 1713400504
transform 1 0 2728 0 -1 770
box -8 -3 40 105
use top_module_VIA0  top_module_VIA0_0
timestamp 1713400504
transform 1 0 3064 0 1 3017
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_1
timestamp 1713400504
transform 1 0 3064 0 1 23
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_2
timestamp 1713400504
transform 1 0 24 0 1 3017
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_3
timestamp 1713400504
transform 1 0 24 0 1 23
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_4
timestamp 1713400504
transform 1 0 3040 0 1 2993
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_5
timestamp 1713400504
transform 1 0 3040 0 1 47
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_6
timestamp 1713400504
transform 1 0 48 0 1 2993
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_7
timestamp 1713400504
transform 1 0 48 0 1 47
box -10 -10 10 10
use top_module_VIA1  top_module_VIA1_0
timestamp 1713400504
transform 1 0 3064 0 1 2870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_1
timestamp 1713400504
transform 1 0 3064 0 1 2670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_2
timestamp 1713400504
transform 1 0 3064 0 1 2470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_3
timestamp 1713400504
transform 1 0 3064 0 1 2270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_4
timestamp 1713400504
transform 1 0 3064 0 1 2070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_5
timestamp 1713400504
transform 1 0 3064 0 1 1870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_6
timestamp 1713400504
transform 1 0 3064 0 1 1670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_7
timestamp 1713400504
transform 1 0 3064 0 1 1470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_8
timestamp 1713400504
transform 1 0 3064 0 1 1270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_9
timestamp 1713400504
transform 1 0 3064 0 1 1070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_10
timestamp 1713400504
transform 1 0 3064 0 1 870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_11
timestamp 1713400504
transform 1 0 3064 0 1 670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_12
timestamp 1713400504
transform 1 0 3064 0 1 470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_13
timestamp 1713400504
transform 1 0 3064 0 1 270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_14
timestamp 1713400504
transform 1 0 3064 0 1 70
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_15
timestamp 1713400504
transform 1 0 24 0 1 2870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_16
timestamp 1713400504
transform 1 0 24 0 1 2670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_17
timestamp 1713400504
transform 1 0 24 0 1 2470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_18
timestamp 1713400504
transform 1 0 24 0 1 2270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_19
timestamp 1713400504
transform 1 0 24 0 1 2070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_20
timestamp 1713400504
transform 1 0 24 0 1 1870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_21
timestamp 1713400504
transform 1 0 24 0 1 1670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_22
timestamp 1713400504
transform 1 0 24 0 1 1470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_23
timestamp 1713400504
transform 1 0 24 0 1 1270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_24
timestamp 1713400504
transform 1 0 24 0 1 1070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_25
timestamp 1713400504
transform 1 0 24 0 1 870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_26
timestamp 1713400504
transform 1 0 24 0 1 670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_27
timestamp 1713400504
transform 1 0 24 0 1 470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_28
timestamp 1713400504
transform 1 0 24 0 1 270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_29
timestamp 1713400504
transform 1 0 24 0 1 70
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_30
timestamp 1713400504
transform 1 0 48 0 1 170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_31
timestamp 1713400504
transform 1 0 48 0 1 370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_32
timestamp 1713400504
transform 1 0 48 0 1 570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_33
timestamp 1713400504
transform 1 0 48 0 1 770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_34
timestamp 1713400504
transform 1 0 48 0 1 970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_35
timestamp 1713400504
transform 1 0 48 0 1 1170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_36
timestamp 1713400504
transform 1 0 48 0 1 1370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_37
timestamp 1713400504
transform 1 0 48 0 1 1570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_38
timestamp 1713400504
transform 1 0 48 0 1 1770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_39
timestamp 1713400504
transform 1 0 48 0 1 1970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_40
timestamp 1713400504
transform 1 0 48 0 1 2170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_41
timestamp 1713400504
transform 1 0 48 0 1 2370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_42
timestamp 1713400504
transform 1 0 48 0 1 2570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_43
timestamp 1713400504
transform 1 0 48 0 1 2770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_44
timestamp 1713400504
transform 1 0 48 0 1 2970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_45
timestamp 1713400504
transform 1 0 3040 0 1 170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_46
timestamp 1713400504
transform 1 0 3040 0 1 370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_47
timestamp 1713400504
transform 1 0 3040 0 1 570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_48
timestamp 1713400504
transform 1 0 3040 0 1 770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_49
timestamp 1713400504
transform 1 0 3040 0 1 970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_50
timestamp 1713400504
transform 1 0 3040 0 1 1170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_51
timestamp 1713400504
transform 1 0 3040 0 1 1370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_52
timestamp 1713400504
transform 1 0 3040 0 1 1570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_53
timestamp 1713400504
transform 1 0 3040 0 1 1770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_54
timestamp 1713400504
transform 1 0 3040 0 1 1970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_55
timestamp 1713400504
transform 1 0 3040 0 1 2170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_56
timestamp 1713400504
transform 1 0 3040 0 1 2370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_57
timestamp 1713400504
transform 1 0 3040 0 1 2570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_58
timestamp 1713400504
transform 1 0 3040 0 1 2770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_59
timestamp 1713400504
transform 1 0 3040 0 1 2970
box -10 -3 10 3
use XNOR2X1  XNOR2X1_0
timestamp 1713400504
transform 1 0 192 0 1 1770
box -8 -3 64 105
use XNOR2X1  XNOR2X1_1
timestamp 1713400504
transform 1 0 152 0 -1 1970
box -8 -3 64 105
use XNOR2X1  XNOR2X1_2
timestamp 1713400504
transform 1 0 216 0 1 2370
box -8 -3 64 105
use XNOR2X1  XNOR2X1_3
timestamp 1713400504
transform 1 0 112 0 1 2570
box -8 -3 64 105
use XNOR2X1  XNOR2X1_4
timestamp 1713400504
transform 1 0 304 0 1 2570
box -8 -3 64 105
use XNOR2X1  XNOR2X1_5
timestamp 1713400504
transform 1 0 352 0 -1 2770
box -8 -3 64 105
use XNOR2X1  XNOR2X1_6
timestamp 1713400504
transform 1 0 512 0 -1 2770
box -8 -3 64 105
use XNOR2X1  XNOR2X1_7
timestamp 1713400504
transform 1 0 576 0 1 2770
box -8 -3 64 105
use XNOR2X1  XNOR2X1_8
timestamp 1713400504
transform 1 0 656 0 -1 2770
box -8 -3 64 105
use XNOR2X1  XNOR2X1_9
timestamp 1713400504
transform 1 0 760 0 -1 2770
box -8 -3 64 105
use XNOR2X1  XNOR2X1_10
timestamp 1713400504
transform 1 0 992 0 1 2570
box -8 -3 64 105
use XNOR2X1  XNOR2X1_11
timestamp 1713400504
transform 1 0 1280 0 1 1970
box -8 -3 64 105
use XNOR2X1  XNOR2X1_12
timestamp 1713400504
transform 1 0 1416 0 1 570
box -8 -3 64 105
use XNOR2X1  XNOR2X1_13
timestamp 1713400504
transform 1 0 1320 0 1 1570
box -8 -3 64 105
use XNOR2X1  XNOR2X1_14
timestamp 1713400504
transform 1 0 1208 0 1 1770
box -8 -3 64 105
use XNOR2X1  XNOR2X1_15
timestamp 1713400504
transform 1 0 1264 0 -1 1370
box -8 -3 64 105
use XNOR2X1  XNOR2X1_16
timestamp 1713400504
transform 1 0 1360 0 -1 1970
box -8 -3 64 105
use XNOR2X1  XNOR2X1_17
timestamp 1713400504
transform 1 0 200 0 -1 170
box -8 -3 64 105
use XNOR2X1  XNOR2X1_18
timestamp 1713400504
transform 1 0 272 0 -1 170
box -8 -3 64 105
use XNOR2X1  XNOR2X1_19
timestamp 1713400504
transform 1 0 392 0 -1 170
box -8 -3 64 105
use XNOR2X1  XNOR2X1_20
timestamp 1713400504
transform 1 0 2264 0 1 1170
box -8 -3 64 105
use XNOR2X1  XNOR2X1_21
timestamp 1713400504
transform 1 0 2144 0 -1 1370
box -8 -3 64 105
use XNOR2X1  XNOR2X1_22
timestamp 1713400504
transform 1 0 2288 0 -1 1170
box -8 -3 64 105
use XNOR2X1  XNOR2X1_23
timestamp 1713400504
transform 1 0 2184 0 1 1370
box -8 -3 64 105
use XNOR2X1  XNOR2X1_24
timestamp 1713400504
transform 1 0 2224 0 -1 1170
box -8 -3 64 105
use XNOR2X1  XNOR2X1_25
timestamp 1713400504
transform 1 0 2344 0 -1 370
box -8 -3 64 105
use XOR2X1  XOR2X1_0
timestamp 1713400504
transform 1 0 888 0 -1 2770
box -8 -3 64 105
use XOR2X1  XOR2X1_1
timestamp 1713400504
transform 1 0 2952 0 -1 970
box -8 -3 64 105
use XOR2X1  XOR2X1_2
timestamp 1713400504
transform 1 0 1264 0 -1 1770
box -8 -3 64 105
use XOR2X1  XOR2X1_3
timestamp 1713400504
transform 1 0 1216 0 1 1370
box -8 -3 64 105
use XOR2X1  XOR2X1_4
timestamp 1713400504
transform 1 0 848 0 -1 2570
box -8 -3 64 105
use XOR2X1  XOR2X1_5
timestamp 1713400504
transform 1 0 792 0 1 2570
box -8 -3 64 105
use XOR2X1  XOR2X1_6
timestamp 1713400504
transform 1 0 680 0 1 2570
box -8 -3 64 105
use XOR2X1  XOR2X1_7
timestamp 1713400504
transform 1 0 568 0 -1 2570
box -8 -3 64 105
use XOR2X1  XOR2X1_8
timestamp 1713400504
transform 1 0 432 0 -1 2570
box -8 -3 64 105
use XOR2X1  XOR2X1_9
timestamp 1713400504
transform 1 0 296 0 -1 1970
box -8 -3 64 105
use XOR2X1  XOR2X1_10
timestamp 1713400504
transform 1 0 1448 0 1 1570
box -8 -3 64 105
use XOR2X1  XOR2X1_11
timestamp 1713400504
transform 1 0 1344 0 -1 1370
box -8 -3 64 105
use XOR2X1  XOR2X1_12
timestamp 1713400504
transform 1 0 1648 0 1 570
box -8 -3 64 105
use XOR2X1  XOR2X1_13
timestamp 1713400504
transform 1 0 2112 0 1 1170
box -8 -3 64 105
use XOR2X1  XOR2X1_14
timestamp 1713400504
transform 1 0 2056 0 1 1170
box -8 -3 64 105
use XOR2X1  XOR2X1_15
timestamp 1713400504
transform 1 0 1992 0 -1 1170
box -8 -3 64 105
use XOR2X1  XOR2X1_16
timestamp 1713400504
transform 1 0 2352 0 -1 970
box -8 -3 64 105
use XOR2X1  XOR2X1_17
timestamp 1713400504
transform 1 0 2264 0 1 970
box -8 -3 64 105
use XOR2X1  XOR2X1_18
timestamp 1713400504
transform 1 0 2224 0 1 770
box -8 -3 64 105
use XOR2X1  XOR2X1_19
timestamp 1713400504
transform 1 0 2176 0 -1 970
box -8 -3 64 105
use XOR2X1  XOR2X1_20
timestamp 1713400504
transform 1 0 1960 0 -1 970
box -8 -3 64 105
use XOR2X1  XOR2X1_21
timestamp 1713400504
transform 1 0 2320 0 1 1170
box -8 -3 64 105
use XOR2X1  XOR2X1_22
timestamp 1713400504
transform 1 0 2232 0 -1 1370
box -8 -3 64 105
use XOR2X1  XOR2X1_23
timestamp 1713400504
transform 1 0 2112 0 1 1370
box -8 -3 64 105
use XOR2X1  XOR2X1_24
timestamp 1713400504
transform 1 0 2016 0 -1 1370
box -8 -3 64 105
use XOR2X1  XOR2X1_25
timestamp 1713400504
transform 1 0 2088 0 1 970
box -8 -3 64 105
use XOR2X1  XOR2X1_26
timestamp 1713400504
transform 1 0 2048 0 -1 1170
box -8 -3 64 105
use XOR2X1  XOR2X1_27
timestamp 1713400504
transform 1 0 1952 0 1 970
box -8 -3 64 105
<< labels >>
rlabel metal3 3085 1455 3085 1455 4 in_clka
rlabel metal2 1580 1 1580 1 4 in_clkb
rlabel metal3 3085 725 3085 725 4 in_restart
rlabel metal3 2 2135 2 2135 4 in_mult[2]
rlabel metal3 2 2115 2 2115 4 in_mult[1]
rlabel metal3 2 2005 2 2005 4 in_mult[0]
rlabel metal3 2 2415 2 2415 4 in_incr[2]
rlabel metal3 2 2215 2 2215 4 in_incr[1]
rlabel metal3 2 1965 2 1965 4 in_incr[0]
rlabel metal2 444 1 444 1 4 in_n_mines[2]
rlabel metal2 252 1 252 1 4 in_n_mines[1]
rlabel metal2 324 1 324 1 4 in_n_mines[0]
rlabel metal2 2756 1 2756 1 4 out_state_main[3]
rlabel metal2 2804 1 2804 1 4 out_state_main[2]
rlabel metal2 2772 1 2772 1 4 out_state_main[1]
rlabel metal2 2788 1 2788 1 4 out_state_main[0]
rlabel metal2 2852 1 2852 1 4 in_place
rlabel metal3 3085 485 3085 485 4 in_data_in
rlabel metal2 1876 1 1876 1 4 in_data[4]
rlabel metal2 1828 1 1828 1 4 in_data[3]
rlabel metal2 1724 1 1724 1 4 in_data[2]
rlabel metal2 1756 1 1756 1 4 in_data[1]
rlabel metal2 1796 1 1796 1 4 in_data[0]
rlabel metal2 1812 1 1812 1 4 out_start
rlabel metal2 2084 1 2084 1 4 out_place_done
rlabel metal3 2 1645 2 1645 4 out_mines[24]
rlabel metal3 2 1285 2 1285 4 out_mines[23]
rlabel metal3 2 1325 2 1325 4 out_mines[22]
rlabel metal3 2 1515 2 1515 4 out_mines[21]
rlabel metal3 2 1415 2 1415 4 out_mines[20]
rlabel metal3 2 1345 2 1345 4 out_mines[19]
rlabel metal3 2 1445 2 1445 4 out_mines[18]
rlabel metal3 2 1695 2 1695 4 out_mines[17]
rlabel metal3 2 1855 2 1855 4 out_mines[16]
rlabel metal3 2 1545 2 1545 4 out_mines[15]
rlabel metal3 2 1495 2 1495 4 out_mines[14]
rlabel metal2 1276 3038 1276 3038 4 out_mines[13]
rlabel metal3 2 1585 2 1585 4 out_mines[12]
rlabel metal2 1532 1 1532 1 4 out_mines[11]
rlabel metal2 1564 1 1564 1 4 out_mines[10]
rlabel metal3 2 1365 2 1365 4 out_mines[9]
rlabel metal3 2 1475 2 1475 4 out_mines[8]
rlabel metal2 1484 3038 1484 3038 4 out_mines[7]
rlabel metal3 2 1395 2 1395 4 out_mines[6]
rlabel metal3 2 1305 2 1305 4 out_mines[5]
rlabel metal2 1268 1 1268 1 4 out_mines[4]
rlabel metal2 1468 1 1468 1 4 out_mines[3]
rlabel metal2 1596 1 1596 1 4 out_mines[2]
rlabel metal3 2 1255 2 1255 4 out_mines[1]
rlabel metal3 2 1235 2 1235 4 out_mines[0]
rlabel metal2 1980 1 1980 1 4 out_load
rlabel metal2 1740 1 1740 1 4 out_temp_data_in[4]
rlabel metal2 1652 1 1652 1 4 out_temp_data_in[3]
rlabel metal2 1620 1 1620 1 4 out_temp_data_in[2]
rlabel metal2 1484 1 1484 1 4 out_temp_data_in[1]
rlabel metal3 2 1565 2 1565 4 out_temp_data_in[0]
rlabel metal2 2228 1 2228 1 4 out_decode
rlabel metal2 2100 1 2100 1 4 out_alu
rlabel metal3 3085 655 3085 655 4 out_alu_done
rlabel metal3 3085 905 3085 905 4 out_gameover
rlabel metal3 3085 1365 3085 1365 4 out_win
rlabel metal3 3085 955 3085 955 4 out_global_score[7]
rlabel metal3 3085 785 3085 785 4 out_global_score[6]
rlabel metal3 3085 815 3085 815 4 out_global_score[5]
rlabel metal3 3085 1015 3085 1015 4 out_global_score[4]
rlabel metal3 3085 1125 3085 1125 4 out_global_score[3]
rlabel metal3 3085 1215 3085 1215 4 out_global_score[2]
rlabel metal3 3085 1325 3085 1325 4 out_global_score[1]
rlabel metal3 3085 1385 3085 1385 4 out_global_score[0]
rlabel metal3 3085 925 3085 925 4 out_n_nearby[1]
rlabel metal3 3085 975 3085 975 4 out_n_nearby[0]
rlabel metal3 3085 1905 3085 1905 4 out_temp_decoded[24]
rlabel metal2 1932 3038 1932 3038 4 out_temp_decoded[23]
rlabel metal2 1764 3038 1764 3038 4 out_temp_decoded[22]
rlabel metal2 1796 3038 1796 3038 4 out_temp_decoded[21]
rlabel metal2 1868 3038 1868 3038 4 out_temp_decoded[20]
rlabel metal2 1452 3038 1452 3038 4 out_temp_decoded[19]
rlabel metal2 1436 3038 1436 3038 4 out_temp_decoded[18]
rlabel metal2 1580 3038 1580 3038 4 out_temp_decoded[17]
rlabel metal2 1420 3038 1420 3038 4 out_temp_decoded[16]
rlabel metal2 1508 3038 1508 3038 4 out_temp_decoded[15]
rlabel metal2 1964 3038 1964 3038 4 out_temp_decoded[14]
rlabel metal2 1916 3038 1916 3038 4 out_temp_decoded[13]
rlabel metal2 2076 3038 2076 3038 4 out_temp_decoded[12]
rlabel metal2 2404 3038 2404 3038 4 out_temp_decoded[11]
rlabel metal2 2476 3038 2476 3038 4 out_temp_decoded[10]
rlabel metal2 2260 3038 2260 3038 4 out_temp_decoded[9]
rlabel metal3 3085 2725 3085 2725 4 out_temp_decoded[8]
rlabel metal3 3085 2415 3085 2415 4 out_temp_decoded[7]
rlabel metal3 3085 2245 3085 2245 4 out_temp_decoded[6]
rlabel metal3 3085 2125 3085 2125 4 out_temp_decoded[5]
rlabel metal3 3085 1725 3085 1725 4 out_temp_decoded[4]
rlabel metal3 3085 1745 3085 1745 4 out_temp_decoded[3]
rlabel metal3 3085 2085 3085 2085 4 out_temp_decoded[2]
rlabel metal3 3085 1945 3085 1945 4 out_temp_decoded[1]
rlabel metal3 3085 1575 3085 1575 4 out_temp_decoded[0]
rlabel metal3 3085 1925 3085 1925 4 out_temp_cleared[24]
rlabel metal2 1948 3038 1948 3038 4 out_temp_cleared[23]
rlabel metal2 1620 3038 1620 3038 4 out_temp_cleared[22]
rlabel metal2 1468 3038 1468 3038 4 out_temp_cleared[21]
rlabel metal2 1596 3038 1596 3038 4 out_temp_cleared[20]
rlabel metal2 1388 3038 1388 3038 4 out_temp_cleared[19]
rlabel metal2 1308 3038 1308 3038 4 out_temp_cleared[18]
rlabel metal2 1148 3038 1148 3038 4 out_temp_cleared[17]
rlabel metal2 1132 3038 1132 3038 4 out_temp_cleared[16]
rlabel metal2 1164 3038 1164 3038 4 out_temp_cleared[15]
rlabel metal2 1780 3038 1780 3038 4 out_temp_cleared[14]
rlabel metal2 1852 3038 1852 3038 4 out_temp_cleared[13]
rlabel metal2 1996 3038 1996 3038 4 out_temp_cleared[12]
rlabel metal2 2564 3038 2564 3038 4 out_temp_cleared[11]
rlabel metal2 2620 3038 2620 3038 4 out_temp_cleared[10]
rlabel metal2 2844 3038 2844 3038 4 out_temp_cleared[9]
rlabel metal3 3085 2775 3085 2775 4 out_temp_cleared[8]
rlabel metal3 3085 2605 3085 2605 4 out_temp_cleared[7]
rlabel metal3 3085 2325 3085 2325 4 out_temp_cleared[6]
rlabel metal3 3085 2015 3085 2015 4 out_temp_cleared[5]
rlabel metal3 3085 1525 3085 1525 4 out_temp_cleared[4]
rlabel metal3 3085 1545 3085 1545 4 out_temp_cleared[3]
rlabel metal3 3085 2305 3085 2305 4 out_temp_cleared[2]
rlabel metal3 3085 1765 3085 1765 4 out_temp_cleared[1]
rlabel metal3 3085 1675 3085 1675 4 out_temp_cleared[0]
rlabel metal2 2356 1 2356 1 4 out_display
rlabel metal3 3085 635 3085 635 4 out_display_done
rlabel metal3 2 1765 2 1765 4 out_temp_index[4]
rlabel metal3 2 1675 2 1675 4 out_temp_index[3]
rlabel metal3 2 1605 2 1605 4 out_temp_index[2]
rlabel metal3 2 1745 2 1745 4 out_temp_index[1]
rlabel metal3 2 1715 2 1715 4 out_temp_index[0]
rlabel metal2 428 1 428 1 4 out_temp_mine_cnt[2]
rlabel metal2 188 1 188 1 4 out_temp_mine_cnt[1]
rlabel metal3 2 325 2 325 4 out_temp_mine_cnt[0]
rlabel metal2 38 37 38 37 4 gnd
rlabel metal2 14 13 14 13 4 vdd
<< properties >>
string path 25884.002 10935.000 25884.002 11025.000 
<< end >>
