* SPICE3 file created from top_module.ext - technology: scmos

.option scale=0.3u

M1000 DFFNEGX1_51/a_76_6# BUFX2_14/Y DFFNEGX1_51/a_66_6# Gnd nfet w=10 l=2
+  ad=14.999999p pd=13u as=40p ps=18u
M1001 gnd BUFX2_14/Y DFFNEGX1_51/a_2_6# Gnd nfet w=20 l=2
+  ad=55p pd=26u as=100p ps=50u
M1002 DFFNEGX1_51/a_66_6# DFFNEGX1_51/a_2_6# DFFNEGX1_51/a_61_6# Gnd nfet w=10 l=2
+  ad=40p pd=18u as=14.999999p ps=13u
M1003 out_temp_decoded[15] DFFNEGX1_51/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=55p ps=26u
M1004 DFFNEGX1_51/a_23_6# BUFX2_14/Y DFFNEGX1_51/a_17_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=16u as=20p ps=14u
M1005 DFFNEGX1_51/a_23_6# DFFNEGX1_51/a_2_6# DFFNEGX1_51/a_17_74# vdd pfet w=20 l=2
+  ad=59.999996p pd=26u as=40p ps=24u
M1006 gnd DFFNEGX1_51/a_34_4# DFFNEGX1_51/a_31_6# Gnd nfet w=10 l=2
+  ad=35p pd=17u as=14.999999p ps=13u
M1007 vdd DFFNEGX1_51/a_34_4# DFFNEGX1_51/a_31_74# vdd pfet w=20 l=2
+  ad=59.999996p pd=26u as=40p ps=24u
M1008 DFFNEGX1_51/a_61_74# DFFNEGX1_51/a_34_4# vdd vdd pfet w=20 l=2
+  ad=29.999998p pd=23u as=100p ps=50u
M1009 DFFNEGX1_51/a_34_4# DFFNEGX1_51/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=59.999996p ps=26u
M1010 DFFNEGX1_51/a_34_4# DFFNEGX1_51/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=35p ps=17u
M1011 vdd out_temp_decoded[15] DFFNEGX1_51/a_76_84# vdd pfet w=10 l=2
+  ad=0.105n pd=46u as=14.999999p ps=13u
M1012 gnd out_temp_decoded[15] DFFNEGX1_51/a_76_6# Gnd nfet w=10 l=2
+  ad=55p pd=26u as=14.999999p ps=13u
M1013 DFFNEGX1_51/a_61_6# DFFNEGX1_51/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=14.999999p pd=13u as=50p ps=30u
M1014 DFFNEGX1_51/a_76_84# DFFNEGX1_51/a_2_6# DFFNEGX1_51/a_66_6# vdd pfet w=10 l=2
+  ad=14.999999p pd=13u as=75p ps=28u
M1015 out_temp_decoded[15] DFFNEGX1_51/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.105n ps=46u
M1016 vdd BUFX2_14/Y DFFNEGX1_51/a_2_6# vdd pfet w=40 l=2
+  ad=0.11n pd=46u as=0.2n ps=90u
M1017 DFFNEGX1_51/a_31_6# DFFNEGX1_51/a_2_6# DFFNEGX1_51/a_23_6# Gnd nfet w=10 l=2
+  ad=14.999999p pd=13u as=29.999998p ps=16u
M1018 DFFNEGX1_51/a_66_6# BUFX2_14/Y DFFNEGX1_51/a_61_74# vdd pfet w=20 l=2
+  ad=75p pd=28u as=29.999998p ps=23u
M1019 DFFNEGX1_51/a_17_74# OAI21X1_97/Y vdd vdd pfet w=20 l=2
+  ad=40p pd=24u as=0.11n ps=46u
M1020 DFFNEGX1_51/a_31_74# BUFX2_14/Y DFFNEGX1_51/a_23_6# vdd pfet w=20 l=2
+  ad=40p pd=24u as=59.999996p ps=26u
M1021 DFFNEGX1_51/a_17_6# OAI21X1_97/Y gnd Gnd nfet w=10 l=2
+  ad=20p pd=14u as=55p ps=26u
M1022 DFFNEGX1_40/a_76_6# BUFX2_15/Y DFFNEGX1_40/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1023 gnd BUFX2_15/Y DFFNEGX1_40/a_2_6# Gnd nfet w=20 l=2
+  ad=0.21371u pd=0.103284 as=100p ps=50u
M1024 DFFNEGX1_40/a_66_6# DFFNEGX1_40/a_2_6# DFFNEGX1_40/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1025 out_temp_data_in[1] DFFNEGX1_40/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1026 DFFNEGX1_40/a_23_6# BUFX2_15/Y DFFNEGX1_40/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1027 DFFNEGX1_40/a_23_6# DFFNEGX1_40/a_2_6# DFFNEGX1_40/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1028 gnd DFFNEGX1_40/a_34_4# DFFNEGX1_40/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1029 vdd DFFNEGX1_40/a_34_4# DFFNEGX1_40/a_31_74# vdd pfet w=20 l=2
+  ad=0.431054u pd=0.188526 as=80p ps=48u
M1030 DFFNEGX1_40/a_61_74# DFFNEGX1_40/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1031 DFFNEGX1_40/a_34_4# DFFNEGX1_40/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1032 DFFNEGX1_40/a_34_4# DFFNEGX1_40/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1033 vdd out_temp_data_in[1] DFFNEGX1_40/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1034 gnd out_temp_data_in[1] DFFNEGX1_40/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1035 DFFNEGX1_40/a_61_6# DFFNEGX1_40/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1036 DFFNEGX1_40/a_76_84# DFFNEGX1_40/a_2_6# DFFNEGX1_40/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1037 out_temp_data_in[1] DFFNEGX1_40/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1038 vdd BUFX2_15/Y DFFNEGX1_40/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1039 DFFNEGX1_40/a_31_6# DFFNEGX1_40/a_2_6# DFFNEGX1_40/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1040 DFFNEGX1_40/a_66_6# BUFX2_15/Y DFFNEGX1_40/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1041 DFFNEGX1_40/a_17_74# OAI21X1_108/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1042 DFFNEGX1_40/a_31_74# BUFX2_15/Y DFFNEGX1_40/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1043 DFFNEGX1_40/a_17_6# OAI21X1_108/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1044 DFFNEGX1_95/a_76_6# BUFX2_10/Y DFFNEGX1_95/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1045 gnd BUFX2_10/Y DFFNEGX1_95/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1046 DFFNEGX1_95/a_66_6# DFFNEGX1_95/a_2_6# DFFNEGX1_95/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1047 out_global_score[1] DFFNEGX1_95/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1048 DFFNEGX1_95/a_23_6# BUFX2_10/Y DFFNEGX1_95/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1049 DFFNEGX1_95/a_23_6# DFFNEGX1_95/a_2_6# DFFNEGX1_95/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1050 gnd DFFNEGX1_95/a_34_4# DFFNEGX1_95/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1051 vdd DFFNEGX1_95/a_34_4# DFFNEGX1_95/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1052 DFFNEGX1_95/a_61_74# DFFNEGX1_95/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1053 DFFNEGX1_95/a_34_4# DFFNEGX1_95/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1054 DFFNEGX1_95/a_34_4# DFFNEGX1_95/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1055 vdd out_global_score[1] DFFNEGX1_95/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1056 gnd out_global_score[1] DFFNEGX1_95/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1057 DFFNEGX1_95/a_61_6# DFFNEGX1_95/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1058 DFFNEGX1_95/a_76_84# DFFNEGX1_95/a_2_6# DFFNEGX1_95/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1059 out_global_score[1] DFFNEGX1_95/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1060 vdd BUFX2_10/Y DFFNEGX1_95/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1061 DFFNEGX1_95/a_31_6# DFFNEGX1_95/a_2_6# DFFNEGX1_95/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1062 DFFNEGX1_95/a_66_6# BUFX2_10/Y DFFNEGX1_95/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1063 DFFNEGX1_95/a_17_74# INVX2_215/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1064 DFFNEGX1_95/a_31_74# BUFX2_10/Y DFFNEGX1_95/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1065 DFFNEGX1_95/a_17_6# INVX2_215/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1066 DFFNEGX1_84/a_76_6# BUFX2_11/Y DFFNEGX1_84/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1067 gnd BUFX2_11/Y DFFNEGX1_84/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1068 DFFNEGX1_84/a_66_6# DFFNEGX1_84/a_2_6# DFFNEGX1_84/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1069 out_temp_cleared[7] DFFNEGX1_84/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1070 DFFNEGX1_84/a_23_6# BUFX2_11/Y DFFNEGX1_84/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1071 DFFNEGX1_84/a_23_6# DFFNEGX1_84/a_2_6# DFFNEGX1_84/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1072 gnd DFFNEGX1_84/a_34_4# DFFNEGX1_84/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1073 vdd DFFNEGX1_84/a_34_4# DFFNEGX1_84/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1074 DFFNEGX1_84/a_61_74# DFFNEGX1_84/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1075 DFFNEGX1_84/a_34_4# DFFNEGX1_84/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1076 DFFNEGX1_84/a_34_4# DFFNEGX1_84/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1077 vdd out_temp_cleared[7] DFFNEGX1_84/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1078 gnd out_temp_cleared[7] DFFNEGX1_84/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1079 DFFNEGX1_84/a_61_6# DFFNEGX1_84/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1080 DFFNEGX1_84/a_76_84# DFFNEGX1_84/a_2_6# DFFNEGX1_84/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1081 out_temp_cleared[7] DFFNEGX1_84/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1082 vdd BUFX2_11/Y DFFNEGX1_84/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1083 DFFNEGX1_84/a_31_6# DFFNEGX1_84/a_2_6# DFFNEGX1_84/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1084 DFFNEGX1_84/a_66_6# BUFX2_11/Y DFFNEGX1_84/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1085 DFFNEGX1_84/a_17_74# OAI22X1_21/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1086 DFFNEGX1_84/a_31_74# BUFX2_11/Y DFFNEGX1_84/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1087 DFFNEGX1_84/a_17_6# OAI22X1_21/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1088 DFFNEGX1_73/a_76_6# BUFX2_12/Y DFFNEGX1_73/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1089 gnd BUFX2_12/Y DFFNEGX1_73/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1090 DFFNEGX1_73/a_66_6# DFFNEGX1_73/a_2_6# DFFNEGX1_73/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1091 out_temp_cleared[18] DFFNEGX1_73/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1092 DFFNEGX1_73/a_23_6# BUFX2_12/Y DFFNEGX1_73/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1093 DFFNEGX1_73/a_23_6# DFFNEGX1_73/a_2_6# DFFNEGX1_73/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1094 gnd DFFNEGX1_73/a_34_4# DFFNEGX1_73/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1095 vdd DFFNEGX1_73/a_34_4# DFFNEGX1_73/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1096 DFFNEGX1_73/a_61_74# DFFNEGX1_73/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1097 DFFNEGX1_73/a_34_4# DFFNEGX1_73/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1098 DFFNEGX1_73/a_34_4# DFFNEGX1_73/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1099 vdd out_temp_cleared[18] DFFNEGX1_73/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1100 gnd out_temp_cleared[18] DFFNEGX1_73/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1101 DFFNEGX1_73/a_61_6# DFFNEGX1_73/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1102 DFFNEGX1_73/a_76_84# DFFNEGX1_73/a_2_6# DFFNEGX1_73/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1103 out_temp_cleared[18] DFFNEGX1_73/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1104 vdd BUFX2_12/Y DFFNEGX1_73/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1105 DFFNEGX1_73/a_31_6# DFFNEGX1_73/a_2_6# DFFNEGX1_73/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1106 DFFNEGX1_73/a_66_6# BUFX2_12/Y DFFNEGX1_73/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1107 DFFNEGX1_73/a_17_74# OAI22X1_10/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1108 DFFNEGX1_73/a_31_74# BUFX2_12/Y DFFNEGX1_73/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1109 DFFNEGX1_73/a_17_6# OAI22X1_10/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1110 DFFNEGX1_62/a_76_6# BUFX2_13/Y DFFNEGX1_62/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1111 gnd BUFX2_13/Y DFFNEGX1_62/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1112 DFFNEGX1_62/a_66_6# DFFNEGX1_62/a_2_6# DFFNEGX1_62/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1113 out_temp_decoded[4] DFFNEGX1_62/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1114 DFFNEGX1_62/a_23_6# BUFX2_13/Y DFFNEGX1_62/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1115 DFFNEGX1_62/a_23_6# DFFNEGX1_62/a_2_6# DFFNEGX1_62/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1116 gnd DFFNEGX1_62/a_34_4# DFFNEGX1_62/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1117 vdd DFFNEGX1_62/a_34_4# DFFNEGX1_62/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1118 DFFNEGX1_62/a_61_74# DFFNEGX1_62/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1119 DFFNEGX1_62/a_34_4# DFFNEGX1_62/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1120 DFFNEGX1_62/a_34_4# DFFNEGX1_62/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1121 vdd out_temp_decoded[4] DFFNEGX1_62/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1122 gnd out_temp_decoded[4] DFFNEGX1_62/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1123 DFFNEGX1_62/a_61_6# DFFNEGX1_62/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1124 DFFNEGX1_62/a_76_84# DFFNEGX1_62/a_2_6# DFFNEGX1_62/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1125 out_temp_decoded[4] DFFNEGX1_62/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1126 vdd BUFX2_13/Y DFFNEGX1_62/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1127 DFFNEGX1_62/a_31_6# DFFNEGX1_62/a_2_6# DFFNEGX1_62/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1128 DFFNEGX1_62/a_66_6# BUFX2_13/Y DFFNEGX1_62/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1129 DFFNEGX1_62/a_17_74# OAI21X1_86/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1130 DFFNEGX1_62/a_31_74# BUFX2_13/Y DFFNEGX1_62/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1131 DFFNEGX1_62/a_17_6# OAI21X1_86/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1132 vdd out_global_score[21] HAX1_9/a_2_74# vdd pfet w=20 l=2
+  ad=59.999996p pd=26u as=100p ps=50u
M1133 HAX1_9/a_41_74# HAX1_9/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.11n pd=46u as=59.999996p ps=26u
M1134 HAX1_9/a_9_6# out_global_score[21] gnd Gnd nfet w=20 l=2
+  ad=29.999998p pd=23u as=100p ps=50u
M1135 HAX1_9/a_41_74# HAX1_9/B HAX1_9/a_38_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=26u as=59.999996p ps=26u
M1136 vdd out_global_score[21] HAX1_9/a_49_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=59.999996p ps=43u
M1137 vdd HAX1_9/a_2_74# HAX1_8/B vdd pfet w=20 l=2
+  ad=59.999996p pd=26u as=100p ps=50u
M1138 HAX1_9/a_38_6# HAX1_9/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=26u as=54p ps=26u
M1139 HAX1_9/YS HAX1_9/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1140 HAX1_9/a_38_6# out_global_score[21] HAX1_9/a_41_74# Gnd nfet w=20 l=2
+  ad=96p pd=50u as=59.999996p ps=26u
M1141 HAX1_9/YS HAX1_9/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M1142 HAX1_9/a_2_74# HAX1_9/B vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=59.999996p ps=26u
M1143 HAX1_9/a_2_74# HAX1_9/B HAX1_9/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=29.999998p ps=23u
M1144 HAX1_9/a_49_54# HAX1_9/B HAX1_9/a_41_74# vdd pfet w=40 l=2
+  ad=59.999996p pd=43u as=0.11n ps=46u
M1145 gnd HAX1_9/a_2_74# HAX1_8/B Gnd nfet w=10 l=2
+  ad=54p pd=26u as=50p ps=30u
M1146 AND2X2_5/a_2_6# out_temp_data_in[1] vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=26u as=100p ps=50u
M1147 AND2X2_5/a_9_6# out_temp_data_in[1] AND2X2_5/a_2_6# Gnd nfet w=20 l=2
+  ad=29.999998p pd=23u as=100p ps=50u
M1148 OR2X1_10/B AND2X2_5/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=59.999996p ps=26u
M1149 OR2X1_10/B AND2X2_5/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.108n ps=46u
M1150 vdd out_temp_data_in[2] AND2X2_5/a_2_6# vdd pfet w=20 l=2
+  ad=0.108n pd=46u as=59.999996p ps=26u
M1151 gnd out_temp_data_in[2] AND2X2_5/a_9_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=26u as=29.999998p ps=23u
M1152 gnd XNOR2X1_7/Y MUX2X1_17/a_30_10# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=29.999998p ps=23u
M1153 MUX2X1_17/a_17_50# MUX2X1_17/B vdd vdd pfet w=40 l=2
+  ad=59.999996p pd=43u as=0.104n ps=46u
M1154 MUX2X1_17/Y OR2X1_3/Y MUX2X1_17/a_17_50# vdd pfet w=40 l=2
+  ad=0.124n pd=50u as=59.999996p ps=43u
M1155 MUX2X1_17/a_30_54# MUX2X1_17/a_2_10# MUX2X1_17/Y vdd pfet w=40 l=2
+  ad=59.999996p pd=43u as=0.124n ps=50u
M1156 MUX2X1_17/a_17_10# MUX2X1_17/B gnd Gnd nfet w=20 l=2
+  ad=29.999998p pd=23u as=53p ps=26u
M1157 vdd OR2X1_3/Y MUX2X1_17/a_2_10# vdd pfet w=20 l=2
+  ad=0.104n pd=46u as=100p ps=50u
M1158 MUX2X1_17/a_30_10# OR2X1_3/Y MUX2X1_17/Y Gnd nfet w=20 l=2
+  ad=29.999998p pd=23u as=59.999996p ps=26u
M1159 gnd OR2X1_3/Y MUX2X1_17/a_2_10# Gnd nfet w=10 l=2
+  ad=53p pd=26u as=50p ps=30u
M1160 vdd XNOR2X1_7/Y MUX2X1_17/a_30_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=59.999996p ps=43u
M1161 MUX2X1_17/Y MUX2X1_17/a_2_10# MUX2X1_17/a_17_10# Gnd nfet w=20 l=2
+  ad=59.999996p pd=26u as=29.999998p ps=23u
M1162 DFFNEGX1_141/a_76_6# INVX2_259/Y DFFNEGX1_141/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1163 gnd INVX2_259/Y DFFNEGX1_141/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1164 DFFNEGX1_141/a_66_6# DFFNEGX1_141/a_2_6# DFFNEGX1_141/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1165 out_alu DFFNEGX1_141/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1166 DFFNEGX1_141/a_23_6# INVX2_259/Y DFFNEGX1_141/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1167 DFFNEGX1_141/a_23_6# DFFNEGX1_141/a_2_6# DFFNEGX1_141/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1168 gnd DFFNEGX1_141/a_34_4# DFFNEGX1_141/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1169 vdd DFFNEGX1_141/a_34_4# DFFNEGX1_141/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1170 DFFNEGX1_141/a_61_74# DFFNEGX1_141/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1171 DFFNEGX1_141/a_34_4# DFFNEGX1_141/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1172 DFFNEGX1_141/a_34_4# DFFNEGX1_141/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1173 vdd out_alu DFFNEGX1_141/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1174 gnd out_alu DFFNEGX1_141/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1175 DFFNEGX1_141/a_61_6# DFFNEGX1_141/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1176 DFFNEGX1_141/a_76_84# DFFNEGX1_141/a_2_6# DFFNEGX1_141/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1177 out_alu DFFNEGX1_141/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1178 vdd INVX2_259/Y DFFNEGX1_141/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1179 DFFNEGX1_141/a_31_6# DFFNEGX1_141/a_2_6# DFFNEGX1_141/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1180 DFFNEGX1_141/a_66_6# INVX2_259/Y DFFNEGX1_141/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1181 DFFNEGX1_141/a_17_74# OAI21X1_157/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1182 DFFNEGX1_141/a_31_74# INVX2_259/Y DFFNEGX1_141/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1183 DFFNEGX1_141/a_17_6# OAI21X1_157/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1184 DFFNEGX1_130/a_76_6# INVX2_259/Y DFFNEGX1_130/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1185 gnd INVX2_259/Y DFFNEGX1_130/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1186 DFFNEGX1_130/a_66_6# DFFNEGX1_130/a_2_6# DFFNEGX1_130/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1187 out_state_main[0] DFFNEGX1_130/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1188 DFFNEGX1_130/a_23_6# INVX2_259/Y DFFNEGX1_130/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1189 DFFNEGX1_130/a_23_6# DFFNEGX1_130/a_2_6# DFFNEGX1_130/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1190 gnd DFFNEGX1_130/a_34_4# DFFNEGX1_130/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1191 vdd DFFNEGX1_130/a_34_4# DFFNEGX1_130/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1192 DFFNEGX1_130/a_61_74# DFFNEGX1_130/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1193 DFFNEGX1_130/a_34_4# DFFNEGX1_130/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1194 DFFNEGX1_130/a_34_4# DFFNEGX1_130/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1195 vdd out_state_main[0] DFFNEGX1_130/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1196 gnd out_state_main[0] DFFNEGX1_130/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1197 DFFNEGX1_130/a_61_6# DFFNEGX1_130/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1198 DFFNEGX1_130/a_76_84# DFFNEGX1_130/a_2_6# DFFNEGX1_130/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1199 out_state_main[0] DFFNEGX1_130/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1200 vdd INVX2_259/Y DFFNEGX1_130/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1201 DFFNEGX1_130/a_31_6# DFFNEGX1_130/a_2_6# DFFNEGX1_130/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1202 DFFNEGX1_130/a_66_6# INVX2_259/Y DFFNEGX1_130/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1203 DFFNEGX1_130/a_17_74# INVX2_127/A vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1204 DFFNEGX1_130/a_31_74# INVX2_259/Y DFFNEGX1_130/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1205 DFFNEGX1_130/a_17_6# INVX2_127/A gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1206 gnd XNOR2X1_2/Y MUX2X1_28/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M1207 MUX2X1_28/a_17_50# NOR2X1_1/A vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1208 XNOR2X1_1/A OR2X1_1/Y MUX2X1_28/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M1209 MUX2X1_28/a_30_54# MUX2X1_28/a_2_10# XNOR2X1_1/A vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1210 MUX2X1_28/a_17_10# NOR2X1_1/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1211 vdd OR2X1_1/Y MUX2X1_28/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1212 MUX2X1_28/a_30_10# OR2X1_1/Y XNOR2X1_1/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M1213 gnd OR2X1_1/Y MUX2X1_28/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M1214 vdd XNOR2X1_2/Y MUX2X1_28/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1215 XNOR2X1_1/A MUX2X1_28/a_2_10# MUX2X1_28/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1216 gnd INVX2_86/Y AOI22X1_0/a_28_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=29.999998p ps=23u
M1217 AOI22X1_0/Y XOR2X1_24/Y AOI22X1_0/a_11_6# Gnd nfet w=20 l=2
+  ad=100p pd=30u as=29.999998p ps=23u
M1218 AOI22X1_0/a_11_6# OR2X1_14/B gnd Gnd nfet w=20 l=2
+  ad=29.999998p pd=23u as=100p ps=50u
M1219 AOI22X1_0/a_2_54# XOR2X1_24/Y vdd vdd pfet w=40 l=2
+  ad=0.12n pd=46u as=0.12n ps=46u
M1220 AOI22X1_0/a_28_6# XOR2X1_16/Y AOI22X1_0/Y Gnd nfet w=20 l=2
+  ad=29.999998p pd=23u as=100p ps=30u
M1221 vdd OR2X1_14/B AOI22X1_0/a_2_54# vdd pfet w=40 l=2
+  ad=0.12n pd=46u as=0.2n ps=90u
M1222 AOI22X1_0/Y XOR2X1_16/Y AOI22X1_0/a_2_54# vdd pfet w=40 l=2
+  ad=0.12n pd=46u as=0.12n ps=46u
M1223 AOI22X1_0/a_2_54# INVX2_86/Y AOI22X1_0/Y vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=46u
M1224 OAI21X1_6/A NOR2X1_65/A vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=26u as=100p ps=50u
M1225 NAND2X1_21/a_9_6# NOR2X1_65/A gnd Gnd nfet w=20 l=2
+  ad=29.999998p pd=23u as=100p ps=50u
M1226 vdd NOR2X1_61/Y OAI21X1_6/A vdd pfet w=20 l=2
+  ad=100p pd=50u as=59.999996p ps=26u
M1227 OAI21X1_6/A NOR2X1_61/Y NAND2X1_21/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=29.999998p ps=23u
M1228 OAI21X1_46/B NOR2X1_64/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1229 NAND2X1_43/a_9_6# NOR2X1_64/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1230 vdd NOR2X1_65/A OAI21X1_46/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1231 OAI21X1_46/B NOR2X1_65/A NAND2X1_43/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1232 OAI21X1_31/C out_mines[10] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1233 NAND2X1_32/a_9_6# out_mines[10] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1234 vdd INVX2_242/Y OAI21X1_31/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1235 OAI21X1_31/C INVX2_242/Y NAND2X1_32/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1236 NOR2X1_43/A out_temp_data_in[3] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1237 NAND2X1_10/a_9_6# out_temp_data_in[3] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1238 vdd OAI21X1_1/B NOR2X1_43/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1239 NOR2X1_43/A OAI21X1_1/B NAND2X1_10/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1240 OAI21X1_89/C NOR2X1_37/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1241 NAND2X1_76/a_9_6# NOR2X1_37/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1242 vdd BUFX2_20/Y OAI21X1_89/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1243 OAI21X1_89/C BUFX2_20/Y NAND2X1_76/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1244 OAI21X1_76/B INVX2_111/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1245 NAND2X1_65/a_9_6# INVX2_111/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1246 vdd INVX2_82/Y OAI21X1_76/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1247 OAI21X1_76/B INVX2_82/Y NAND2X1_65/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1248 OAI21X1_58/C out_alu_done vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1249 NAND2X1_54/a_9_6# out_alu_done gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1250 vdd INVX2_184/Y OAI21X1_58/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1251 OAI21X1_58/C INVX2_184/Y NAND2X1_54/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1252 NAND2X1_87/Y NOR2X1_50/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1253 NAND2X1_87/a_9_6# NOR2X1_50/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1254 vdd BUFX2_21/Y NAND2X1_87/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1255 NAND2X1_87/Y BUFX2_21/Y NAND2X1_87/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1256 NAND2X1_98/Y in_data[2] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1257 NAND2X1_98/a_9_6# in_data[2] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1258 vdd NOR2X1_107/Y NAND2X1_98/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1259 NAND2X1_98/Y NOR2X1_107/Y NAND2X1_98/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1260 gnd out_global_score[3] AOI22X1_30/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M1261 INVX2_213/A INVX2_258/Y AOI22X1_30/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M1262 AOI22X1_30/a_11_6# HAX1_27/YS gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1263 AOI22X1_30/a_2_54# INVX2_258/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M1264 AOI22X1_30/a_28_6# INVX2_255/Y INVX2_213/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1265 vdd HAX1_27/YS AOI22X1_30/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1266 INVX2_213/A INVX2_255/Y AOI22X1_30/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M1267 AOI22X1_30/a_2_54# out_global_score[3] INVX2_213/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1268 gnd out_temp_decoded[13] AOI22X1_41/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M1269 OAI21X1_73/C out_mines[12] AOI22X1_41/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M1270 AOI22X1_41/a_11_6# out_temp_decoded[12] gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1271 AOI22X1_41/a_2_54# out_mines[12] vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M1272 AOI22X1_41/a_28_6# out_mines[13] OAI21X1_73/C Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1273 vdd out_temp_decoded[12] AOI22X1_41/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1274 OAI21X1_73/C out_mines[13] AOI22X1_41/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M1275 AOI22X1_41/a_2_54# out_temp_decoded[13] OAI21X1_73/C vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1276 gnd INVX2_39/A AOI22X1_74/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M1277 AOI22X1_74/Y INVX2_39/Y AOI22X1_74/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M1278 AOI22X1_74/a_11_6# AOI22X1_74/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1279 AOI22X1_74/a_2_54# INVX2_39/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M1280 AOI22X1_74/a_28_6# INVX2_23/Y AOI22X1_74/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1281 vdd AOI22X1_74/A AOI22X1_74/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1282 AOI22X1_74/Y INVX2_23/Y AOI22X1_74/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M1283 AOI22X1_74/a_2_54# INVX2_39/A AOI22X1_74/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1284 gnd XOR2X1_18/Y AOI22X1_52/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M1285 XNOR2X1_25/B INVX2_45/A AOI22X1_52/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M1286 AOI22X1_52/a_11_6# XOR2X1_17/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1287 AOI22X1_52/a_2_54# INVX2_45/A vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M1288 AOI22X1_52/a_28_6# INVX2_48/A XNOR2X1_25/B Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1289 vdd XOR2X1_17/Y AOI22X1_52/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1290 XNOR2X1_25/B INVX2_48/A AOI22X1_52/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M1291 AOI22X1_52/a_2_54# XOR2X1_18/Y XNOR2X1_25/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1292 gnd NOR2X1_113/Y AOI22X1_63/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M1293 AOI22X1_63/Y out_mines[11] AOI22X1_63/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M1294 AOI22X1_63/a_11_6# NOR2X1_114/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1295 AOI22X1_63/a_2_54# out_mines[11] vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M1296 AOI22X1_63/a_28_6# out_mines[12] AOI22X1_63/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1297 vdd NOR2X1_114/Y AOI22X1_63/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1298 AOI22X1_63/Y out_mines[12] AOI22X1_63/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M1299 AOI22X1_63/a_2_54# NOR2X1_113/Y AOI22X1_63/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1300 gnd INVX2_10/Y OAI22X1_3/a_2_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=26u as=100p ps=50u
M1301 OAI22X1_3/a_2_6# INVX2_9/Y OAI22X1_3/Y Gnd nfet w=20 l=2
+  ad=100p pd=50u as=59.999996p ps=26u
M1302 OAI22X1_3/Y OAI22X1_3/D OAI22X1_3/a_2_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=26u as=59.999996p ps=26u
M1303 OAI22X1_3/Y OAI22X1_3/B OAI22X1_3/a_9_54# vdd pfet w=40 l=2
+  ad=0.24n pd=52u as=59.999996p ps=43u
M1304 OAI22X1_3/a_28_54# OAI22X1_3/D OAI22X1_3/Y vdd pfet w=40 l=2
+  ad=59.999996p pd=43u as=0.24n ps=52u
M1305 OAI22X1_3/a_9_54# INVX2_10/Y vdd vdd pfet w=40 l=2
+  ad=59.999996p pd=43u as=0.2n ps=90u
M1306 OAI22X1_3/a_2_6# OAI22X1_3/B gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=26u as=59.999996p ps=26u
M1307 vdd INVX2_9/Y OAI22X1_3/a_28_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=59.999996p ps=43u
M1308 INVX2_12/Y out_mines[13] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M1309 INVX2_12/Y out_mines[13] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.2n ps=90u
M1310 INVX2_34/Y INVX2_34/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1311 INVX2_34/Y INVX2_34/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1312 INVX2_23/Y out_mines[24] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1313 INVX2_23/Y out_mines[24] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1314 INVX2_45/Y INVX2_45/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1315 INVX2_45/Y INVX2_45/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1316 INVX2_56/Y out_temp_decoded[23] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1317 INVX2_56/Y out_temp_decoded[23] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1318 INVX2_67/Y out_temp_decoded[14] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1319 INVX2_67/Y out_temp_decoded[14] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1320 INVX2_78/Y out_temp_decoded[5] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1321 INVX2_78/Y out_temp_decoded[5] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1322 INVX2_89/Y out_temp_cleared[24] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1323 INVX2_89/Y out_temp_cleared[24] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1324 gnd INVX2_224/Y OAI21X1_19/a_2_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=26u as=100p ps=50u
M1325 vdd OAI21X1_19/C OAI21X1_19/Y vdd pfet w=20 l=2
+  ad=100p pd=50u as=0.11n ps=46u
M1326 OAI21X1_19/Y OAI21X1_19/C OAI21X1_19/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=59.999996p ps=26u
M1327 OAI21X1_19/Y OAI21X1_9/B OAI21X1_19/a_9_54# vdd pfet w=40 l=2
+  ad=0.11n pd=46u as=59.999996p ps=43u
M1328 OAI21X1_19/a_9_54# INVX2_224/Y vdd vdd pfet w=40 l=2
+  ad=59.999996p pd=43u as=0.2n ps=90u
M1329 OAI21X1_19/a_2_6# OAI21X1_9/B gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=26u as=59.999996p ps=26u
M1330 INVX2_190/Y INVX2_190/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1331 INVX2_190/Y INVX2_190/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1332 gnd NOR2X1_3/A XNOR2X1_6/a_2_6# Gnd nfet w=20 l=2
+  ad=70p pd=27u as=100p ps=50u
M1333 XNOR2X1_6/Y NOR2X1_3/A XNOR2X1_6/a_18_6# Gnd nfet w=20 l=2
+  ad=100p pd=30u as=29.999998p ps=23u
M1334 XNOR2X1_6/a_12_41# FAX1_1/YS gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=70p ps=27u
M1335 XNOR2X1_6/a_18_54# XNOR2X1_6/a_12_41# vdd vdd pfet w=40 l=2
+  ad=59.999996p pd=43u as=0.14n ps=47u
M1336 XNOR2X1_6/a_35_6# XNOR2X1_6/a_2_6# XNOR2X1_6/Y Gnd nfet w=20 l=2
+  ad=29.999998p pd=23u as=100p ps=30u
M1337 XNOR2X1_6/a_18_6# XNOR2X1_6/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=29.999998p pd=23u as=70p ps=27u
M1338 vdd NOR2X1_3/A XNOR2X1_6/a_2_6# vdd pfet w=40 l=2
+  ad=0.14n pd=47u as=0.2n ps=90u
M1339 vdd FAX1_1/YS XNOR2X1_6/a_35_54# vdd pfet w=40 l=2
+  ad=0.14n pd=47u as=59.999996p ps=43u
M1340 XNOR2X1_6/Y XNOR2X1_6/a_2_6# XNOR2X1_6/a_18_54# vdd pfet w=40 l=2
+  ad=0.2n pd=50u as=59.999996p ps=43u
M1341 XNOR2X1_6/a_35_54# NOR2X1_3/A XNOR2X1_6/Y vdd pfet w=40 l=2
+  ad=59.999996p pd=43u as=0.2n ps=50u
M1342 XNOR2X1_6/a_12_41# FAX1_1/YS vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.14n ps=47u
M1343 gnd FAX1_1/YS XNOR2X1_6/a_35_6# Gnd nfet w=20 l=2
+  ad=70p pd=27u as=29.999998p ps=23u
M1344 DFFNEGX1_30/a_76_6# BUFX2_15/Y DFFNEGX1_30/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1345 gnd BUFX2_15/Y DFFNEGX1_30/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1346 DFFNEGX1_30/a_66_6# DFFNEGX1_30/a_2_6# DFFNEGX1_30/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1347 out_mines[2] DFFNEGX1_30/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1348 DFFNEGX1_30/a_23_6# BUFX2_15/Y DFFNEGX1_30/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1349 DFFNEGX1_30/a_23_6# DFFNEGX1_30/a_2_6# DFFNEGX1_30/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1350 gnd DFFNEGX1_30/a_34_4# DFFNEGX1_30/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1351 vdd DFFNEGX1_30/a_34_4# DFFNEGX1_30/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1352 DFFNEGX1_30/a_61_74# DFFNEGX1_30/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1353 DFFNEGX1_30/a_34_4# DFFNEGX1_30/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1354 DFFNEGX1_30/a_34_4# DFFNEGX1_30/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1355 vdd out_mines[2] DFFNEGX1_30/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1356 gnd out_mines[2] DFFNEGX1_30/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1357 DFFNEGX1_30/a_61_6# DFFNEGX1_30/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1358 DFFNEGX1_30/a_76_84# DFFNEGX1_30/a_2_6# DFFNEGX1_30/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1359 out_mines[2] DFFNEGX1_30/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1360 vdd BUFX2_15/Y DFFNEGX1_30/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1361 DFFNEGX1_30/a_31_6# DFFNEGX1_30/a_2_6# DFFNEGX1_30/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1362 DFFNEGX1_30/a_66_6# BUFX2_15/Y DFFNEGX1_30/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1363 DFFNEGX1_30/a_17_74# OAI21X1_47/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1364 DFFNEGX1_30/a_31_74# BUFX2_15/Y DFFNEGX1_30/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1365 DFFNEGX1_30/a_17_6# OAI21X1_47/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1366 DFFNEGX1_52/a_76_6# BUFX2_14/Y DFFNEGX1_52/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1367 gnd BUFX2_14/Y DFFNEGX1_52/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1368 DFFNEGX1_52/a_66_6# DFFNEGX1_52/a_2_6# DFFNEGX1_52/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1369 out_temp_decoded[14] DFFNEGX1_52/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1370 DFFNEGX1_52/a_23_6# BUFX2_14/Y DFFNEGX1_52/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1371 DFFNEGX1_52/a_23_6# DFFNEGX1_52/a_2_6# DFFNEGX1_52/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1372 gnd DFFNEGX1_52/a_34_4# DFFNEGX1_52/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1373 vdd DFFNEGX1_52/a_34_4# DFFNEGX1_52/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1374 DFFNEGX1_52/a_61_74# DFFNEGX1_52/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1375 DFFNEGX1_52/a_34_4# DFFNEGX1_52/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1376 DFFNEGX1_52/a_34_4# DFFNEGX1_52/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1377 vdd out_temp_decoded[14] DFFNEGX1_52/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1378 gnd out_temp_decoded[14] DFFNEGX1_52/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1379 DFFNEGX1_52/a_61_6# DFFNEGX1_52/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1380 DFFNEGX1_52/a_76_84# DFFNEGX1_52/a_2_6# DFFNEGX1_52/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1381 out_temp_decoded[14] DFFNEGX1_52/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1382 vdd BUFX2_14/Y DFFNEGX1_52/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1383 DFFNEGX1_52/a_31_6# DFFNEGX1_52/a_2_6# DFFNEGX1_52/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1384 DFFNEGX1_52/a_66_6# BUFX2_14/Y DFFNEGX1_52/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1385 DFFNEGX1_52/a_17_74# OAI21X1_96/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1386 DFFNEGX1_52/a_31_74# BUFX2_14/Y DFFNEGX1_52/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1387 DFFNEGX1_52/a_17_6# OAI21X1_96/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1388 DFFNEGX1_41/a_76_6# BUFX2_14/Y DFFNEGX1_41/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1389 gnd BUFX2_14/Y DFFNEGX1_41/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1390 DFFNEGX1_41/a_66_6# DFFNEGX1_41/a_2_6# DFFNEGX1_41/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1391 out_temp_data_in[0] DFFNEGX1_41/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1392 DFFNEGX1_41/a_23_6# BUFX2_14/Y DFFNEGX1_41/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1393 DFFNEGX1_41/a_23_6# DFFNEGX1_41/a_2_6# DFFNEGX1_41/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1394 gnd DFFNEGX1_41/a_34_4# DFFNEGX1_41/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1395 vdd DFFNEGX1_41/a_34_4# DFFNEGX1_41/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1396 DFFNEGX1_41/a_61_74# DFFNEGX1_41/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1397 DFFNEGX1_41/a_34_4# DFFNEGX1_41/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1398 DFFNEGX1_41/a_34_4# DFFNEGX1_41/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1399 vdd out_temp_data_in[0] DFFNEGX1_41/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1400 gnd out_temp_data_in[0] DFFNEGX1_41/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1401 DFFNEGX1_41/a_61_6# DFFNEGX1_41/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1402 DFFNEGX1_41/a_76_84# DFFNEGX1_41/a_2_6# DFFNEGX1_41/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1403 out_temp_data_in[0] DFFNEGX1_41/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1404 vdd BUFX2_14/Y DFFNEGX1_41/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1405 DFFNEGX1_41/a_31_6# DFFNEGX1_41/a_2_6# DFFNEGX1_41/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1406 DFFNEGX1_41/a_66_6# BUFX2_14/Y DFFNEGX1_41/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1407 DFFNEGX1_41/a_17_74# OAI21X1_107/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1408 DFFNEGX1_41/a_31_74# BUFX2_14/Y DFFNEGX1_41/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1409 DFFNEGX1_41/a_17_6# OAI21X1_107/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1410 DFFNEGX1_74/a_76_6# BUFX2_12/Y DFFNEGX1_74/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1411 gnd BUFX2_12/Y DFFNEGX1_74/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1412 DFFNEGX1_74/a_66_6# DFFNEGX1_74/a_2_6# DFFNEGX1_74/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1413 out_temp_cleared[17] DFFNEGX1_74/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1414 DFFNEGX1_74/a_23_6# BUFX2_12/Y DFFNEGX1_74/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1415 DFFNEGX1_74/a_23_6# DFFNEGX1_74/a_2_6# DFFNEGX1_74/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1416 gnd DFFNEGX1_74/a_34_4# DFFNEGX1_74/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1417 vdd DFFNEGX1_74/a_34_4# DFFNEGX1_74/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1418 DFFNEGX1_74/a_61_74# DFFNEGX1_74/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1419 DFFNEGX1_74/a_34_4# DFFNEGX1_74/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1420 DFFNEGX1_74/a_34_4# DFFNEGX1_74/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1421 vdd out_temp_cleared[17] DFFNEGX1_74/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1422 gnd out_temp_cleared[17] DFFNEGX1_74/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1423 DFFNEGX1_74/a_61_6# DFFNEGX1_74/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1424 DFFNEGX1_74/a_76_84# DFFNEGX1_74/a_2_6# DFFNEGX1_74/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1425 out_temp_cleared[17] DFFNEGX1_74/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1426 vdd BUFX2_12/Y DFFNEGX1_74/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1427 DFFNEGX1_74/a_31_6# DFFNEGX1_74/a_2_6# DFFNEGX1_74/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1428 DFFNEGX1_74/a_66_6# BUFX2_12/Y DFFNEGX1_74/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1429 DFFNEGX1_74/a_17_74# OAI22X1_11/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1430 DFFNEGX1_74/a_31_74# BUFX2_12/Y DFFNEGX1_74/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1431 DFFNEGX1_74/a_17_6# OAI22X1_11/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1432 DFFNEGX1_85/a_76_6# BUFX2_11/Y DFFNEGX1_85/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1433 gnd BUFX2_11/Y DFFNEGX1_85/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1434 DFFNEGX1_85/a_66_6# DFFNEGX1_85/a_2_6# DFFNEGX1_85/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1435 out_temp_cleared[6] DFFNEGX1_85/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1436 DFFNEGX1_85/a_23_6# BUFX2_11/Y DFFNEGX1_85/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1437 DFFNEGX1_85/a_23_6# DFFNEGX1_85/a_2_6# DFFNEGX1_85/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1438 gnd DFFNEGX1_85/a_34_4# DFFNEGX1_85/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1439 vdd DFFNEGX1_85/a_34_4# DFFNEGX1_85/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1440 DFFNEGX1_85/a_61_74# DFFNEGX1_85/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1441 DFFNEGX1_85/a_34_4# DFFNEGX1_85/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1442 DFFNEGX1_85/a_34_4# DFFNEGX1_85/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1443 vdd out_temp_cleared[6] DFFNEGX1_85/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1444 gnd out_temp_cleared[6] DFFNEGX1_85/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1445 DFFNEGX1_85/a_61_6# DFFNEGX1_85/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1446 DFFNEGX1_85/a_76_84# DFFNEGX1_85/a_2_6# DFFNEGX1_85/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1447 out_temp_cleared[6] DFFNEGX1_85/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1448 vdd BUFX2_11/Y DFFNEGX1_85/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1449 DFFNEGX1_85/a_31_6# DFFNEGX1_85/a_2_6# DFFNEGX1_85/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1450 DFFNEGX1_85/a_66_6# BUFX2_11/Y DFFNEGX1_85/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1451 DFFNEGX1_85/a_17_74# OAI22X1_22/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1452 DFFNEGX1_85/a_31_74# BUFX2_11/Y DFFNEGX1_85/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1453 DFFNEGX1_85/a_17_6# OAI22X1_22/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1454 DFFNEGX1_63/a_76_6# BUFX2_13/Y DFFNEGX1_63/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1455 gnd BUFX2_13/Y DFFNEGX1_63/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1456 DFFNEGX1_63/a_66_6# DFFNEGX1_63/a_2_6# DFFNEGX1_63/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1457 out_temp_decoded[3] DFFNEGX1_63/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1458 DFFNEGX1_63/a_23_6# BUFX2_13/Y DFFNEGX1_63/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1459 DFFNEGX1_63/a_23_6# DFFNEGX1_63/a_2_6# DFFNEGX1_63/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1460 gnd DFFNEGX1_63/a_34_4# DFFNEGX1_63/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1461 vdd DFFNEGX1_63/a_34_4# DFFNEGX1_63/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1462 DFFNEGX1_63/a_61_74# DFFNEGX1_63/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1463 DFFNEGX1_63/a_34_4# DFFNEGX1_63/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1464 DFFNEGX1_63/a_34_4# DFFNEGX1_63/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1465 vdd out_temp_decoded[3] DFFNEGX1_63/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1466 gnd out_temp_decoded[3] DFFNEGX1_63/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1467 DFFNEGX1_63/a_61_6# DFFNEGX1_63/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1468 DFFNEGX1_63/a_76_84# DFFNEGX1_63/a_2_6# DFFNEGX1_63/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1469 out_temp_decoded[3] DFFNEGX1_63/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1470 vdd BUFX2_13/Y DFFNEGX1_63/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1471 DFFNEGX1_63/a_31_6# DFFNEGX1_63/a_2_6# DFFNEGX1_63/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1472 DFFNEGX1_63/a_66_6# BUFX2_13/Y DFFNEGX1_63/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1473 DFFNEGX1_63/a_17_74# OAI21X1_85/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1474 DFFNEGX1_63/a_31_74# BUFX2_13/Y DFFNEGX1_63/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1475 DFFNEGX1_63/a_17_6# OAI21X1_85/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1476 DFFNEGX1_96/a_76_6# BUFX2_10/Y DFFNEGX1_96/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1477 gnd BUFX2_10/Y DFFNEGX1_96/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1478 DFFNEGX1_96/a_66_6# DFFNEGX1_96/a_2_6# DFFNEGX1_96/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1479 out_global_score[2] DFFNEGX1_96/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1480 DFFNEGX1_96/a_23_6# BUFX2_10/Y DFFNEGX1_96/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1481 DFFNEGX1_96/a_23_6# DFFNEGX1_96/a_2_6# DFFNEGX1_96/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1482 gnd DFFNEGX1_96/a_34_4# DFFNEGX1_96/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1483 vdd DFFNEGX1_96/a_34_4# DFFNEGX1_96/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1484 DFFNEGX1_96/a_61_74# DFFNEGX1_96/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1485 DFFNEGX1_96/a_34_4# DFFNEGX1_96/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1486 DFFNEGX1_96/a_34_4# DFFNEGX1_96/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1487 vdd out_global_score[2] DFFNEGX1_96/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1488 gnd out_global_score[2] DFFNEGX1_96/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1489 DFFNEGX1_96/a_61_6# DFFNEGX1_96/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1490 DFFNEGX1_96/a_76_84# DFFNEGX1_96/a_2_6# DFFNEGX1_96/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1491 out_global_score[2] DFFNEGX1_96/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1492 vdd BUFX2_10/Y DFFNEGX1_96/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1493 DFFNEGX1_96/a_31_6# DFFNEGX1_96/a_2_6# DFFNEGX1_96/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1494 DFFNEGX1_96/a_66_6# BUFX2_10/Y DFFNEGX1_96/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1495 DFFNEGX1_96/a_17_74# INVX2_214/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1496 DFFNEGX1_96/a_31_74# BUFX2_10/Y DFFNEGX1_96/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1497 DFFNEGX1_96/a_17_6# INVX2_214/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1498 AND2X2_6/a_2_6# out_temp_data_in[4] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1499 AND2X2_6/a_9_6# out_temp_data_in[4] AND2X2_6/a_2_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=100p ps=50u
M1500 AND2X2_6/Y AND2X2_6/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1501 AND2X2_6/Y AND2X2_6/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1502 vdd AND2X2_6/B AND2X2_6/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1503 gnd AND2X2_6/B AND2X2_6/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1504 DFFNEGX1_120/a_76_6# BUFX2_5/Y DFFNEGX1_120/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1505 gnd BUFX2_5/Y DFFNEGX1_120/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1506 DFFNEGX1_120/a_66_6# DFFNEGX1_120/a_2_6# DFFNEGX1_120/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1507 out_global_score[26] DFFNEGX1_120/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1508 DFFNEGX1_120/a_23_6# BUFX2_5/Y DFFNEGX1_120/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1509 DFFNEGX1_120/a_23_6# DFFNEGX1_120/a_2_6# DFFNEGX1_120/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1510 gnd DFFNEGX1_120/a_34_4# DFFNEGX1_120/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1511 vdd DFFNEGX1_120/a_34_4# DFFNEGX1_120/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1512 DFFNEGX1_120/a_61_74# DFFNEGX1_120/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1513 DFFNEGX1_120/a_34_4# DFFNEGX1_120/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1514 DFFNEGX1_120/a_34_4# DFFNEGX1_120/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1515 vdd out_global_score[26] DFFNEGX1_120/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1516 gnd out_global_score[26] DFFNEGX1_120/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1517 DFFNEGX1_120/a_61_6# DFFNEGX1_120/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1518 DFFNEGX1_120/a_76_84# DFFNEGX1_120/a_2_6# DFFNEGX1_120/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1519 out_global_score[26] DFFNEGX1_120/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1520 vdd BUFX2_5/Y DFFNEGX1_120/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1521 DFFNEGX1_120/a_31_6# DFFNEGX1_120/a_2_6# DFFNEGX1_120/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1522 DFFNEGX1_120/a_66_6# BUFX2_5/Y DFFNEGX1_120/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1523 DFFNEGX1_120/a_17_74# INVX2_190/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1524 DFFNEGX1_120/a_31_74# BUFX2_5/Y DFFNEGX1_120/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1525 DFFNEGX1_120/a_17_6# INVX2_190/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1526 gnd XNOR2X1_6/Y MUX2X1_18/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M1527 MUX2X1_18/a_17_50# NOR2X1_3/A vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1528 XNOR2X1_5/A OR2X1_3/Y MUX2X1_18/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M1529 MUX2X1_18/a_30_54# MUX2X1_18/a_2_10# XNOR2X1_5/A vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1530 MUX2X1_18/a_17_10# NOR2X1_3/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1531 vdd OR2X1_3/Y MUX2X1_18/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1532 MUX2X1_18/a_30_10# OR2X1_3/Y XNOR2X1_5/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M1533 gnd OR2X1_3/Y MUX2X1_18/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M1534 vdd XNOR2X1_6/Y MUX2X1_18/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1535 XNOR2X1_5/A MUX2X1_18/a_2_10# MUX2X1_18/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1536 DFFNEGX1_142/a_76_6# INVX2_259/Y DFFNEGX1_142/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1537 gnd INVX2_259/Y DFFNEGX1_142/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1538 DFFNEGX1_142/a_66_6# DFFNEGX1_142/a_2_6# DFFNEGX1_142/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1539 out_display DFFNEGX1_142/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1540 DFFNEGX1_142/a_23_6# INVX2_259/Y DFFNEGX1_142/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1541 DFFNEGX1_142/a_23_6# DFFNEGX1_142/a_2_6# DFFNEGX1_142/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1542 gnd DFFNEGX1_142/a_34_4# DFFNEGX1_142/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1543 vdd DFFNEGX1_142/a_34_4# DFFNEGX1_142/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1544 DFFNEGX1_142/a_61_74# DFFNEGX1_142/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1545 DFFNEGX1_142/a_34_4# DFFNEGX1_142/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1546 DFFNEGX1_142/a_34_4# DFFNEGX1_142/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1547 vdd out_display DFFNEGX1_142/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1548 gnd out_display DFFNEGX1_142/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1549 DFFNEGX1_142/a_61_6# DFFNEGX1_142/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1550 DFFNEGX1_142/a_76_84# DFFNEGX1_142/a_2_6# DFFNEGX1_142/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1551 out_display DFFNEGX1_142/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1552 vdd INVX2_259/Y DFFNEGX1_142/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1553 DFFNEGX1_142/a_31_6# DFFNEGX1_142/a_2_6# DFFNEGX1_142/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1554 DFFNEGX1_142/a_66_6# INVX2_259/Y DFFNEGX1_142/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1555 DFFNEGX1_142/a_17_74# OAI21X1_155/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1556 DFFNEGX1_142/a_31_74# INVX2_259/Y DFFNEGX1_142/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1557 DFFNEGX1_142/a_17_6# OAI21X1_155/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1558 DFFNEGX1_131/a_76_6# BUFX2_5/Y DFFNEGX1_131/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1559 gnd BUFX2_5/Y DFFNEGX1_131/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1560 DFFNEGX1_131/a_66_6# DFFNEGX1_131/a_2_6# DFFNEGX1_131/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1561 INVX2_117/A DFFNEGX1_131/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1562 DFFNEGX1_131/a_23_6# BUFX2_5/Y DFFNEGX1_131/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1563 DFFNEGX1_131/a_23_6# DFFNEGX1_131/a_2_6# DFFNEGX1_131/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1564 gnd DFFNEGX1_131/a_34_4# DFFNEGX1_131/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1565 vdd DFFNEGX1_131/a_34_4# DFFNEGX1_131/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1566 DFFNEGX1_131/a_61_74# DFFNEGX1_131/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1567 DFFNEGX1_131/a_34_4# DFFNEGX1_131/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1568 DFFNEGX1_131/a_34_4# DFFNEGX1_131/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1569 vdd INVX2_117/A DFFNEGX1_131/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1570 gnd INVX2_117/A DFFNEGX1_131/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1571 DFFNEGX1_131/a_61_6# DFFNEGX1_131/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1572 DFFNEGX1_131/a_76_84# DFFNEGX1_131/a_2_6# DFFNEGX1_131/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1573 INVX2_117/A DFFNEGX1_131/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1574 vdd BUFX2_5/Y DFFNEGX1_131/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1575 DFFNEGX1_131/a_31_6# DFFNEGX1_131/a_2_6# DFFNEGX1_131/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1576 DFFNEGX1_131/a_66_6# BUFX2_5/Y DFFNEGX1_131/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1577 DFFNEGX1_131/a_17_74# AOI21X1_20/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1578 DFFNEGX1_131/a_31_74# BUFX2_5/Y DFFNEGX1_131/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1579 DFFNEGX1_131/a_17_6# AOI21X1_20/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1580 gnd MUX2X1_29/A MUX2X1_29/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M1581 MUX2X1_29/a_17_50# FAX1_3/YS vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1582 MUX2X1_29/Y OR2X1_1/Y MUX2X1_29/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M1583 MUX2X1_29/a_30_54# MUX2X1_29/a_2_10# MUX2X1_29/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1584 MUX2X1_29/a_17_10# FAX1_3/YS gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1585 vdd OR2X1_1/Y MUX2X1_29/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1586 MUX2X1_29/a_30_10# OR2X1_1/Y MUX2X1_29/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M1587 gnd OR2X1_1/Y MUX2X1_29/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M1588 vdd MUX2X1_29/A MUX2X1_29/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1589 MUX2X1_29/Y MUX2X1_29/a_2_10# MUX2X1_29/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1590 gnd OR2X1_14/B AOI22X1_1/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M1591 INVX2_88/A INVX2_86/Y AOI22X1_1/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M1592 AOI22X1_1/a_11_6# AOI22X1_1/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1593 AOI22X1_1/a_2_54# INVX2_86/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M1594 AOI22X1_1/a_28_6# XOR2X1_23/Y INVX2_88/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1595 vdd AOI22X1_1/A AOI22X1_1/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1596 INVX2_88/A XOR2X1_23/Y AOI22X1_1/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M1597 AOI22X1_1/a_2_54# OR2X1_14/B INVX2_88/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1598 OAI21X1_32/B NOR2X1_62/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1599 NAND2X1_33/a_9_6# NOR2X1_62/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1600 vdd NOR2X1_63/B OAI21X1_32/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1601 OAI21X1_32/B NOR2X1_63/B NAND2X1_33/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1602 OAI21X1_15/C out_mines[18] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1603 NAND2X1_22/a_9_6# out_mines[18] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1604 vdd INVX2_240/Y OAI21X1_15/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1605 OAI21X1_15/C INVX2_240/Y NAND2X1_22/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1606 NOR2X1_55/A out_temp_data_in[0] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1607 NAND2X1_11/a_9_6# out_temp_data_in[0] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1608 vdd OR2X1_6/A NOR2X1_55/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1609 NOR2X1_55/A OR2X1_6/A NAND2X1_11/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1610 OAI21X1_47/C out_mines[2] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1611 NAND2X1_44/a_9_6# out_mines[2] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1612 vdd INVX2_244/Y OAI21X1_47/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1613 OAI21X1_47/C INVX2_244/Y NAND2X1_44/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1614 OAI21X1_90/C NOR2X1_36/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1615 NAND2X1_77/a_9_6# NOR2X1_36/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1616 vdd BUFX2_20/Y OAI21X1_90/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1617 OAI21X1_90/C BUFX2_20/Y NAND2X1_77/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1618 OAI21X1_77/B INVX2_91/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1619 NAND2X1_66/a_9_6# INVX2_91/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1620 vdd INVX2_57/Y OAI21X1_77/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1621 OAI21X1_77/B INVX2_57/Y NAND2X1_66/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1622 OAI21X1_59/C out_display_done vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1623 NAND2X1_55/a_9_6# out_display_done gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1624 vdd INVX2_184/Y OAI21X1_59/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1625 OAI21X1_59/C INVX2_184/Y NAND2X1_55/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1626 NAND2X1_88/Y NOR2X1_49/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1627 NAND2X1_88/a_9_6# NOR2X1_49/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1628 vdd BUFX2_21/Y NAND2X1_88/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1629 NAND2X1_88/Y BUFX2_21/Y NAND2X1_88/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1630 NAND2X1_99/Y in_data[3] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1631 NAND2X1_99/a_9_6# in_data[3] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1632 vdd NOR2X1_107/Y NAND2X1_99/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1633 NAND2X1_99/Y NOR2X1_107/Y NAND2X1_99/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1634 gnd out_global_score[13] AOI22X1_20/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M1635 INVX2_203/A INVX2_257/Y AOI22X1_20/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M1636 AOI22X1_20/a_11_6# HAX1_17/YS gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1637 AOI22X1_20/a_2_54# INVX2_257/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M1638 AOI22X1_20/a_28_6# OR2X1_11/B INVX2_203/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1639 vdd HAX1_17/YS AOI22X1_20/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1640 INVX2_203/A OR2X1_11/B AOI22X1_20/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M1641 AOI22X1_20/a_2_54# out_global_score[13] INVX2_203/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1642 gnd out_global_score[2] AOI22X1_31/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M1643 INVX2_214/A INVX2_258/Y AOI22X1_31/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M1644 AOI22X1_31/a_11_6# HAX1_28/YS gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1645 AOI22X1_31/a_2_54# INVX2_258/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M1646 AOI22X1_31/a_28_6# OR2X1_11/B INVX2_214/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1647 vdd HAX1_28/YS AOI22X1_31/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1648 INVX2_214/A OR2X1_11/B AOI22X1_31/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M1649 AOI22X1_31/a_2_54# out_global_score[2] INVX2_214/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1650 gnd out_temp_cleared[11] AOI22X1_42/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M1651 OAI21X1_74/C out_mines[10] AOI22X1_42/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M1652 AOI22X1_42/a_11_6# out_temp_cleared[10] gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1653 AOI22X1_42/a_2_54# out_mines[10] vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M1654 AOI22X1_42/a_28_6# out_mines[11] OAI21X1_74/C Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1655 vdd out_temp_cleared[10] AOI22X1_42/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1656 OAI21X1_74/C out_mines[11] AOI22X1_42/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M1657 AOI22X1_42/a_2_54# out_temp_cleared[11] OAI21X1_74/C vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1658 gnd INVX2_36/A AOI22X1_75/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M1659 AOI22X1_75/Y INVX2_36/Y AOI22X1_75/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M1660 AOI22X1_75/a_11_6# AOI22X1_75/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1661 AOI22X1_75/a_2_54# INVX2_36/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M1662 AOI22X1_75/a_28_6# INVX2_23/Y AOI22X1_75/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1663 vdd AOI22X1_75/A AOI22X1_75/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1664 AOI22X1_75/Y INVX2_23/Y AOI22X1_75/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M1665 AOI22X1_75/a_2_54# INVX2_36/A AOI22X1_75/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1666 gnd XOR2X1_28/Y AOI22X1_53/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M1667 XNOR2X1_27/B INVX2_48/A AOI22X1_53/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M1668 AOI22X1_53/a_11_6# XOR2X1_27/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1669 AOI22X1_53/a_2_54# INVX2_48/A vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M1670 AOI22X1_53/a_28_6# INVX2_44/A XNOR2X1_27/B Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1671 vdd XOR2X1_27/Y AOI22X1_53/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1672 XNOR2X1_27/B INVX2_44/A AOI22X1_53/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M1673 AOI22X1_53/a_2_54# XOR2X1_28/Y XNOR2X1_27/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1674 gnd NOR2X1_111/Y AOI22X1_64/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M1675 AOI22X1_64/Y out_mines[17] AOI22X1_64/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M1676 AOI22X1_64/a_11_6# NOR2X1_112/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1677 AOI22X1_64/a_2_54# out_mines[17] vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M1678 AOI22X1_64/a_28_6# out_mines[18] AOI22X1_64/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1679 vdd NOR2X1_112/Y AOI22X1_64/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1680 AOI22X1_64/Y out_mines[18] AOI22X1_64/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M1681 AOI22X1_64/a_2_54# NOR2X1_111/Y AOI22X1_64/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1682 gnd BUFX2_25/A OAI22X1_4/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M1683 OAI22X1_4/a_2_6# OR2X1_11/A OAI22X1_4/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M1684 OAI22X1_4/Y INVX2_55/Y OAI22X1_4/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1685 OAI22X1_4/Y INVX2_89/Y OAI22X1_4/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M1686 OAI22X1_4/a_28_54# INVX2_55/Y OAI22X1_4/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1687 OAI22X1_4/a_9_54# BUFX2_25/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1688 OAI22X1_4/a_2_6# INVX2_89/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1689 vdd OR2X1_11/A OAI22X1_4/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1690 INVX2_13/Y out_mines[14] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1691 INVX2_13/Y out_mines[14] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1692 INVX2_24/Y out_mines[19] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1693 INVX2_24/Y out_mines[19] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1694 INVX2_35/Y XOR2X1_4/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1695 INVX2_35/Y XOR2X1_4/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1696 INVX2_68/Y out_temp_decoded[13] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1697 INVX2_68/Y out_temp_decoded[13] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1698 INVX2_57/Y out_temp_decoded[22] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1699 INVX2_57/Y out_temp_decoded[22] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1700 INVX2_79/Y out_temp_decoded[4] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1701 INVX2_79/Y out_temp_decoded[4] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1702 INVX2_46/Y INVX2_46/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1703 INVX2_46/Y INVX2_46/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1704 INVX2_180/Y NOR2X1_61/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1705 INVX2_180/Y NOR2X1_61/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1706 INVX2_191/Y INVX2_191/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1707 INVX2_191/Y INVX2_191/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1708 gnd XNOR2X1_7/A XNOR2X1_7/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1709 XNOR2X1_7/Y XNOR2X1_7/A XNOR2X1_7/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M1710 XNOR2X1_7/a_12_41# NOR2X1_3/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1711 XNOR2X1_7/a_18_54# XNOR2X1_7/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1712 XNOR2X1_7/a_35_6# XNOR2X1_7/a_2_6# XNOR2X1_7/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1713 XNOR2X1_7/a_18_6# XNOR2X1_7/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1714 vdd XNOR2X1_7/A XNOR2X1_7/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1715 vdd NOR2X1_3/Y XNOR2X1_7/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M1716 XNOR2X1_7/Y XNOR2X1_7/a_2_6# XNOR2X1_7/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M1717 XNOR2X1_7/a_35_54# XNOR2X1_7/A XNOR2X1_7/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1718 XNOR2X1_7/a_12_41# NOR2X1_3/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1719 gnd NOR2X1_3/Y XNOR2X1_7/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1720 DFFNEGX1_31/a_76_6# BUFX2_15/Y DFFNEGX1_31/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1721 gnd BUFX2_15/Y DFFNEGX1_31/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1722 DFFNEGX1_31/a_66_6# DFFNEGX1_31/a_2_6# DFFNEGX1_31/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1723 out_temp_mine_cnt[0] DFFNEGX1_31/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1724 DFFNEGX1_31/a_23_6# BUFX2_15/Y DFFNEGX1_31/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1725 DFFNEGX1_31/a_23_6# DFFNEGX1_31/a_2_6# DFFNEGX1_31/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1726 gnd DFFNEGX1_31/a_34_4# DFFNEGX1_31/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1727 vdd DFFNEGX1_31/a_34_4# DFFNEGX1_31/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1728 DFFNEGX1_31/a_61_74# DFFNEGX1_31/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1729 DFFNEGX1_31/a_34_4# DFFNEGX1_31/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1730 DFFNEGX1_31/a_34_4# DFFNEGX1_31/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1731 vdd out_temp_mine_cnt[0] DFFNEGX1_31/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1732 gnd out_temp_mine_cnt[0] DFFNEGX1_31/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1733 DFFNEGX1_31/a_61_6# DFFNEGX1_31/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1734 DFFNEGX1_31/a_76_84# DFFNEGX1_31/a_2_6# DFFNEGX1_31/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1735 out_temp_mine_cnt[0] DFFNEGX1_31/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1736 vdd BUFX2_15/Y DFFNEGX1_31/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1737 DFFNEGX1_31/a_31_6# DFFNEGX1_31/a_2_6# DFFNEGX1_31/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1738 DFFNEGX1_31/a_66_6# BUFX2_15/Y DFFNEGX1_31/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1739 DFFNEGX1_31/a_17_74# AND2X2_13/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1740 DFFNEGX1_31/a_31_74# BUFX2_15/Y DFFNEGX1_31/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1741 DFFNEGX1_31/a_17_6# AND2X2_13/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1742 DFFNEGX1_20/a_76_6# BUFX2_16/Y DFFNEGX1_20/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1743 gnd BUFX2_16/Y DFFNEGX1_20/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1744 DFFNEGX1_20/a_66_6# DFFNEGX1_20/a_2_6# DFFNEGX1_20/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1745 out_mines[22] DFFNEGX1_20/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1746 DFFNEGX1_20/a_23_6# BUFX2_16/Y DFFNEGX1_20/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1747 DFFNEGX1_20/a_23_6# DFFNEGX1_20/a_2_6# DFFNEGX1_20/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1748 gnd DFFNEGX1_20/a_34_4# DFFNEGX1_20/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1749 vdd DFFNEGX1_20/a_34_4# DFFNEGX1_20/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1750 DFFNEGX1_20/a_61_74# DFFNEGX1_20/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1751 DFFNEGX1_20/a_34_4# DFFNEGX1_20/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1752 DFFNEGX1_20/a_34_4# DFFNEGX1_20/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1753 vdd out_mines[22] DFFNEGX1_20/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1754 gnd out_mines[22] DFFNEGX1_20/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1755 DFFNEGX1_20/a_61_6# DFFNEGX1_20/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1756 DFFNEGX1_20/a_76_84# DFFNEGX1_20/a_2_6# DFFNEGX1_20/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1757 out_mines[22] DFFNEGX1_20/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1758 vdd BUFX2_16/Y DFFNEGX1_20/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1759 DFFNEGX1_20/a_31_6# DFFNEGX1_20/a_2_6# DFFNEGX1_20/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1760 DFFNEGX1_20/a_66_6# BUFX2_16/Y DFFNEGX1_20/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1761 DFFNEGX1_20/a_17_74# OAI21X1_7/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1762 DFFNEGX1_20/a_31_74# BUFX2_16/Y DFFNEGX1_20/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1763 DFFNEGX1_20/a_17_6# OAI21X1_7/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1764 DFFNEGX1_42/a_76_6# BUFX2_14/Y DFFNEGX1_42/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1765 gnd BUFX2_14/Y DFFNEGX1_42/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1766 DFFNEGX1_42/a_66_6# DFFNEGX1_42/a_2_6# DFFNEGX1_42/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1767 out_temp_decoded[24] DFFNEGX1_42/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1768 DFFNEGX1_42/a_23_6# BUFX2_14/Y DFFNEGX1_42/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1769 DFFNEGX1_42/a_23_6# DFFNEGX1_42/a_2_6# DFFNEGX1_42/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1770 gnd DFFNEGX1_42/a_34_4# DFFNEGX1_42/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1771 vdd DFFNEGX1_42/a_34_4# DFFNEGX1_42/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1772 DFFNEGX1_42/a_61_74# DFFNEGX1_42/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1773 DFFNEGX1_42/a_34_4# DFFNEGX1_42/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1774 DFFNEGX1_42/a_34_4# DFFNEGX1_42/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1775 vdd out_temp_decoded[24] DFFNEGX1_42/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1776 gnd out_temp_decoded[24] DFFNEGX1_42/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1777 DFFNEGX1_42/a_61_6# DFFNEGX1_42/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1778 DFFNEGX1_42/a_76_84# DFFNEGX1_42/a_2_6# DFFNEGX1_42/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1779 out_temp_decoded[24] DFFNEGX1_42/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1780 vdd BUFX2_14/Y DFFNEGX1_42/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1781 DFFNEGX1_42/a_31_6# DFFNEGX1_42/a_2_6# DFFNEGX1_42/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1782 DFFNEGX1_42/a_66_6# BUFX2_14/Y DFFNEGX1_42/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1783 DFFNEGX1_42/a_17_74# OAI21X1_106/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1784 DFFNEGX1_42/a_31_74# BUFX2_14/Y DFFNEGX1_42/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1785 DFFNEGX1_42/a_17_6# OAI21X1_106/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1786 DFFNEGX1_53/a_76_6# BUFX2_14/Y DFFNEGX1_53/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1787 gnd BUFX2_14/Y DFFNEGX1_53/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1788 DFFNEGX1_53/a_66_6# DFFNEGX1_53/a_2_6# DFFNEGX1_53/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1789 out_temp_decoded[13] DFFNEGX1_53/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1790 DFFNEGX1_53/a_23_6# BUFX2_14/Y DFFNEGX1_53/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1791 DFFNEGX1_53/a_23_6# DFFNEGX1_53/a_2_6# DFFNEGX1_53/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1792 gnd DFFNEGX1_53/a_34_4# DFFNEGX1_53/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1793 vdd DFFNEGX1_53/a_34_4# DFFNEGX1_53/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1794 DFFNEGX1_53/a_61_74# DFFNEGX1_53/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1795 DFFNEGX1_53/a_34_4# DFFNEGX1_53/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1796 DFFNEGX1_53/a_34_4# DFFNEGX1_53/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1797 vdd out_temp_decoded[13] DFFNEGX1_53/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1798 gnd out_temp_decoded[13] DFFNEGX1_53/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1799 DFFNEGX1_53/a_61_6# DFFNEGX1_53/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1800 DFFNEGX1_53/a_76_84# DFFNEGX1_53/a_2_6# DFFNEGX1_53/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1801 out_temp_decoded[13] DFFNEGX1_53/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1802 vdd BUFX2_14/Y DFFNEGX1_53/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1803 DFFNEGX1_53/a_31_6# DFFNEGX1_53/a_2_6# DFFNEGX1_53/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1804 DFFNEGX1_53/a_66_6# BUFX2_14/Y DFFNEGX1_53/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1805 DFFNEGX1_53/a_17_74# OAI21X1_95/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1806 DFFNEGX1_53/a_31_74# BUFX2_14/Y DFFNEGX1_53/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1807 DFFNEGX1_53/a_17_6# OAI21X1_95/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1808 DFFNEGX1_75/a_76_6# BUFX2_12/Y DFFNEGX1_75/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1809 gnd BUFX2_12/Y DFFNEGX1_75/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1810 DFFNEGX1_75/a_66_6# DFFNEGX1_75/a_2_6# DFFNEGX1_75/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1811 out_temp_cleared[16] DFFNEGX1_75/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1812 DFFNEGX1_75/a_23_6# BUFX2_12/Y DFFNEGX1_75/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1813 DFFNEGX1_75/a_23_6# DFFNEGX1_75/a_2_6# DFFNEGX1_75/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1814 gnd DFFNEGX1_75/a_34_4# DFFNEGX1_75/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1815 vdd DFFNEGX1_75/a_34_4# DFFNEGX1_75/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1816 DFFNEGX1_75/a_61_74# DFFNEGX1_75/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1817 DFFNEGX1_75/a_34_4# DFFNEGX1_75/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1818 DFFNEGX1_75/a_34_4# DFFNEGX1_75/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1819 vdd out_temp_cleared[16] DFFNEGX1_75/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1820 gnd out_temp_cleared[16] DFFNEGX1_75/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1821 DFFNEGX1_75/a_61_6# DFFNEGX1_75/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1822 DFFNEGX1_75/a_76_84# DFFNEGX1_75/a_2_6# DFFNEGX1_75/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1823 out_temp_cleared[16] DFFNEGX1_75/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1824 vdd BUFX2_12/Y DFFNEGX1_75/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1825 DFFNEGX1_75/a_31_6# DFFNEGX1_75/a_2_6# DFFNEGX1_75/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1826 DFFNEGX1_75/a_66_6# BUFX2_12/Y DFFNEGX1_75/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1827 DFFNEGX1_75/a_17_74# OAI22X1_12/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1828 DFFNEGX1_75/a_31_74# BUFX2_12/Y DFFNEGX1_75/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1829 DFFNEGX1_75/a_17_6# OAI22X1_12/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1830 DFFNEGX1_64/a_76_6# BUFX2_13/Y DFFNEGX1_64/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1831 gnd BUFX2_13/Y DFFNEGX1_64/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1832 DFFNEGX1_64/a_66_6# DFFNEGX1_64/a_2_6# DFFNEGX1_64/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1833 out_temp_decoded[2] DFFNEGX1_64/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1834 DFFNEGX1_64/a_23_6# BUFX2_13/Y DFFNEGX1_64/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1835 DFFNEGX1_64/a_23_6# DFFNEGX1_64/a_2_6# DFFNEGX1_64/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1836 gnd DFFNEGX1_64/a_34_4# DFFNEGX1_64/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1837 vdd DFFNEGX1_64/a_34_4# DFFNEGX1_64/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1838 DFFNEGX1_64/a_61_74# DFFNEGX1_64/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1839 DFFNEGX1_64/a_34_4# DFFNEGX1_64/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1840 DFFNEGX1_64/a_34_4# DFFNEGX1_64/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1841 vdd out_temp_decoded[2] DFFNEGX1_64/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1842 gnd out_temp_decoded[2] DFFNEGX1_64/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1843 DFFNEGX1_64/a_61_6# DFFNEGX1_64/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1844 DFFNEGX1_64/a_76_84# DFFNEGX1_64/a_2_6# DFFNEGX1_64/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1845 out_temp_decoded[2] DFFNEGX1_64/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1846 vdd BUFX2_13/Y DFFNEGX1_64/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1847 DFFNEGX1_64/a_31_6# DFFNEGX1_64/a_2_6# DFFNEGX1_64/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1848 DFFNEGX1_64/a_66_6# BUFX2_13/Y DFFNEGX1_64/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1849 DFFNEGX1_64/a_17_74# OAI21X1_84/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1850 DFFNEGX1_64/a_31_74# BUFX2_13/Y DFFNEGX1_64/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1851 DFFNEGX1_64/a_17_6# OAI21X1_84/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1852 DFFNEGX1_86/a_76_6# BUFX2_11/Y DFFNEGX1_86/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1853 gnd BUFX2_11/Y DFFNEGX1_86/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1854 DFFNEGX1_86/a_66_6# DFFNEGX1_86/a_2_6# DFFNEGX1_86/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1855 out_temp_cleared[5] DFFNEGX1_86/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1856 DFFNEGX1_86/a_23_6# BUFX2_11/Y DFFNEGX1_86/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1857 DFFNEGX1_86/a_23_6# DFFNEGX1_86/a_2_6# DFFNEGX1_86/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1858 gnd DFFNEGX1_86/a_34_4# DFFNEGX1_86/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1859 vdd DFFNEGX1_86/a_34_4# DFFNEGX1_86/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1860 DFFNEGX1_86/a_61_74# DFFNEGX1_86/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1861 DFFNEGX1_86/a_34_4# DFFNEGX1_86/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1862 DFFNEGX1_86/a_34_4# DFFNEGX1_86/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1863 vdd out_temp_cleared[5] DFFNEGX1_86/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1864 gnd out_temp_cleared[5] DFFNEGX1_86/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1865 DFFNEGX1_86/a_61_6# DFFNEGX1_86/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1866 DFFNEGX1_86/a_76_84# DFFNEGX1_86/a_2_6# DFFNEGX1_86/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1867 out_temp_cleared[5] DFFNEGX1_86/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1868 vdd BUFX2_11/Y DFFNEGX1_86/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1869 DFFNEGX1_86/a_31_6# DFFNEGX1_86/a_2_6# DFFNEGX1_86/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1870 DFFNEGX1_86/a_66_6# BUFX2_11/Y DFFNEGX1_86/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1871 DFFNEGX1_86/a_17_74# OAI22X1_23/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1872 DFFNEGX1_86/a_31_74# BUFX2_11/Y DFFNEGX1_86/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1873 DFFNEGX1_86/a_17_6# OAI22X1_23/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1874 DFFNEGX1_97/a_76_6# BUFX2_10/Y DFFNEGX1_97/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1875 gnd BUFX2_10/Y DFFNEGX1_97/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1876 DFFNEGX1_97/a_66_6# DFFNEGX1_97/a_2_6# DFFNEGX1_97/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1877 out_global_score[3] DFFNEGX1_97/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1878 DFFNEGX1_97/a_23_6# BUFX2_10/Y DFFNEGX1_97/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1879 DFFNEGX1_97/a_23_6# DFFNEGX1_97/a_2_6# DFFNEGX1_97/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1880 gnd DFFNEGX1_97/a_34_4# DFFNEGX1_97/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1881 vdd DFFNEGX1_97/a_34_4# DFFNEGX1_97/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1882 DFFNEGX1_97/a_61_74# DFFNEGX1_97/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1883 DFFNEGX1_97/a_34_4# DFFNEGX1_97/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1884 DFFNEGX1_97/a_34_4# DFFNEGX1_97/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1885 vdd out_global_score[3] DFFNEGX1_97/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1886 gnd out_global_score[3] DFFNEGX1_97/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1887 DFFNEGX1_97/a_61_6# DFFNEGX1_97/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1888 DFFNEGX1_97/a_76_84# DFFNEGX1_97/a_2_6# DFFNEGX1_97/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1889 out_global_score[3] DFFNEGX1_97/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1890 vdd BUFX2_10/Y DFFNEGX1_97/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1891 DFFNEGX1_97/a_31_6# DFFNEGX1_97/a_2_6# DFFNEGX1_97/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1892 DFFNEGX1_97/a_66_6# BUFX2_10/Y DFFNEGX1_97/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1893 DFFNEGX1_97/a_17_74# INVX2_213/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1894 DFFNEGX1_97/a_31_74# BUFX2_10/Y DFFNEGX1_97/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1895 DFFNEGX1_97/a_17_6# INVX2_213/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1896 AND2X2_7/a_2_6# XOR2X1_6/A vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1897 AND2X2_7/a_9_6# XOR2X1_6/A AND2X2_7/a_2_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=100p ps=50u
M1898 XOR2X1_5/A AND2X2_7/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1899 XOR2X1_5/A AND2X2_7/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1900 vdd FAX1_4/YS AND2X2_7/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1901 gnd FAX1_4/YS AND2X2_7/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1902 DFFNEGX1_110/a_76_6# BUFX2_9/Y DFFNEGX1_110/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1903 gnd BUFX2_9/Y DFFNEGX1_110/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1904 DFFNEGX1_110/a_66_6# DFFNEGX1_110/a_2_6# DFFNEGX1_110/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1905 out_global_score[16] DFFNEGX1_110/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1906 DFFNEGX1_110/a_23_6# BUFX2_9/Y DFFNEGX1_110/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1907 DFFNEGX1_110/a_23_6# DFFNEGX1_110/a_2_6# DFFNEGX1_110/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1908 gnd DFFNEGX1_110/a_34_4# DFFNEGX1_110/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1909 vdd DFFNEGX1_110/a_34_4# DFFNEGX1_110/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1910 DFFNEGX1_110/a_61_74# DFFNEGX1_110/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1911 DFFNEGX1_110/a_34_4# DFFNEGX1_110/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1912 DFFNEGX1_110/a_34_4# DFFNEGX1_110/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1913 vdd out_global_score[16] DFFNEGX1_110/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1914 gnd out_global_score[16] DFFNEGX1_110/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1915 DFFNEGX1_110/a_61_6# DFFNEGX1_110/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1916 DFFNEGX1_110/a_76_84# DFFNEGX1_110/a_2_6# DFFNEGX1_110/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1917 out_global_score[16] DFFNEGX1_110/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1918 vdd BUFX2_9/Y DFFNEGX1_110/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1919 DFFNEGX1_110/a_31_6# DFFNEGX1_110/a_2_6# DFFNEGX1_110/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1920 DFFNEGX1_110/a_66_6# BUFX2_9/Y DFFNEGX1_110/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1921 DFFNEGX1_110/a_17_74# INVX2_200/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1922 DFFNEGX1_110/a_31_74# BUFX2_9/Y DFFNEGX1_110/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1923 DFFNEGX1_110/a_17_6# INVX2_200/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1924 DFFNEGX1_121/a_76_6# BUFX2_5/Y DFFNEGX1_121/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1925 gnd BUFX2_5/Y DFFNEGX1_121/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1926 DFFNEGX1_121/a_66_6# DFFNEGX1_121/a_2_6# DFFNEGX1_121/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1927 out_global_score[27] DFFNEGX1_121/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1928 DFFNEGX1_121/a_23_6# BUFX2_5/Y DFFNEGX1_121/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1929 DFFNEGX1_121/a_23_6# DFFNEGX1_121/a_2_6# DFFNEGX1_121/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1930 gnd DFFNEGX1_121/a_34_4# DFFNEGX1_121/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1931 vdd DFFNEGX1_121/a_34_4# DFFNEGX1_121/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1932 DFFNEGX1_121/a_61_74# DFFNEGX1_121/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1933 DFFNEGX1_121/a_34_4# DFFNEGX1_121/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1934 DFFNEGX1_121/a_34_4# DFFNEGX1_121/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1935 vdd out_global_score[27] DFFNEGX1_121/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1936 gnd out_global_score[27] DFFNEGX1_121/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1937 DFFNEGX1_121/a_61_6# DFFNEGX1_121/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1938 DFFNEGX1_121/a_76_84# DFFNEGX1_121/a_2_6# DFFNEGX1_121/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1939 out_global_score[27] DFFNEGX1_121/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1940 vdd BUFX2_5/Y DFFNEGX1_121/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1941 DFFNEGX1_121/a_31_6# DFFNEGX1_121/a_2_6# DFFNEGX1_121/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1942 DFFNEGX1_121/a_66_6# BUFX2_5/Y DFFNEGX1_121/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1943 DFFNEGX1_121/a_17_74# INVX2_189/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1944 DFFNEGX1_121/a_31_74# BUFX2_5/Y DFFNEGX1_121/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1945 DFFNEGX1_121/a_17_6# INVX2_189/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1946 DFFNEGX1_132/a_76_6# INVX2_259/Y DFFNEGX1_132/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M1947 gnd INVX2_259/Y DFFNEGX1_132/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1948 DFFNEGX1_132/a_66_6# DFFNEGX1_132/a_2_6# DFFNEGX1_132/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1949 out_state_main[3] DFFNEGX1_132/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1950 DFFNEGX1_132/a_23_6# INVX2_259/Y DFFNEGX1_132/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M1951 DFFNEGX1_132/a_23_6# DFFNEGX1_132/a_2_6# DFFNEGX1_132/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M1952 gnd DFFNEGX1_132/a_34_4# DFFNEGX1_132/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1953 vdd DFFNEGX1_132/a_34_4# DFFNEGX1_132/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M1954 DFFNEGX1_132/a_61_74# DFFNEGX1_132/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1955 DFFNEGX1_132/a_34_4# DFFNEGX1_132/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1956 DFFNEGX1_132/a_34_4# DFFNEGX1_132/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M1957 vdd out_state_main[3] DFFNEGX1_132/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M1958 gnd out_state_main[3] DFFNEGX1_132/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1959 DFFNEGX1_132/a_61_6# DFFNEGX1_132/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1960 DFFNEGX1_132/a_76_84# DFFNEGX1_132/a_2_6# DFFNEGX1_132/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M1961 out_state_main[3] DFFNEGX1_132/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M1962 vdd INVX2_259/Y DFFNEGX1_132/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M1963 DFFNEGX1_132/a_31_6# DFFNEGX1_132/a_2_6# DFFNEGX1_132/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1964 DFFNEGX1_132/a_66_6# INVX2_259/Y DFFNEGX1_132/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1965 DFFNEGX1_132/a_17_74# INVX2_117/A vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1966 DFFNEGX1_132/a_31_74# INVX2_259/Y DFFNEGX1_132/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1967 DFFNEGX1_132/a_17_6# INVX2_117/A gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1968 gnd MUX2X1_19/A MUX2X1_19/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M1969 MUX2X1_19/a_17_50# FAX1_1/YS vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1970 MUX2X1_19/Y OR2X1_3/Y MUX2X1_19/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M1971 MUX2X1_19/a_30_54# MUX2X1_19/a_2_10# MUX2X1_19/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M1972 MUX2X1_19/a_17_10# FAX1_1/YS gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1973 vdd OR2X1_3/Y MUX2X1_19/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M1974 MUX2X1_19/a_30_10# OR2X1_3/Y MUX2X1_19/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M1975 gnd OR2X1_3/Y MUX2X1_19/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M1976 vdd MUX2X1_19/A MUX2X1_19/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1977 MUX2X1_19/Y MUX2X1_19/a_2_10# MUX2X1_19/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1978 gnd out_global_score[31] AOI22X1_2/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M1979 INVX2_185/A INVX2_258/Y AOI22X1_2/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M1980 AOI22X1_2/a_11_6# XOR2X1_2/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1981 AOI22X1_2/a_2_54# INVX2_258/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M1982 AOI22X1_2/a_28_6# INVX2_255/Y INVX2_185/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1983 vdd XOR2X1_2/Y AOI22X1_2/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1984 INVX2_185/A INVX2_255/Y AOI22X1_2/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M1985 AOI22X1_2/a_2_54# out_global_score[31] INVX2_185/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1986 OAI21X1_8/B NOR2X1_61/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1987 NAND2X1_23/a_9_6# NOR2X1_61/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1988 vdd NOR2X1_63/B OAI21X1_8/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1989 OAI21X1_8/B NOR2X1_63/B NAND2X1_23/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1990 OAI21X1_33/C out_mines[9] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1991 NAND2X1_34/a_9_6# out_mines[9] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1992 vdd INVX2_221/Y OAI21X1_33/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1993 OAI21X1_33/C INVX2_221/Y NAND2X1_34/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1994 NOR2X1_57/B out_temp_data_in[1] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1995 NAND2X1_12/a_9_6# out_temp_data_in[1] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M1996 vdd out_temp_data_in[0] NOR2X1_57/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1997 NOR2X1_57/B out_temp_data_in[0] NAND2X1_12/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M1998 OAI21X1_48/B NOR2X1_64/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M1999 NAND2X1_45/a_9_6# NOR2X1_64/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2000 vdd NOR2X1_63/B OAI21X1_48/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2001 OAI21X1_48/B NOR2X1_63/B NAND2X1_45/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2002 OAI21X1_79/B INVX2_97/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M2003 NAND2X1_67/a_9_6# INVX2_97/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2004 vdd INVX2_65/Y OAI21X1_79/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2005 OAI21X1_79/B INVX2_65/Y NAND2X1_67/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2006 OAI21X1_59/B AND2X2_14/B vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M2007 NAND2X1_56/a_9_6# AND2X2_14/B gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2008 vdd INVX2_184/A OAI21X1_59/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2009 OAI21X1_59/B INVX2_184/A NAND2X1_56/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2010 NAND2X1_89/Y NOR2X1_47/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M2011 NAND2X1_89/a_9_6# NOR2X1_47/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2012 vdd BUFX2_21/Y NAND2X1_89/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2013 NAND2X1_89/Y BUFX2_21/Y NAND2X1_89/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2014 OAI21X1_91/C NOR2X1_35/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M2015 NAND2X1_78/a_9_6# NOR2X1_35/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2016 vdd BUFX2_20/Y OAI21X1_91/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2017 OAI21X1_91/C BUFX2_20/Y NAND2X1_78/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2018 gnd out_global_score[12] AOI22X1_21/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M2019 INVX2_204/A INVX2_258/Y AOI22X1_21/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2020 AOI22X1_21/a_11_6# HAX1_18/YS gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2021 AOI22X1_21/a_2_54# INVX2_258/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M2022 AOI22X1_21/a_28_6# OR2X1_11/B INVX2_204/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2023 vdd HAX1_18/YS AOI22X1_21/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2024 INVX2_204/A OR2X1_11/B AOI22X1_21/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M2025 AOI22X1_21/a_2_54# out_global_score[12] INVX2_204/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2026 gnd out_global_score[1] AOI22X1_32/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M2027 INVX2_215/A INVX2_258/Y AOI22X1_32/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2028 AOI22X1_32/a_11_6# HAX1_29/YS gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2029 AOI22X1_32/a_2_54# INVX2_258/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M2030 AOI22X1_32/a_28_6# INVX2_255/Y INVX2_215/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2031 vdd HAX1_29/YS AOI22X1_32/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2032 INVX2_215/A INVX2_255/Y AOI22X1_32/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M2033 AOI22X1_32/a_2_54# out_global_score[1] INVX2_215/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2034 gnd out_global_score[23] AOI22X1_10/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M2035 INVX2_193/A INVX2_257/Y AOI22X1_10/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2036 AOI22X1_10/a_11_6# HAX1_7/YS gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2037 AOI22X1_10/a_2_54# INVX2_257/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M2038 AOI22X1_10/a_28_6# INVX2_255/Y INVX2_193/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2039 vdd HAX1_7/YS AOI22X1_10/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2040 INVX2_193/A INVX2_255/Y AOI22X1_10/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M2041 AOI22X1_10/a_2_54# out_global_score[23] INVX2_193/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2042 gnd NOR2X1_88/Y AOI22X1_43/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M2043 NAND3X1_34/C out_mines[2] AOI22X1_43/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2044 AOI22X1_43/a_11_6# out_temp_cleared[2] gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2045 AOI22X1_43/a_2_54# out_mines[2] vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M2046 AOI22X1_43/a_28_6# INVX2_27/Y NAND3X1_34/C Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2047 vdd out_temp_cleared[2] AOI22X1_43/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2048 NAND3X1_34/C INVX2_27/Y AOI22X1_43/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M2049 AOI22X1_43/a_2_54# NOR2X1_88/Y NAND3X1_34/C vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2050 gnd INVX2_42/Y AOI22X1_54/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M2051 OAI22X1_34/C AOI22X1_54/B AOI22X1_54/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2052 AOI22X1_54/a_11_6# out_temp_data_in[2] gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2053 AOI22X1_54/a_2_54# AOI22X1_54/B vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M2054 AOI22X1_54/a_28_6# OAI21X1_1/B OAI22X1_34/C Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2055 vdd out_temp_data_in[2] AOI22X1_54/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2056 OAI22X1_34/C OAI21X1_1/B AOI22X1_54/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M2057 AOI22X1_54/a_2_54# INVX2_42/Y OAI22X1_34/C vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2058 gnd NOR2X1_113/Y AOI22X1_65/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M2059 AOI22X1_65/Y out_mines[19] AOI22X1_65/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2060 AOI22X1_65/a_11_6# NOR2X1_114/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2061 AOI22X1_65/a_2_54# out_mines[19] vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M2062 AOI22X1_65/a_28_6# out_mines[20] AOI22X1_65/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2063 vdd NOR2X1_114/Y AOI22X1_65/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2064 AOI22X1_65/Y out_mines[20] AOI22X1_65/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M2065 AOI22X1_65/a_2_54# NOR2X1_113/Y AOI22X1_65/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2066 gnd INVX2_123/Y AOI22X1_76/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M2067 NOR2X1_118/B INVX2_118/Y AOI22X1_76/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2068 AOI22X1_76/a_11_6# INVX2_126/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2069 AOI22X1_76/a_2_54# INVX2_118/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M2070 AOI22X1_76/a_28_6# OR2X1_16/Y NOR2X1_118/B Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2071 vdd INVX2_126/Y AOI22X1_76/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2072 NOR2X1_118/B OR2X1_16/Y AOI22X1_76/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M2073 AOI22X1_76/a_2_54# INVX2_123/Y NOR2X1_118/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2074 gnd BUFX2_25/Y OAI22X1_5/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M2075 OAI22X1_5/a_2_6# OAI22X1_5/C OAI22X1_5/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M2076 OAI22X1_5/Y INVX2_56/Y OAI22X1_5/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2077 OAI22X1_5/Y INVX2_90/Y OAI22X1_5/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M2078 OAI22X1_5/a_28_54# INVX2_56/Y OAI22X1_5/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2079 OAI22X1_5/a_9_54# BUFX2_25/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2080 OAI22X1_5/a_2_6# INVX2_90/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2081 vdd OAI22X1_5/C OAI22X1_5/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2082 INVX2_25/Y out_mines[18] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2083 INVX2_25/Y out_mines[18] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2084 INVX2_14/Y out_mines[12] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2085 INVX2_14/Y out_mines[12] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2086 INVX2_36/Y INVX2_36/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2087 INVX2_36/Y INVX2_36/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2088 INVX2_69/Y out_temp_decoded[12] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2089 INVX2_69/Y out_temp_decoded[12] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2090 INVX2_58/Y INVX2_58/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2091 INVX2_58/Y INVX2_58/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2092 INVX2_47/Y INVX2_47/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2093 INVX2_47/Y INVX2_47/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2094 HAX1_46/A MUX2X1_22/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2095 HAX1_46/A MUX2X1_22/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2096 INVX2_181/Y NOR2X1_62/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2097 INVX2_181/Y NOR2X1_62/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2098 INVX2_192/Y INVX2_192/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2099 INVX2_192/Y INVX2_192/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2100 gnd NOR2X1_4/A XNOR2X1_8/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2101 XNOR2X1_8/Y NOR2X1_4/A XNOR2X1_8/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2102 XNOR2X1_8/a_12_41# FAX1_0/YS gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2103 XNOR2X1_8/a_18_54# XNOR2X1_8/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2104 XNOR2X1_8/a_35_6# XNOR2X1_8/a_2_6# XNOR2X1_8/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2105 XNOR2X1_8/a_18_6# XNOR2X1_8/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2106 vdd NOR2X1_4/A XNOR2X1_8/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2107 vdd FAX1_0/YS XNOR2X1_8/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2108 XNOR2X1_8/Y XNOR2X1_8/a_2_6# XNOR2X1_8/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2109 XNOR2X1_8/a_35_54# NOR2X1_4/A XNOR2X1_8/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2110 XNOR2X1_8/a_12_41# FAX1_0/YS vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2111 gnd FAX1_0/YS XNOR2X1_8/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2112 DFFNEGX1_32/a_76_6# BUFX2_15/Y DFFNEGX1_32/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2113 gnd BUFX2_15/Y DFFNEGX1_32/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2114 DFFNEGX1_32/a_66_6# DFFNEGX1_32/a_2_6# DFFNEGX1_32/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2115 out_temp_mine_cnt[1] DFFNEGX1_32/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2116 DFFNEGX1_32/a_23_6# BUFX2_15/Y DFFNEGX1_32/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2117 DFFNEGX1_32/a_23_6# DFFNEGX1_32/a_2_6# DFFNEGX1_32/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2118 gnd DFFNEGX1_32/a_34_4# DFFNEGX1_32/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2119 vdd DFFNEGX1_32/a_34_4# DFFNEGX1_32/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2120 DFFNEGX1_32/a_61_74# DFFNEGX1_32/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2121 DFFNEGX1_32/a_34_4# DFFNEGX1_32/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2122 DFFNEGX1_32/a_34_4# DFFNEGX1_32/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2123 vdd out_temp_mine_cnt[1] DFFNEGX1_32/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2124 gnd out_temp_mine_cnt[1] DFFNEGX1_32/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2125 DFFNEGX1_32/a_61_6# DFFNEGX1_32/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2126 DFFNEGX1_32/a_76_84# DFFNEGX1_32/a_2_6# DFFNEGX1_32/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2127 out_temp_mine_cnt[1] DFFNEGX1_32/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2128 vdd BUFX2_15/Y DFFNEGX1_32/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2129 DFFNEGX1_32/a_31_6# DFFNEGX1_32/a_2_6# DFFNEGX1_32/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2130 DFFNEGX1_32/a_66_6# BUFX2_15/Y DFFNEGX1_32/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2131 DFFNEGX1_32/a_17_74# AND2X2_12/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2132 DFFNEGX1_32/a_31_74# BUFX2_15/Y DFFNEGX1_32/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2133 DFFNEGX1_32/a_17_6# AND2X2_12/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2134 DFFNEGX1_10/a_76_6# BUFX2_17/Y DFFNEGX1_10/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2135 gnd BUFX2_17/Y DFFNEGX1_10/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2136 DFFNEGX1_10/a_66_6# DFFNEGX1_10/a_2_6# DFFNEGX1_10/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2137 out_mines[1] DFFNEGX1_10/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2138 DFFNEGX1_10/a_23_6# BUFX2_17/Y DFFNEGX1_10/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2139 DFFNEGX1_10/a_23_6# DFFNEGX1_10/a_2_6# DFFNEGX1_10/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2140 gnd DFFNEGX1_10/a_34_4# DFFNEGX1_10/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2141 vdd DFFNEGX1_10/a_34_4# DFFNEGX1_10/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2142 DFFNEGX1_10/a_61_74# DFFNEGX1_10/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2143 DFFNEGX1_10/a_34_4# DFFNEGX1_10/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2144 DFFNEGX1_10/a_34_4# DFFNEGX1_10/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2145 vdd out_mines[1] DFFNEGX1_10/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2146 gnd out_mines[1] DFFNEGX1_10/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2147 DFFNEGX1_10/a_61_6# DFFNEGX1_10/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2148 DFFNEGX1_10/a_76_84# DFFNEGX1_10/a_2_6# DFFNEGX1_10/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2149 out_mines[1] DFFNEGX1_10/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2150 vdd BUFX2_17/Y DFFNEGX1_10/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2151 DFFNEGX1_10/a_31_6# DFFNEGX1_10/a_2_6# DFFNEGX1_10/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2152 DFFNEGX1_10/a_66_6# BUFX2_17/Y DFFNEGX1_10/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2153 DFFNEGX1_10/a_17_74# OAI21X1_49/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2154 DFFNEGX1_10/a_31_74# BUFX2_17/Y DFFNEGX1_10/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2155 DFFNEGX1_10/a_17_6# OAI21X1_49/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2156 DFFNEGX1_21/a_76_6# BUFX2_16/Y DFFNEGX1_21/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2157 gnd BUFX2_16/Y DFFNEGX1_21/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2158 DFFNEGX1_21/a_66_6# DFFNEGX1_21/a_2_6# DFFNEGX1_21/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2159 out_mines[20] DFFNEGX1_21/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2160 DFFNEGX1_21/a_23_6# BUFX2_16/Y DFFNEGX1_21/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2161 DFFNEGX1_21/a_23_6# DFFNEGX1_21/a_2_6# DFFNEGX1_21/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2162 gnd DFFNEGX1_21/a_34_4# DFFNEGX1_21/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2163 vdd DFFNEGX1_21/a_34_4# DFFNEGX1_21/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2164 DFFNEGX1_21/a_61_74# DFFNEGX1_21/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2165 DFFNEGX1_21/a_34_4# DFFNEGX1_21/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2166 DFFNEGX1_21/a_34_4# DFFNEGX1_21/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2167 vdd out_mines[20] DFFNEGX1_21/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2168 gnd out_mines[20] DFFNEGX1_21/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2169 DFFNEGX1_21/a_61_6# DFFNEGX1_21/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2170 DFFNEGX1_21/a_76_84# DFFNEGX1_21/a_2_6# DFFNEGX1_21/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2171 out_mines[20] DFFNEGX1_21/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2172 vdd BUFX2_16/Y DFFNEGX1_21/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2173 DFFNEGX1_21/a_31_6# DFFNEGX1_21/a_2_6# DFFNEGX1_21/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2174 DFFNEGX1_21/a_66_6# BUFX2_16/Y DFFNEGX1_21/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2175 DFFNEGX1_21/a_17_74# OAI21X1_11/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2176 DFFNEGX1_21/a_31_74# BUFX2_16/Y DFFNEGX1_21/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2177 DFFNEGX1_21/a_17_6# OAI21X1_11/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2178 DFFNEGX1_43/a_76_6# BUFX2_14/Y DFFNEGX1_43/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2179 gnd BUFX2_14/Y DFFNEGX1_43/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2180 DFFNEGX1_43/a_66_6# DFFNEGX1_43/a_2_6# DFFNEGX1_43/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2181 out_temp_decoded[23] DFFNEGX1_43/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2182 DFFNEGX1_43/a_23_6# BUFX2_14/Y DFFNEGX1_43/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2183 DFFNEGX1_43/a_23_6# DFFNEGX1_43/a_2_6# DFFNEGX1_43/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2184 gnd DFFNEGX1_43/a_34_4# DFFNEGX1_43/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2185 vdd DFFNEGX1_43/a_34_4# DFFNEGX1_43/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2186 DFFNEGX1_43/a_61_74# DFFNEGX1_43/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2187 DFFNEGX1_43/a_34_4# DFFNEGX1_43/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2188 DFFNEGX1_43/a_34_4# DFFNEGX1_43/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2189 vdd out_temp_decoded[23] DFFNEGX1_43/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2190 gnd out_temp_decoded[23] DFFNEGX1_43/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2191 DFFNEGX1_43/a_61_6# DFFNEGX1_43/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2192 DFFNEGX1_43/a_76_84# DFFNEGX1_43/a_2_6# DFFNEGX1_43/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2193 out_temp_decoded[23] DFFNEGX1_43/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2194 vdd BUFX2_14/Y DFFNEGX1_43/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2195 DFFNEGX1_43/a_31_6# DFFNEGX1_43/a_2_6# DFFNEGX1_43/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2196 DFFNEGX1_43/a_66_6# BUFX2_14/Y DFFNEGX1_43/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2197 DFFNEGX1_43/a_17_74# OAI21X1_105/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2198 DFFNEGX1_43/a_31_74# BUFX2_14/Y DFFNEGX1_43/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2199 DFFNEGX1_43/a_17_6# OAI21X1_105/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2200 DFFNEGX1_54/a_76_6# BUFX2_13/Y DFFNEGX1_54/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2201 gnd BUFX2_13/Y DFFNEGX1_54/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2202 DFFNEGX1_54/a_66_6# DFFNEGX1_54/a_2_6# DFFNEGX1_54/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2203 out_temp_decoded[12] DFFNEGX1_54/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2204 DFFNEGX1_54/a_23_6# BUFX2_13/Y DFFNEGX1_54/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2205 DFFNEGX1_54/a_23_6# DFFNEGX1_54/a_2_6# DFFNEGX1_54/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2206 gnd DFFNEGX1_54/a_34_4# DFFNEGX1_54/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2207 vdd DFFNEGX1_54/a_34_4# DFFNEGX1_54/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2208 DFFNEGX1_54/a_61_74# DFFNEGX1_54/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2209 DFFNEGX1_54/a_34_4# DFFNEGX1_54/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2210 DFFNEGX1_54/a_34_4# DFFNEGX1_54/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2211 vdd out_temp_decoded[12] DFFNEGX1_54/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2212 gnd out_temp_decoded[12] DFFNEGX1_54/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2213 DFFNEGX1_54/a_61_6# DFFNEGX1_54/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2214 DFFNEGX1_54/a_76_84# DFFNEGX1_54/a_2_6# DFFNEGX1_54/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2215 out_temp_decoded[12] DFFNEGX1_54/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2216 vdd BUFX2_13/Y DFFNEGX1_54/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2217 DFFNEGX1_54/a_31_6# DFFNEGX1_54/a_2_6# DFFNEGX1_54/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2218 DFFNEGX1_54/a_66_6# BUFX2_13/Y DFFNEGX1_54/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2219 DFFNEGX1_54/a_17_74# OAI21X1_94/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2220 DFFNEGX1_54/a_31_74# BUFX2_13/Y DFFNEGX1_54/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2221 DFFNEGX1_54/a_17_6# OAI21X1_94/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2222 DFFNEGX1_76/a_76_6# BUFX2_12/Y DFFNEGX1_76/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2223 gnd BUFX2_12/Y DFFNEGX1_76/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2224 DFFNEGX1_76/a_66_6# DFFNEGX1_76/a_2_6# DFFNEGX1_76/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2225 out_temp_cleared[15] DFFNEGX1_76/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2226 DFFNEGX1_76/a_23_6# BUFX2_12/Y DFFNEGX1_76/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2227 DFFNEGX1_76/a_23_6# DFFNEGX1_76/a_2_6# DFFNEGX1_76/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2228 gnd DFFNEGX1_76/a_34_4# DFFNEGX1_76/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2229 vdd DFFNEGX1_76/a_34_4# DFFNEGX1_76/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2230 DFFNEGX1_76/a_61_74# DFFNEGX1_76/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2231 DFFNEGX1_76/a_34_4# DFFNEGX1_76/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2232 DFFNEGX1_76/a_34_4# DFFNEGX1_76/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2233 vdd out_temp_cleared[15] DFFNEGX1_76/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2234 gnd out_temp_cleared[15] DFFNEGX1_76/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2235 DFFNEGX1_76/a_61_6# DFFNEGX1_76/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2236 DFFNEGX1_76/a_76_84# DFFNEGX1_76/a_2_6# DFFNEGX1_76/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2237 out_temp_cleared[15] DFFNEGX1_76/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2238 vdd BUFX2_12/Y DFFNEGX1_76/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2239 DFFNEGX1_76/a_31_6# DFFNEGX1_76/a_2_6# DFFNEGX1_76/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2240 DFFNEGX1_76/a_66_6# BUFX2_12/Y DFFNEGX1_76/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2241 DFFNEGX1_76/a_17_74# OAI22X1_13/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2242 DFFNEGX1_76/a_31_74# BUFX2_12/Y DFFNEGX1_76/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2243 DFFNEGX1_76/a_17_6# OAI22X1_13/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2244 DFFNEGX1_65/a_76_6# BUFX2_13/Y DFFNEGX1_65/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2245 gnd BUFX2_13/Y DFFNEGX1_65/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2246 DFFNEGX1_65/a_66_6# DFFNEGX1_65/a_2_6# DFFNEGX1_65/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2247 out_temp_decoded[1] DFFNEGX1_65/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2248 DFFNEGX1_65/a_23_6# BUFX2_13/Y DFFNEGX1_65/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2249 DFFNEGX1_65/a_23_6# DFFNEGX1_65/a_2_6# DFFNEGX1_65/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2250 gnd DFFNEGX1_65/a_34_4# DFFNEGX1_65/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2251 vdd DFFNEGX1_65/a_34_4# DFFNEGX1_65/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2252 DFFNEGX1_65/a_61_74# DFFNEGX1_65/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2253 DFFNEGX1_65/a_34_4# DFFNEGX1_65/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2254 DFFNEGX1_65/a_34_4# DFFNEGX1_65/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2255 vdd out_temp_decoded[1] DFFNEGX1_65/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2256 gnd out_temp_decoded[1] DFFNEGX1_65/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2257 DFFNEGX1_65/a_61_6# DFFNEGX1_65/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2258 DFFNEGX1_65/a_76_84# DFFNEGX1_65/a_2_6# DFFNEGX1_65/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2259 out_temp_decoded[1] DFFNEGX1_65/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2260 vdd BUFX2_13/Y DFFNEGX1_65/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2261 DFFNEGX1_65/a_31_6# DFFNEGX1_65/a_2_6# DFFNEGX1_65/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2262 DFFNEGX1_65/a_66_6# BUFX2_13/Y DFFNEGX1_65/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2263 DFFNEGX1_65/a_17_74# OAI21X1_83/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2264 DFFNEGX1_65/a_31_74# BUFX2_13/Y DFFNEGX1_65/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2265 DFFNEGX1_65/a_17_6# OAI21X1_83/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2266 DFFNEGX1_98/a_76_6# BUFX2_10/Y DFFNEGX1_98/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2267 gnd BUFX2_10/Y DFFNEGX1_98/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2268 DFFNEGX1_98/a_66_6# DFFNEGX1_98/a_2_6# DFFNEGX1_98/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2269 out_global_score[4] DFFNEGX1_98/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2270 DFFNEGX1_98/a_23_6# BUFX2_10/Y DFFNEGX1_98/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2271 DFFNEGX1_98/a_23_6# DFFNEGX1_98/a_2_6# DFFNEGX1_98/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2272 gnd DFFNEGX1_98/a_34_4# DFFNEGX1_98/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2273 vdd DFFNEGX1_98/a_34_4# DFFNEGX1_98/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2274 DFFNEGX1_98/a_61_74# DFFNEGX1_98/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2275 DFFNEGX1_98/a_34_4# DFFNEGX1_98/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2276 DFFNEGX1_98/a_34_4# DFFNEGX1_98/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2277 vdd out_global_score[4] DFFNEGX1_98/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2278 gnd out_global_score[4] DFFNEGX1_98/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2279 DFFNEGX1_98/a_61_6# DFFNEGX1_98/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2280 DFFNEGX1_98/a_76_84# DFFNEGX1_98/a_2_6# DFFNEGX1_98/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2281 out_global_score[4] DFFNEGX1_98/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2282 vdd BUFX2_10/Y DFFNEGX1_98/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2283 DFFNEGX1_98/a_31_6# DFFNEGX1_98/a_2_6# DFFNEGX1_98/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2284 DFFNEGX1_98/a_66_6# BUFX2_10/Y DFFNEGX1_98/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2285 DFFNEGX1_98/a_17_74# INVX2_212/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2286 DFFNEGX1_98/a_31_74# BUFX2_10/Y DFFNEGX1_98/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2287 DFFNEGX1_98/a_17_6# INVX2_212/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2288 DFFNEGX1_87/a_76_6# BUFX2_11/Y DFFNEGX1_87/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2289 gnd BUFX2_11/Y DFFNEGX1_87/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2290 DFFNEGX1_87/a_66_6# DFFNEGX1_87/a_2_6# DFFNEGX1_87/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2291 out_temp_cleared[4] DFFNEGX1_87/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2292 DFFNEGX1_87/a_23_6# BUFX2_11/Y DFFNEGX1_87/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2293 DFFNEGX1_87/a_23_6# DFFNEGX1_87/a_2_6# DFFNEGX1_87/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2294 gnd DFFNEGX1_87/a_34_4# DFFNEGX1_87/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2295 vdd DFFNEGX1_87/a_34_4# DFFNEGX1_87/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2296 DFFNEGX1_87/a_61_74# DFFNEGX1_87/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2297 DFFNEGX1_87/a_34_4# DFFNEGX1_87/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2298 DFFNEGX1_87/a_34_4# DFFNEGX1_87/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2299 vdd out_temp_cleared[4] DFFNEGX1_87/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2300 gnd out_temp_cleared[4] DFFNEGX1_87/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2301 DFFNEGX1_87/a_61_6# DFFNEGX1_87/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2302 DFFNEGX1_87/a_76_84# DFFNEGX1_87/a_2_6# DFFNEGX1_87/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2303 out_temp_cleared[4] DFFNEGX1_87/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2304 vdd BUFX2_11/Y DFFNEGX1_87/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2305 DFFNEGX1_87/a_31_6# DFFNEGX1_87/a_2_6# DFFNEGX1_87/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2306 DFFNEGX1_87/a_66_6# BUFX2_11/Y DFFNEGX1_87/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2307 DFFNEGX1_87/a_17_74# OAI22X1_24/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2308 DFFNEGX1_87/a_31_74# BUFX2_11/Y DFFNEGX1_87/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2309 DFFNEGX1_87/a_17_6# OAI22X1_24/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2310 AND2X2_8/a_2_6# AND2X2_8/A vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M2311 AND2X2_8/a_9_6# AND2X2_8/A AND2X2_8/a_2_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=100p ps=50u
M2312 BUFX2_19/A AND2X2_8/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2313 BUFX2_19/A AND2X2_8/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2314 vdd AND2X2_8/B AND2X2_8/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2315 gnd AND2X2_8/B AND2X2_8/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2316 DFFNEGX1_111/a_76_6# BUFX2_9/Y DFFNEGX1_111/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2317 gnd BUFX2_9/Y DFFNEGX1_111/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2318 DFFNEGX1_111/a_66_6# DFFNEGX1_111/a_2_6# DFFNEGX1_111/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2319 out_global_score[17] DFFNEGX1_111/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2320 DFFNEGX1_111/a_23_6# BUFX2_9/Y DFFNEGX1_111/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2321 DFFNEGX1_111/a_23_6# DFFNEGX1_111/a_2_6# DFFNEGX1_111/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2322 gnd DFFNEGX1_111/a_34_4# DFFNEGX1_111/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2323 vdd DFFNEGX1_111/a_34_4# DFFNEGX1_111/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2324 DFFNEGX1_111/a_61_74# DFFNEGX1_111/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2325 DFFNEGX1_111/a_34_4# DFFNEGX1_111/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2326 DFFNEGX1_111/a_34_4# DFFNEGX1_111/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2327 vdd out_global_score[17] DFFNEGX1_111/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2328 gnd out_global_score[17] DFFNEGX1_111/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2329 DFFNEGX1_111/a_61_6# DFFNEGX1_111/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2330 DFFNEGX1_111/a_76_84# DFFNEGX1_111/a_2_6# DFFNEGX1_111/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2331 out_global_score[17] DFFNEGX1_111/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2332 vdd BUFX2_9/Y DFFNEGX1_111/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2333 DFFNEGX1_111/a_31_6# DFFNEGX1_111/a_2_6# DFFNEGX1_111/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2334 DFFNEGX1_111/a_66_6# BUFX2_9/Y DFFNEGX1_111/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2335 DFFNEGX1_111/a_17_74# INVX2_199/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2336 DFFNEGX1_111/a_31_74# BUFX2_9/Y DFFNEGX1_111/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2337 DFFNEGX1_111/a_17_6# INVX2_199/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2338 DFFNEGX1_100/a_76_6# BUFX2_10/Y DFFNEGX1_100/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2339 gnd BUFX2_10/Y DFFNEGX1_100/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2340 DFFNEGX1_100/a_66_6# DFFNEGX1_100/a_2_6# DFFNEGX1_100/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2341 out_global_score[6] DFFNEGX1_100/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2342 DFFNEGX1_100/a_23_6# BUFX2_10/Y DFFNEGX1_100/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2343 DFFNEGX1_100/a_23_6# DFFNEGX1_100/a_2_6# DFFNEGX1_100/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2344 gnd DFFNEGX1_100/a_34_4# DFFNEGX1_100/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2345 vdd DFFNEGX1_100/a_34_4# DFFNEGX1_100/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2346 DFFNEGX1_100/a_61_74# DFFNEGX1_100/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2347 DFFNEGX1_100/a_34_4# DFFNEGX1_100/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2348 DFFNEGX1_100/a_34_4# DFFNEGX1_100/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2349 vdd out_global_score[6] DFFNEGX1_100/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2350 gnd out_global_score[6] DFFNEGX1_100/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2351 DFFNEGX1_100/a_61_6# DFFNEGX1_100/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2352 DFFNEGX1_100/a_76_84# DFFNEGX1_100/a_2_6# DFFNEGX1_100/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2353 out_global_score[6] DFFNEGX1_100/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2354 vdd BUFX2_10/Y DFFNEGX1_100/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2355 DFFNEGX1_100/a_31_6# DFFNEGX1_100/a_2_6# DFFNEGX1_100/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2356 DFFNEGX1_100/a_66_6# BUFX2_10/Y DFFNEGX1_100/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2357 DFFNEGX1_100/a_17_74# INVX2_210/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2358 DFFNEGX1_100/a_31_74# BUFX2_10/Y DFFNEGX1_100/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2359 DFFNEGX1_100/a_17_6# INVX2_210/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2360 DFFNEGX1_133/a_76_6# BUFX2_5/Y DFFNEGX1_133/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2361 gnd BUFX2_5/Y DFFNEGX1_133/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2362 DFFNEGX1_133/a_66_6# DFFNEGX1_133/a_2_6# DFFNEGX1_133/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2363 INVX2_119/A DFFNEGX1_133/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2364 DFFNEGX1_133/a_23_6# BUFX2_5/Y DFFNEGX1_133/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2365 DFFNEGX1_133/a_23_6# DFFNEGX1_133/a_2_6# DFFNEGX1_133/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2366 gnd DFFNEGX1_133/a_34_4# DFFNEGX1_133/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2367 vdd DFFNEGX1_133/a_34_4# DFFNEGX1_133/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2368 DFFNEGX1_133/a_61_74# DFFNEGX1_133/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2369 DFFNEGX1_133/a_34_4# DFFNEGX1_133/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2370 DFFNEGX1_133/a_34_4# DFFNEGX1_133/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2371 vdd INVX2_119/A DFFNEGX1_133/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2372 gnd INVX2_119/A DFFNEGX1_133/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2373 DFFNEGX1_133/a_61_6# DFFNEGX1_133/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2374 DFFNEGX1_133/a_76_84# DFFNEGX1_133/a_2_6# DFFNEGX1_133/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2375 INVX2_119/A DFFNEGX1_133/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2376 vdd BUFX2_5/Y DFFNEGX1_133/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2377 DFFNEGX1_133/a_31_6# DFFNEGX1_133/a_2_6# DFFNEGX1_133/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2378 DFFNEGX1_133/a_66_6# BUFX2_5/Y DFFNEGX1_133/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2379 DFFNEGX1_133/a_17_74# NOR2X1_118/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2380 DFFNEGX1_133/a_31_74# BUFX2_5/Y DFFNEGX1_133/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2381 DFFNEGX1_133/a_17_6# NOR2X1_118/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2382 DFFNEGX1_122/a_76_6# BUFX2_5/Y DFFNEGX1_122/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2383 gnd BUFX2_5/Y DFFNEGX1_122/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2384 DFFNEGX1_122/a_66_6# DFFNEGX1_122/a_2_6# DFFNEGX1_122/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2385 out_global_score[28] DFFNEGX1_122/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2386 DFFNEGX1_122/a_23_6# BUFX2_5/Y DFFNEGX1_122/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2387 DFFNEGX1_122/a_23_6# DFFNEGX1_122/a_2_6# DFFNEGX1_122/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2388 gnd DFFNEGX1_122/a_34_4# DFFNEGX1_122/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2389 vdd DFFNEGX1_122/a_34_4# DFFNEGX1_122/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2390 DFFNEGX1_122/a_61_74# DFFNEGX1_122/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2391 DFFNEGX1_122/a_34_4# DFFNEGX1_122/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2392 DFFNEGX1_122/a_34_4# DFFNEGX1_122/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2393 vdd out_global_score[28] DFFNEGX1_122/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2394 gnd out_global_score[28] DFFNEGX1_122/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2395 DFFNEGX1_122/a_61_6# DFFNEGX1_122/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2396 DFFNEGX1_122/a_76_84# DFFNEGX1_122/a_2_6# DFFNEGX1_122/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2397 out_global_score[28] DFFNEGX1_122/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2398 vdd BUFX2_5/Y DFFNEGX1_122/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2399 DFFNEGX1_122/a_31_6# DFFNEGX1_122/a_2_6# DFFNEGX1_122/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2400 DFFNEGX1_122/a_66_6# BUFX2_5/Y DFFNEGX1_122/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2401 DFFNEGX1_122/a_17_74# INVX2_188/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2402 DFFNEGX1_122/a_31_74# BUFX2_5/Y DFFNEGX1_122/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2403 DFFNEGX1_122/a_17_6# INVX2_188/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2404 gnd out_global_score[30] AOI22X1_3/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M2405 INVX2_186/A INVX2_257/Y AOI22X1_3/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2406 AOI22X1_3/a_11_6# HAX1_0/YS gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2407 AOI22X1_3/a_2_54# INVX2_257/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M2408 AOI22X1_3/a_28_6# INVX2_255/Y INVX2_186/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2409 vdd HAX1_0/YS AOI22X1_3/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2410 INVX2_186/A INVX2_255/Y AOI22X1_3/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M2411 AOI22X1_3/a_2_54# out_global_score[30] INVX2_186/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2412 gnd NOR2X1_116/Y OAI21X1_160/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M2413 vdd AND2X2_17/A OAI21X1_160/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M2414 OAI21X1_160/Y AND2X2_17/A OAI21X1_160/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2415 OAI21X1_160/Y INVX2_117/Y OAI21X1_160/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2416 OAI21X1_160/a_9_54# NOR2X1_116/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2417 OAI21X1_160/a_2_6# INVX2_117/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2418 NOR2X1_7/A XOR2X1_5/A vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M2419 NAND2X1_13/a_9_6# XOR2X1_5/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2420 vdd FAX1_4/YC NOR2X1_7/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2421 NOR2X1_7/A FAX1_4/YC NAND2X1_13/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2422 OAI21X1_17/C out_mines[17] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M2423 NAND2X1_24/a_9_6# out_mines[17] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2424 vdd INVX2_220/Y OAI21X1_17/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2425 OAI21X1_17/C INVX2_220/Y NAND2X1_24/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2426 OAI21X1_49/C out_mines[1] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M2427 NAND2X1_46/a_9_6# out_mines[1] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2428 vdd INVX2_222/Y OAI21X1_49/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2429 OAI21X1_49/C INVX2_222/Y NAND2X1_46/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2430 OAI21X1_35/C out_mines[8] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M2431 NAND2X1_35/a_9_6# out_mines[8] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2432 vdd INVX2_225/Y OAI21X1_35/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2433 OAI21X1_35/C INVX2_225/Y NAND2X1_35/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2434 OAI21X1_80/B OAI22X1_2/B vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M2435 NAND2X1_68/a_9_6# OAI22X1_2/B gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2436 vdd INVX2_79/Y OAI21X1_80/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2437 OAI21X1_80/B INVX2_79/Y NAND2X1_68/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2438 OAI21X1_60/C out_n_nearby[0] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M2439 NAND2X1_57/a_9_6# out_n_nearby[0] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2440 vdd AOI21X1_2/A OAI21X1_60/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2441 OAI21X1_60/C AOI21X1_2/A NAND2X1_57/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2442 OAI21X1_92/C NOR2X1_58/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M2443 NAND2X1_79/a_9_6# NOR2X1_58/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2444 vdd BUFX2_20/Y OAI21X1_92/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2445 OAI21X1_92/C BUFX2_20/Y NAND2X1_79/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2446 gnd out_global_score[11] AOI22X1_22/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M2447 INVX2_205/A INVX2_258/Y AOI22X1_22/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2448 AOI22X1_22/a_11_6# HAX1_19/YS gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2449 AOI22X1_22/a_2_54# INVX2_258/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M2450 AOI22X1_22/a_28_6# OR2X1_11/B INVX2_205/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2451 vdd HAX1_19/YS AOI22X1_22/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2452 INVX2_205/A OR2X1_11/B AOI22X1_22/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M2453 AOI22X1_22/a_2_54# out_global_score[11] INVX2_205/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2454 gnd out_global_score[0] AOI22X1_33/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M2455 INVX2_216/A INVX2_258/Y AOI22X1_33/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2456 AOI22X1_33/a_11_6# INVX2_114/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2457 AOI22X1_33/a_2_54# INVX2_258/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M2458 AOI22X1_33/a_28_6# OR2X1_11/B INVX2_216/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2459 vdd INVX2_114/Y AOI22X1_33/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2460 INVX2_216/A OR2X1_11/B AOI22X1_33/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M2461 AOI22X1_33/a_2_54# out_global_score[0] INVX2_216/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2462 gnd out_global_score[22] AOI22X1_11/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M2463 INVX2_194/A INVX2_257/Y AOI22X1_11/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2464 AOI22X1_11/a_11_6# HAX1_8/YS gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2465 AOI22X1_11/a_2_54# INVX2_257/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M2466 AOI22X1_11/a_28_6# INVX2_255/Y INVX2_194/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2467 vdd HAX1_8/YS AOI22X1_11/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2468 INVX2_194/A INVX2_255/Y AOI22X1_11/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M2469 AOI22X1_11/a_2_54# out_global_score[22] INVX2_194/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2470 gnd out_temp_cleared[12] AOI22X1_44/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M2471 NAND3X1_39/B INVX2_13/Y AOI22X1_44/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2472 AOI22X1_44/a_11_6# NOR2X1_93/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2473 AOI22X1_44/a_2_54# INVX2_13/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M2474 AOI22X1_44/a_28_6# out_mines[12] NAND3X1_39/B Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2475 vdd NOR2X1_93/Y AOI22X1_44/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2476 NAND3X1_39/B out_mines[12] AOI22X1_44/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M2477 AOI22X1_44/a_2_54# out_temp_cleared[12] NAND3X1_39/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2478 gnd INVX2_41/Y AOI22X1_55/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M2479 AOI22X1_55/Y INVX2_251/Y AOI22X1_55/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2480 AOI22X1_55/a_11_6# OAI22X1_35/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2481 AOI22X1_55/a_2_54# INVX2_251/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M2482 AOI22X1_55/a_28_6# out_mines[13] AOI22X1_55/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2483 vdd OAI22X1_35/Y AOI22X1_55/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2484 AOI22X1_55/Y out_mines[13] AOI22X1_55/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M2485 AOI22X1_55/a_2_54# INVX2_41/Y AOI22X1_55/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2486 gnd NOR2X1_111/Y AOI22X1_66/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M2487 AND2X2_16/B INVX2_33/A AOI22X1_66/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2488 AOI22X1_66/a_11_6# NOR2X1_112/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2489 AOI22X1_66/a_2_54# INVX2_33/A vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M2490 AOI22X1_66/a_28_6# AOI22X1_66/D AND2X2_16/B Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2491 vdd NOR2X1_112/Y AOI22X1_66/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2492 AND2X2_16/B AOI22X1_66/D AOI22X1_66/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M2493 AOI22X1_66/a_2_54# NOR2X1_111/Y AND2X2_16/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2494 gnd out_state_main[0] AOI22X1_77/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M2495 INVX2_126/A out_state_main[2] AOI22X1_77/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2496 AOI22X1_77/a_11_6# INVX2_125/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2497 AOI22X1_77/a_2_54# out_state_main[2] vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M2498 AOI22X1_77/a_28_6# NOR2X1_121/Y INVX2_126/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2499 vdd INVX2_125/Y AOI22X1_77/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2500 INVX2_126/A NOR2X1_121/Y AOI22X1_77/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M2501 AOI22X1_77/a_2_54# out_state_main[0] INVX2_126/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2502 gnd BUFX2_25/Y OAI22X1_6/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M2503 OAI22X1_6/a_2_6# OR2X1_11/A OAI22X1_6/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M2504 OAI22X1_6/Y INVX2_57/Y OAI22X1_6/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2505 OAI22X1_6/Y INVX2_91/Y OAI22X1_6/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M2506 OAI22X1_6/a_28_54# INVX2_57/Y OAI22X1_6/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2507 OAI22X1_6/a_9_54# BUFX2_25/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2508 OAI22X1_6/a_2_6# INVX2_91/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2509 vdd OR2X1_11/A OAI22X1_6/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2510 INVX2_26/Y out_mines[11] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2511 INVX2_26/Y out_mines[11] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2512 INVX2_15/Y out_mines[8] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2513 INVX2_15/Y out_mines[8] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2514 INVX2_59/Y out_temp_decoded[21] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2515 INVX2_59/Y out_temp_decoded[21] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2516 INVX2_48/Y INVX2_48/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2517 INVX2_48/Y INVX2_48/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2518 INVX2_37/Y INVX2_37/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2519 INVX2_37/Y INVX2_37/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2520 NOR2X1_3/A MUX2X1_14/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2521 NOR2X1_3/A MUX2X1_14/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2522 MUX2X1_27/B XNOR2X1_3/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2523 MUX2X1_27/B XNOR2X1_3/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2524 NAND3X1_7/C NAND3X1_9/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2525 NAND3X1_7/C NAND3X1_9/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2526 INVX2_193/Y INVX2_193/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2527 INVX2_193/Y INVX2_193/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2528 gnd MUX2X1_8/Y XNOR2X1_9/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2529 XNOR2X1_9/Y MUX2X1_8/Y XNOR2X1_9/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2530 XNOR2X1_9/a_12_41# NOR2X1_4/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2531 XNOR2X1_9/a_18_54# XNOR2X1_9/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2532 XNOR2X1_9/a_35_6# XNOR2X1_9/a_2_6# XNOR2X1_9/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2533 XNOR2X1_9/a_18_6# XNOR2X1_9/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2534 vdd MUX2X1_8/Y XNOR2X1_9/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2535 vdd NOR2X1_4/Y XNOR2X1_9/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2536 XNOR2X1_9/Y XNOR2X1_9/a_2_6# XNOR2X1_9/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M2537 XNOR2X1_9/a_35_54# MUX2X1_8/Y XNOR2X1_9/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2538 XNOR2X1_9/a_12_41# NOR2X1_4/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2539 gnd NOR2X1_4/Y XNOR2X1_9/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2540 DFFNEGX1_33/a_76_6# BUFX2_15/Y DFFNEGX1_33/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2541 gnd BUFX2_15/Y DFFNEGX1_33/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2542 DFFNEGX1_33/a_66_6# DFFNEGX1_33/a_2_6# DFFNEGX1_33/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2543 out_temp_mine_cnt[2] DFFNEGX1_33/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2544 DFFNEGX1_33/a_23_6# BUFX2_15/Y DFFNEGX1_33/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2545 DFFNEGX1_33/a_23_6# DFFNEGX1_33/a_2_6# DFFNEGX1_33/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2546 gnd DFFNEGX1_33/a_34_4# DFFNEGX1_33/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2547 vdd DFFNEGX1_33/a_34_4# DFFNEGX1_33/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2548 DFFNEGX1_33/a_61_74# DFFNEGX1_33/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2549 DFFNEGX1_33/a_34_4# DFFNEGX1_33/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2550 DFFNEGX1_33/a_34_4# DFFNEGX1_33/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2551 vdd out_temp_mine_cnt[2] DFFNEGX1_33/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2552 gnd out_temp_mine_cnt[2] DFFNEGX1_33/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2553 DFFNEGX1_33/a_61_6# DFFNEGX1_33/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2554 DFFNEGX1_33/a_76_84# DFFNEGX1_33/a_2_6# DFFNEGX1_33/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2555 out_temp_mine_cnt[2] DFFNEGX1_33/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2556 vdd BUFX2_15/Y DFFNEGX1_33/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2557 DFFNEGX1_33/a_31_6# DFFNEGX1_33/a_2_6# DFFNEGX1_33/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2558 DFFNEGX1_33/a_66_6# BUFX2_15/Y DFFNEGX1_33/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2559 DFFNEGX1_33/a_17_74# AND2X2_11/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2560 DFFNEGX1_33/a_31_74# BUFX2_15/Y DFFNEGX1_33/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2561 DFFNEGX1_33/a_17_6# AND2X2_11/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2562 DFFNEGX1_22/a_76_6# BUFX2_16/Y DFFNEGX1_22/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2563 gnd BUFX2_16/Y DFFNEGX1_22/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2564 DFFNEGX1_22/a_66_6# DFFNEGX1_22/a_2_6# DFFNEGX1_22/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2565 out_mines[16] DFFNEGX1_22/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2566 DFFNEGX1_22/a_23_6# BUFX2_16/Y DFFNEGX1_22/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2567 DFFNEGX1_22/a_23_6# DFFNEGX1_22/a_2_6# DFFNEGX1_22/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2568 gnd DFFNEGX1_22/a_34_4# DFFNEGX1_22/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2569 vdd DFFNEGX1_22/a_34_4# DFFNEGX1_22/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2570 DFFNEGX1_22/a_61_74# DFFNEGX1_22/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2571 DFFNEGX1_22/a_34_4# DFFNEGX1_22/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2572 DFFNEGX1_22/a_34_4# DFFNEGX1_22/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2573 vdd out_mines[16] DFFNEGX1_22/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2574 gnd out_mines[16] DFFNEGX1_22/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2575 DFFNEGX1_22/a_61_6# DFFNEGX1_22/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2576 DFFNEGX1_22/a_76_84# DFFNEGX1_22/a_2_6# DFFNEGX1_22/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2577 out_mines[16] DFFNEGX1_22/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2578 vdd BUFX2_16/Y DFFNEGX1_22/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2579 DFFNEGX1_22/a_31_6# DFFNEGX1_22/a_2_6# DFFNEGX1_22/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2580 DFFNEGX1_22/a_66_6# BUFX2_16/Y DFFNEGX1_22/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2581 DFFNEGX1_22/a_17_74# OAI21X1_19/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2582 DFFNEGX1_22/a_31_74# BUFX2_16/Y DFFNEGX1_22/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2583 DFFNEGX1_22/a_17_6# OAI21X1_19/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2584 DFFNEGX1_11/a_76_6# BUFX2_17/Y DFFNEGX1_11/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2585 gnd BUFX2_17/Y DFFNEGX1_11/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2586 DFFNEGX1_11/a_66_6# DFFNEGX1_11/a_2_6# DFFNEGX1_11/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2587 out_mines[15] DFFNEGX1_11/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2588 DFFNEGX1_11/a_23_6# BUFX2_17/Y DFFNEGX1_11/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2589 DFFNEGX1_11/a_23_6# DFFNEGX1_11/a_2_6# DFFNEGX1_11/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2590 gnd DFFNEGX1_11/a_34_4# DFFNEGX1_11/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2591 vdd DFFNEGX1_11/a_34_4# DFFNEGX1_11/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2592 DFFNEGX1_11/a_61_74# DFFNEGX1_11/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2593 DFFNEGX1_11/a_34_4# DFFNEGX1_11/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2594 DFFNEGX1_11/a_34_4# DFFNEGX1_11/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2595 vdd out_mines[15] DFFNEGX1_11/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2596 gnd out_mines[15] DFFNEGX1_11/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2597 DFFNEGX1_11/a_61_6# DFFNEGX1_11/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2598 DFFNEGX1_11/a_76_84# DFFNEGX1_11/a_2_6# DFFNEGX1_11/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2599 out_mines[15] DFFNEGX1_11/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2600 vdd BUFX2_17/Y DFFNEGX1_11/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2601 DFFNEGX1_11/a_31_6# DFFNEGX1_11/a_2_6# DFFNEGX1_11/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2602 DFFNEGX1_11/a_66_6# BUFX2_17/Y DFFNEGX1_11/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2603 DFFNEGX1_11/a_17_74# OAI21X1_21/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2604 DFFNEGX1_11/a_31_74# BUFX2_17/Y DFFNEGX1_11/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2605 DFFNEGX1_11/a_17_6# OAI21X1_21/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2606 DFFNEGX1_44/a_76_6# BUFX2_14/Y DFFNEGX1_44/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2607 gnd BUFX2_14/Y DFFNEGX1_44/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2608 DFFNEGX1_44/a_66_6# DFFNEGX1_44/a_2_6# DFFNEGX1_44/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2609 out_temp_decoded[22] DFFNEGX1_44/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2610 DFFNEGX1_44/a_23_6# BUFX2_14/Y DFFNEGX1_44/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2611 DFFNEGX1_44/a_23_6# DFFNEGX1_44/a_2_6# DFFNEGX1_44/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2612 gnd DFFNEGX1_44/a_34_4# DFFNEGX1_44/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2613 vdd DFFNEGX1_44/a_34_4# DFFNEGX1_44/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2614 DFFNEGX1_44/a_61_74# DFFNEGX1_44/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2615 DFFNEGX1_44/a_34_4# DFFNEGX1_44/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2616 DFFNEGX1_44/a_34_4# DFFNEGX1_44/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2617 vdd out_temp_decoded[22] DFFNEGX1_44/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2618 gnd out_temp_decoded[22] DFFNEGX1_44/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2619 DFFNEGX1_44/a_61_6# DFFNEGX1_44/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2620 DFFNEGX1_44/a_76_84# DFFNEGX1_44/a_2_6# DFFNEGX1_44/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2621 out_temp_decoded[22] DFFNEGX1_44/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2622 vdd BUFX2_14/Y DFFNEGX1_44/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2623 DFFNEGX1_44/a_31_6# DFFNEGX1_44/a_2_6# DFFNEGX1_44/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2624 DFFNEGX1_44/a_66_6# BUFX2_14/Y DFFNEGX1_44/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2625 DFFNEGX1_44/a_17_74# OAI21X1_104/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2626 DFFNEGX1_44/a_31_74# BUFX2_14/Y DFFNEGX1_44/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2627 DFFNEGX1_44/a_17_6# OAI21X1_104/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2628 DFFNEGX1_55/a_76_6# BUFX2_13/Y DFFNEGX1_55/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2629 gnd BUFX2_13/Y DFFNEGX1_55/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2630 DFFNEGX1_55/a_66_6# DFFNEGX1_55/a_2_6# DFFNEGX1_55/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2631 out_temp_decoded[11] DFFNEGX1_55/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2632 DFFNEGX1_55/a_23_6# BUFX2_13/Y DFFNEGX1_55/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2633 DFFNEGX1_55/a_23_6# DFFNEGX1_55/a_2_6# DFFNEGX1_55/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2634 gnd DFFNEGX1_55/a_34_4# DFFNEGX1_55/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2635 vdd DFFNEGX1_55/a_34_4# DFFNEGX1_55/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2636 DFFNEGX1_55/a_61_74# DFFNEGX1_55/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2637 DFFNEGX1_55/a_34_4# DFFNEGX1_55/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2638 DFFNEGX1_55/a_34_4# DFFNEGX1_55/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2639 vdd out_temp_decoded[11] DFFNEGX1_55/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2640 gnd out_temp_decoded[11] DFFNEGX1_55/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2641 DFFNEGX1_55/a_61_6# DFFNEGX1_55/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2642 DFFNEGX1_55/a_76_84# DFFNEGX1_55/a_2_6# DFFNEGX1_55/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2643 out_temp_decoded[11] DFFNEGX1_55/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2644 vdd BUFX2_13/Y DFFNEGX1_55/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2645 DFFNEGX1_55/a_31_6# DFFNEGX1_55/a_2_6# DFFNEGX1_55/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2646 DFFNEGX1_55/a_66_6# BUFX2_13/Y DFFNEGX1_55/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2647 DFFNEGX1_55/a_17_74# OAI21X1_93/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2648 DFFNEGX1_55/a_31_74# BUFX2_13/Y DFFNEGX1_55/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2649 DFFNEGX1_55/a_17_6# OAI21X1_93/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2650 DFFNEGX1_77/a_76_6# BUFX2_12/Y DFFNEGX1_77/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2651 gnd BUFX2_12/Y DFFNEGX1_77/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2652 DFFNEGX1_77/a_66_6# DFFNEGX1_77/a_2_6# DFFNEGX1_77/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2653 out_temp_cleared[14] DFFNEGX1_77/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2654 DFFNEGX1_77/a_23_6# BUFX2_12/Y DFFNEGX1_77/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2655 DFFNEGX1_77/a_23_6# DFFNEGX1_77/a_2_6# DFFNEGX1_77/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2656 gnd DFFNEGX1_77/a_34_4# DFFNEGX1_77/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2657 vdd DFFNEGX1_77/a_34_4# DFFNEGX1_77/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2658 DFFNEGX1_77/a_61_74# DFFNEGX1_77/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2659 DFFNEGX1_77/a_34_4# DFFNEGX1_77/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2660 DFFNEGX1_77/a_34_4# DFFNEGX1_77/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2661 vdd out_temp_cleared[14] DFFNEGX1_77/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2662 gnd out_temp_cleared[14] DFFNEGX1_77/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2663 DFFNEGX1_77/a_61_6# DFFNEGX1_77/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2664 DFFNEGX1_77/a_76_84# DFFNEGX1_77/a_2_6# DFFNEGX1_77/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2665 out_temp_cleared[14] DFFNEGX1_77/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2666 vdd BUFX2_12/Y DFFNEGX1_77/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2667 DFFNEGX1_77/a_31_6# DFFNEGX1_77/a_2_6# DFFNEGX1_77/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2668 DFFNEGX1_77/a_66_6# BUFX2_12/Y DFFNEGX1_77/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2669 DFFNEGX1_77/a_17_74# OAI22X1_14/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2670 DFFNEGX1_77/a_31_74# BUFX2_12/Y DFFNEGX1_77/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2671 DFFNEGX1_77/a_17_6# OAI22X1_14/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2672 DFFNEGX1_66/a_76_6# BUFX2_13/Y DFFNEGX1_66/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2673 gnd BUFX2_13/Y DFFNEGX1_66/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2674 DFFNEGX1_66/a_66_6# DFFNEGX1_66/a_2_6# DFFNEGX1_66/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2675 out_temp_decoded[0] DFFNEGX1_66/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2676 DFFNEGX1_66/a_23_6# BUFX2_13/Y DFFNEGX1_66/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2677 DFFNEGX1_66/a_23_6# DFFNEGX1_66/a_2_6# DFFNEGX1_66/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2678 gnd DFFNEGX1_66/a_34_4# DFFNEGX1_66/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2679 vdd DFFNEGX1_66/a_34_4# DFFNEGX1_66/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2680 DFFNEGX1_66/a_61_74# DFFNEGX1_66/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2681 DFFNEGX1_66/a_34_4# DFFNEGX1_66/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2682 DFFNEGX1_66/a_34_4# DFFNEGX1_66/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2683 vdd out_temp_decoded[0] DFFNEGX1_66/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2684 gnd out_temp_decoded[0] DFFNEGX1_66/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2685 DFFNEGX1_66/a_61_6# DFFNEGX1_66/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2686 DFFNEGX1_66/a_76_84# DFFNEGX1_66/a_2_6# DFFNEGX1_66/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2687 out_temp_decoded[0] DFFNEGX1_66/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2688 vdd BUFX2_13/Y DFFNEGX1_66/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2689 DFFNEGX1_66/a_31_6# DFFNEGX1_66/a_2_6# DFFNEGX1_66/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2690 DFFNEGX1_66/a_66_6# BUFX2_13/Y DFFNEGX1_66/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2691 DFFNEGX1_66/a_17_74# OAI21X1_82/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2692 DFFNEGX1_66/a_31_74# BUFX2_13/Y DFFNEGX1_66/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2693 DFFNEGX1_66/a_17_6# OAI21X1_82/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2694 DFFNEGX1_99/a_76_6# BUFX2_10/Y DFFNEGX1_99/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2695 gnd BUFX2_10/Y DFFNEGX1_99/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2696 DFFNEGX1_99/a_66_6# DFFNEGX1_99/a_2_6# DFFNEGX1_99/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2697 out_global_score[5] DFFNEGX1_99/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2698 DFFNEGX1_99/a_23_6# BUFX2_10/Y DFFNEGX1_99/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2699 DFFNEGX1_99/a_23_6# DFFNEGX1_99/a_2_6# DFFNEGX1_99/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2700 gnd DFFNEGX1_99/a_34_4# DFFNEGX1_99/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2701 vdd DFFNEGX1_99/a_34_4# DFFNEGX1_99/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2702 DFFNEGX1_99/a_61_74# DFFNEGX1_99/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2703 DFFNEGX1_99/a_34_4# DFFNEGX1_99/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2704 DFFNEGX1_99/a_34_4# DFFNEGX1_99/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2705 vdd out_global_score[5] DFFNEGX1_99/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2706 gnd out_global_score[5] DFFNEGX1_99/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2707 DFFNEGX1_99/a_61_6# DFFNEGX1_99/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2708 DFFNEGX1_99/a_76_84# DFFNEGX1_99/a_2_6# DFFNEGX1_99/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2709 out_global_score[5] DFFNEGX1_99/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2710 vdd BUFX2_10/Y DFFNEGX1_99/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2711 DFFNEGX1_99/a_31_6# DFFNEGX1_99/a_2_6# DFFNEGX1_99/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2712 DFFNEGX1_99/a_66_6# BUFX2_10/Y DFFNEGX1_99/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2713 DFFNEGX1_99/a_17_74# INVX2_211/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2714 DFFNEGX1_99/a_31_74# BUFX2_10/Y DFFNEGX1_99/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2715 DFFNEGX1_99/a_17_6# INVX2_211/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2716 DFFNEGX1_88/a_76_6# BUFX2_11/Y DFFNEGX1_88/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2717 gnd BUFX2_11/Y DFFNEGX1_88/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2718 DFFNEGX1_88/a_66_6# DFFNEGX1_88/a_2_6# DFFNEGX1_88/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2719 out_temp_cleared[3] DFFNEGX1_88/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2720 DFFNEGX1_88/a_23_6# BUFX2_11/Y DFFNEGX1_88/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2721 DFFNEGX1_88/a_23_6# DFFNEGX1_88/a_2_6# DFFNEGX1_88/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2722 gnd DFFNEGX1_88/a_34_4# DFFNEGX1_88/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2723 vdd DFFNEGX1_88/a_34_4# DFFNEGX1_88/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2724 DFFNEGX1_88/a_61_74# DFFNEGX1_88/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2725 DFFNEGX1_88/a_34_4# DFFNEGX1_88/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2726 DFFNEGX1_88/a_34_4# DFFNEGX1_88/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2727 vdd out_temp_cleared[3] DFFNEGX1_88/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2728 gnd out_temp_cleared[3] DFFNEGX1_88/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2729 DFFNEGX1_88/a_61_6# DFFNEGX1_88/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2730 DFFNEGX1_88/a_76_84# DFFNEGX1_88/a_2_6# DFFNEGX1_88/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2731 out_temp_cleared[3] DFFNEGX1_88/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2732 vdd BUFX2_11/Y DFFNEGX1_88/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2733 DFFNEGX1_88/a_31_6# DFFNEGX1_88/a_2_6# DFFNEGX1_88/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2734 DFFNEGX1_88/a_66_6# BUFX2_11/Y DFFNEGX1_88/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2735 DFFNEGX1_88/a_17_74# OAI22X1_25/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2736 DFFNEGX1_88/a_31_74# BUFX2_11/Y DFFNEGX1_88/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2737 DFFNEGX1_88/a_17_6# OAI22X1_25/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2738 AND2X2_9/a_2_6# XOR2X1_1/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M2739 AND2X2_9/a_9_6# XOR2X1_1/Y AND2X2_9/a_2_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=100p ps=50u
M2740 AND2X2_9/Y AND2X2_9/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2741 AND2X2_9/Y AND2X2_9/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2742 vdd BUFX2_8/Y AND2X2_9/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2743 gnd BUFX2_8/Y AND2X2_9/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2744 gnd INVX2_49/Y XOR2X1_20/a_2_6# Gnd nfet w=20 l=2
+  ad=70p pd=27u as=100p ps=50u
M2745 XOR2X1_20/Y XOR2X1_20/a_2_6# XOR2X1_20/a_18_6# Gnd nfet w=20 l=2
+  ad=100p pd=30u as=29.999998p ps=23u
M2746 XOR2X1_20/a_13_43# INVX2_44/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=70p ps=27u
M2747 XOR2X1_20/a_18_54# XOR2X1_20/a_13_43# vdd vdd pfet w=40 l=2
+  ad=59.999996p pd=43u as=0.14n ps=47u
M2748 XOR2X1_20/a_35_6# INVX2_49/Y XOR2X1_20/Y Gnd nfet w=20 l=2
+  ad=29.999998p pd=23u as=100p ps=30u
M2749 XOR2X1_20/a_18_6# XOR2X1_20/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=29.999998p pd=23u as=70p ps=27u
M2750 vdd INVX2_49/Y XOR2X1_20/a_2_6# vdd pfet w=40 l=2
+  ad=0.14n pd=47u as=0.2n ps=90u
M2751 vdd INVX2_44/Y XOR2X1_20/a_35_54# vdd pfet w=40 l=2
+  ad=0.14n pd=47u as=59.999996p ps=43u
M2752 XOR2X1_20/Y INVX2_49/Y XOR2X1_20/a_18_54# vdd pfet w=40 l=2
+  ad=0.2n pd=50u as=59.999996p ps=43u
M2753 XOR2X1_20/a_35_54# XOR2X1_20/a_2_6# XOR2X1_20/Y vdd pfet w=40 l=2
+  ad=59.999996p pd=43u as=0.2n ps=50u
M2754 XOR2X1_20/a_13_43# INVX2_44/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.14n ps=47u
M2755 gnd INVX2_44/Y XOR2X1_20/a_35_6# Gnd nfet w=20 l=2
+  ad=70p pd=27u as=29.999998p ps=23u
M2756 DFFNEGX1_101/a_76_6# BUFX2_10/Y DFFNEGX1_101/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2757 gnd BUFX2_10/Y DFFNEGX1_101/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2758 DFFNEGX1_101/a_66_6# DFFNEGX1_101/a_2_6# DFFNEGX1_101/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2759 out_global_score[7] DFFNEGX1_101/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2760 DFFNEGX1_101/a_23_6# BUFX2_10/Y DFFNEGX1_101/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2761 DFFNEGX1_101/a_23_6# DFFNEGX1_101/a_2_6# DFFNEGX1_101/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2762 gnd DFFNEGX1_101/a_34_4# DFFNEGX1_101/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2763 vdd DFFNEGX1_101/a_34_4# DFFNEGX1_101/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2764 DFFNEGX1_101/a_61_74# DFFNEGX1_101/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2765 DFFNEGX1_101/a_34_4# DFFNEGX1_101/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2766 DFFNEGX1_101/a_34_4# DFFNEGX1_101/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2767 vdd out_global_score[7] DFFNEGX1_101/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2768 gnd out_global_score[7] DFFNEGX1_101/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2769 DFFNEGX1_101/a_61_6# DFFNEGX1_101/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2770 DFFNEGX1_101/a_76_84# DFFNEGX1_101/a_2_6# DFFNEGX1_101/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2771 out_global_score[7] DFFNEGX1_101/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2772 vdd BUFX2_10/Y DFFNEGX1_101/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2773 DFFNEGX1_101/a_31_6# DFFNEGX1_101/a_2_6# DFFNEGX1_101/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2774 DFFNEGX1_101/a_66_6# BUFX2_10/Y DFFNEGX1_101/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2775 DFFNEGX1_101/a_17_74# INVX2_209/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2776 DFFNEGX1_101/a_31_74# BUFX2_10/Y DFFNEGX1_101/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2777 DFFNEGX1_101/a_17_6# INVX2_209/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2778 DFFNEGX1_112/a_76_6# BUFX2_9/Y DFFNEGX1_112/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2779 gnd BUFX2_9/Y DFFNEGX1_112/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2780 DFFNEGX1_112/a_66_6# DFFNEGX1_112/a_2_6# DFFNEGX1_112/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2781 out_global_score[18] DFFNEGX1_112/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2782 DFFNEGX1_112/a_23_6# BUFX2_9/Y DFFNEGX1_112/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2783 DFFNEGX1_112/a_23_6# DFFNEGX1_112/a_2_6# DFFNEGX1_112/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2784 gnd DFFNEGX1_112/a_34_4# DFFNEGX1_112/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2785 vdd DFFNEGX1_112/a_34_4# DFFNEGX1_112/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2786 DFFNEGX1_112/a_61_74# DFFNEGX1_112/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2787 DFFNEGX1_112/a_34_4# DFFNEGX1_112/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2788 DFFNEGX1_112/a_34_4# DFFNEGX1_112/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2789 vdd out_global_score[18] DFFNEGX1_112/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2790 gnd out_global_score[18] DFFNEGX1_112/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2791 DFFNEGX1_112/a_61_6# DFFNEGX1_112/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2792 DFFNEGX1_112/a_76_84# DFFNEGX1_112/a_2_6# DFFNEGX1_112/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2793 out_global_score[18] DFFNEGX1_112/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2794 vdd BUFX2_9/Y DFFNEGX1_112/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2795 DFFNEGX1_112/a_31_6# DFFNEGX1_112/a_2_6# DFFNEGX1_112/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2796 DFFNEGX1_112/a_66_6# BUFX2_9/Y DFFNEGX1_112/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2797 DFFNEGX1_112/a_17_74# INVX2_198/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2798 DFFNEGX1_112/a_31_74# BUFX2_9/Y DFFNEGX1_112/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2799 DFFNEGX1_112/a_17_6# INVX2_198/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2800 DFFNEGX1_134/a_76_6# INVX2_259/Y DFFNEGX1_134/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2801 gnd INVX2_259/Y DFFNEGX1_134/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2802 DFFNEGX1_134/a_66_6# DFFNEGX1_134/a_2_6# DFFNEGX1_134/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2803 out_state_main[2] DFFNEGX1_134/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2804 DFFNEGX1_134/a_23_6# INVX2_259/Y DFFNEGX1_134/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2805 DFFNEGX1_134/a_23_6# DFFNEGX1_134/a_2_6# DFFNEGX1_134/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2806 gnd DFFNEGX1_134/a_34_4# DFFNEGX1_134/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2807 vdd DFFNEGX1_134/a_34_4# DFFNEGX1_134/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2808 DFFNEGX1_134/a_61_74# DFFNEGX1_134/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2809 DFFNEGX1_134/a_34_4# DFFNEGX1_134/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2810 DFFNEGX1_134/a_34_4# DFFNEGX1_134/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2811 vdd out_state_main[2] DFFNEGX1_134/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2812 gnd out_state_main[2] DFFNEGX1_134/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2813 DFFNEGX1_134/a_61_6# DFFNEGX1_134/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2814 DFFNEGX1_134/a_76_84# DFFNEGX1_134/a_2_6# DFFNEGX1_134/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2815 out_state_main[2] DFFNEGX1_134/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2816 vdd INVX2_259/Y DFFNEGX1_134/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2817 DFFNEGX1_134/a_31_6# DFFNEGX1_134/a_2_6# DFFNEGX1_134/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2818 DFFNEGX1_134/a_66_6# INVX2_259/Y DFFNEGX1_134/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2819 DFFNEGX1_134/a_17_74# INVX2_119/A vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2820 DFFNEGX1_134/a_31_74# INVX2_259/Y DFFNEGX1_134/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2821 DFFNEGX1_134/a_17_6# INVX2_119/A gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2822 DFFNEGX1_123/a_76_6# BUFX2_5/Y DFFNEGX1_123/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2823 gnd BUFX2_5/Y DFFNEGX1_123/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2824 DFFNEGX1_123/a_66_6# DFFNEGX1_123/a_2_6# DFFNEGX1_123/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2825 out_global_score[29] DFFNEGX1_123/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2826 DFFNEGX1_123/a_23_6# BUFX2_5/Y DFFNEGX1_123/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2827 DFFNEGX1_123/a_23_6# DFFNEGX1_123/a_2_6# DFFNEGX1_123/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2828 gnd DFFNEGX1_123/a_34_4# DFFNEGX1_123/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2829 vdd DFFNEGX1_123/a_34_4# DFFNEGX1_123/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2830 DFFNEGX1_123/a_61_74# DFFNEGX1_123/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2831 DFFNEGX1_123/a_34_4# DFFNEGX1_123/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2832 DFFNEGX1_123/a_34_4# DFFNEGX1_123/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2833 vdd out_global_score[29] DFFNEGX1_123/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2834 gnd out_global_score[29] DFFNEGX1_123/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2835 DFFNEGX1_123/a_61_6# DFFNEGX1_123/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2836 DFFNEGX1_123/a_76_84# DFFNEGX1_123/a_2_6# DFFNEGX1_123/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2837 out_global_score[29] DFFNEGX1_123/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2838 vdd BUFX2_5/Y DFFNEGX1_123/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2839 DFFNEGX1_123/a_31_6# DFFNEGX1_123/a_2_6# DFFNEGX1_123/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2840 DFFNEGX1_123/a_66_6# BUFX2_5/Y DFFNEGX1_123/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2841 DFFNEGX1_123/a_17_74# INVX2_187/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2842 DFFNEGX1_123/a_31_74# BUFX2_5/Y DFFNEGX1_123/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2843 DFFNEGX1_123/a_17_6# INVX2_187/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2844 gnd out_global_score[29] AOI22X1_4/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M2845 INVX2_187/A INVX2_258/Y AOI22X1_4/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2846 AOI22X1_4/a_11_6# HAX1_1/YS gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2847 AOI22X1_4/a_2_54# INVX2_258/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M2848 AOI22X1_4/a_28_6# INVX2_255/Y INVX2_187/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2849 vdd HAX1_1/YS AOI22X1_4/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2850 INVX2_187/A INVX2_255/Y AOI22X1_4/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M2851 AOI22X1_4/a_2_54# out_global_score[29] INVX2_187/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2852 gnd OAI22X1_80/Y OAI21X1_150/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M2853 vdd XOR2X1_4/Y AOI21X1_17/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M2854 AOI21X1_17/A XOR2X1_4/Y OAI21X1_150/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2855 AOI21X1_17/A OAI22X1_79/Y OAI21X1_150/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2856 OAI21X1_150/a_9_54# OAI22X1_80/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2857 OAI21X1_150/a_2_6# OAI22X1_79/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2858 gnd out_state_main[3] OAI21X1_161/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M2859 vdd AND2X2_19/B AOI21X1_23/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M2860 AOI21X1_23/C AND2X2_19/B OAI21X1_161/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2861 AOI21X1_23/C AOI22X1_78/Y OAI21X1_161/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M2862 OAI21X1_161/a_9_54# out_state_main[3] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2863 OAI21X1_161/a_2_6# AOI22X1_78/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2864 OAI21X1_19/C out_mines[16] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M2865 NAND2X1_25/a_9_6# out_mines[16] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2866 vdd INVX2_224/Y OAI21X1_19/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2867 OAI21X1_19/C INVX2_224/Y NAND2X1_25/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2868 NAND2X1_14/Y NAND3X1_6/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M2869 NAND2X1_14/a_9_6# NAND3X1_6/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2870 vdd OR2X1_13/Y NAND2X1_14/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2871 NAND2X1_14/Y OR2X1_13/Y NAND2X1_14/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2872 OAI21X1_51/C out_mines[0] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M2873 NAND2X1_47/a_9_6# out_mines[0] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2874 vdd INVX2_226/Y OAI21X1_51/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2875 OAI21X1_51/C INVX2_226/Y NAND2X1_47/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2876 OAI21X1_37/C out_mines[7] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M2877 NAND2X1_36/a_9_6# out_mines[7] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2878 vdd INVX2_231/Y OAI21X1_37/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2879 OAI21X1_37/C INVX2_231/Y NAND2X1_36/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2880 OAI21X1_60/A OAI21X1_61/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M2881 NAND2X1_58/a_9_6# OAI21X1_61/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2882 vdd AOI21X1_3/A OAI21X1_60/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2883 OAI21X1_60/A AOI21X1_3/A NAND2X1_58/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2884 OAI21X1_82/C NOR2X1_59/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M2885 NAND2X1_69/a_9_6# NOR2X1_59/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2886 vdd BUFX2_21/A OAI21X1_82/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2887 OAI21X1_82/C BUFX2_21/A NAND2X1_69/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2888 gnd out_global_score[10] AOI22X1_23/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M2889 INVX2_206/A INVX2_258/Y AOI22X1_23/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2890 AOI22X1_23/a_11_6# HAX1_20/YS gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2891 AOI22X1_23/a_2_54# INVX2_258/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M2892 AOI22X1_23/a_28_6# OR2X1_11/B INVX2_206/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2893 vdd HAX1_20/YS AOI22X1_23/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2894 INVX2_206/A OR2X1_11/B AOI22X1_23/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M2895 AOI22X1_23/a_2_54# out_global_score[10] INVX2_206/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2896 gnd out_global_score[21] AOI22X1_12/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M2897 INVX2_195/A INVX2_257/Y AOI22X1_12/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2898 AOI22X1_12/a_11_6# HAX1_9/YS gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2899 AOI22X1_12/a_2_54# INVX2_257/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M2900 AOI22X1_12/a_28_6# INVX2_255/Y INVX2_195/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2901 vdd HAX1_9/YS AOI22X1_12/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2902 INVX2_195/A INVX2_255/Y AOI22X1_12/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M2903 AOI22X1_12/a_2_54# out_global_score[21] INVX2_195/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2904 gnd out_temp_cleared[14] AOI22X1_45/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M2905 NAND3X1_39/A out_mines[13] AOI22X1_45/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2906 AOI22X1_45/a_11_6# out_temp_cleared[13] gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2907 AOI22X1_45/a_2_54# out_mines[13] vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M2908 AOI22X1_45/a_28_6# out_mines[14] NAND3X1_39/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2909 vdd out_temp_cleared[13] AOI22X1_45/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2910 NAND3X1_39/A out_mines[14] AOI22X1_45/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M2911 AOI22X1_45/a_2_54# out_temp_cleared[14] NAND3X1_39/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2912 gnd out_temp_decoded[22] AOI22X1_34/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M2913 NAND2X1_63/B out_mines[21] AOI22X1_34/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2914 AOI22X1_34/a_11_6# out_temp_decoded[21] gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2915 AOI22X1_34/a_2_54# out_mines[21] vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M2916 AOI22X1_34/a_28_6# out_mines[22] NAND2X1_63/B Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2917 vdd out_temp_decoded[21] AOI22X1_34/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2918 NAND2X1_63/B out_mines[22] AOI22X1_34/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M2919 AOI22X1_34/a_2_54# out_temp_decoded[22] NAND2X1_63/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2920 gnd INVX2_31/Y AOI22X1_56/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M2921 OAI22X1_36/C AOI21X1_9/A AOI22X1_56/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2922 AOI22X1_56/a_11_6# INVX2_32/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2923 AOI22X1_56/a_2_54# AOI21X1_9/A vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M2924 AOI22X1_56/a_28_6# INVX2_47/A OAI22X1_36/C Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2925 vdd INVX2_32/Y AOI22X1_56/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2926 OAI22X1_36/C INVX2_47/A AOI22X1_56/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M2927 AOI22X1_56/a_2_54# INVX2_31/Y OAI22X1_36/C vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2928 gnd out_state_main[0] AOI22X1_78/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M2929 AOI22X1_78/Y INVX2_116/Y AOI22X1_78/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2930 AOI22X1_78/a_11_6# NOR2X1_121/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2931 AOI22X1_78/a_2_54# INVX2_116/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M2932 AOI22X1_78/a_28_6# INVX2_125/Y AOI22X1_78/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2933 vdd NOR2X1_121/Y AOI22X1_78/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2934 AOI22X1_78/Y INVX2_125/Y AOI22X1_78/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M2935 AOI22X1_78/a_2_54# out_state_main[0] AOI22X1_78/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2936 gnd INVX2_31/Y AOI22X1_67/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M2937 AOI22X1_67/Y out_mines[6] AOI22X1_67/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M2938 AOI22X1_67/a_11_6# INVX2_32/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2939 AOI22X1_67/a_2_54# out_mines[6] vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M2940 AOI22X1_67/a_28_6# out_mines[14] AOI22X1_67/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2941 vdd INVX2_32/Y AOI22X1_67/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2942 AOI22X1_67/Y out_mines[14] AOI22X1_67/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M2943 AOI22X1_67/a_2_54# INVX2_31/Y AOI22X1_67/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2944 gnd BUFX2_25/Y OAI22X1_7/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M2945 OAI22X1_7/a_2_6# OR2X1_11/A OAI22X1_7/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M2946 OAI22X1_7/Y INVX2_59/Y OAI22X1_7/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2947 OAI22X1_7/Y INVX2_92/Y OAI22X1_7/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M2948 OAI22X1_7/a_28_54# INVX2_59/Y OAI22X1_7/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2949 OAI22X1_7/a_9_54# BUFX2_25/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2950 OAI22X1_7/a_2_6# INVX2_92/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2951 vdd OR2X1_11/A OAI22X1_7/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2952 INVX2_27/Y out_mines[10] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2953 INVX2_27/Y out_mines[10] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2954 INVX2_16/Y out_mines[9] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2955 INVX2_16/Y out_mines[9] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2956 INVX2_38/Y XOR2X1_3/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2957 INVX2_38/Y XOR2X1_3/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2958 INVX2_49/Y INVX2_49/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2959 INVX2_49/Y INVX2_49/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2960 gnd MUX2X1_0/A MUX2X1_0/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M2961 MUX2X1_0/a_17_50# MUX2X1_0/B vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2962 MUX2X1_0/Y NOR2X1_7/Y MUX2X1_0/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M2963 MUX2X1_0/a_30_54# MUX2X1_0/a_2_10# MUX2X1_0/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M2964 MUX2X1_0/a_17_10# MUX2X1_0/B gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2965 vdd NOR2X1_7/Y MUX2X1_0/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2966 MUX2X1_0/a_30_10# NOR2X1_7/Y MUX2X1_0/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M2967 gnd NOR2X1_7/Y MUX2X1_0/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M2968 vdd MUX2X1_0/A MUX2X1_0/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M2969 MUX2X1_0/Y MUX2X1_0/a_2_10# MUX2X1_0/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2970 MUX2X1_7/B MUX2X1_3/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2971 MUX2X1_7/B MUX2X1_3/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2972 OR2X1_0/A MUX2X1_25/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2973 OR2X1_0/A MUX2X1_25/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2974 HAX1_42/A MUX2X1_12/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2975 HAX1_42/A MUX2X1_12/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2976 NOR2X1_65/A NOR2X1_63/B gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2977 NOR2X1_65/A NOR2X1_63/B vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2978 INVX2_194/Y INVX2_194/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2979 INVX2_194/Y INVX2_194/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2980 DFFNEGX1_23/a_76_6# BUFX2_16/Y DFFNEGX1_23/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M2981 gnd BUFX2_16/Y DFFNEGX1_23/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M2982 DFFNEGX1_23/a_66_6# DFFNEGX1_23/a_2_6# DFFNEGX1_23/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2983 out_mines[17] DFFNEGX1_23/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2984 DFFNEGX1_23/a_23_6# BUFX2_16/Y DFFNEGX1_23/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M2985 DFFNEGX1_23/a_23_6# DFFNEGX1_23/a_2_6# DFFNEGX1_23/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M2986 gnd DFFNEGX1_23/a_34_4# DFFNEGX1_23/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2987 vdd DFFNEGX1_23/a_34_4# DFFNEGX1_23/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M2988 DFFNEGX1_23/a_61_74# DFFNEGX1_23/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M2989 DFFNEGX1_23/a_34_4# DFFNEGX1_23/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M2990 DFFNEGX1_23/a_34_4# DFFNEGX1_23/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M2991 vdd out_mines[17] DFFNEGX1_23/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M2992 gnd out_mines[17] DFFNEGX1_23/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2993 DFFNEGX1_23/a_61_6# DFFNEGX1_23/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2994 DFFNEGX1_23/a_76_84# DFFNEGX1_23/a_2_6# DFFNEGX1_23/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M2995 out_mines[17] DFFNEGX1_23/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M2996 vdd BUFX2_16/Y DFFNEGX1_23/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M2997 DFFNEGX1_23/a_31_6# DFFNEGX1_23/a_2_6# DFFNEGX1_23/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M2998 DFFNEGX1_23/a_66_6# BUFX2_16/Y DFFNEGX1_23/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M2999 DFFNEGX1_23/a_17_74# OAI21X1_17/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3000 DFFNEGX1_23/a_31_74# BUFX2_16/Y DFFNEGX1_23/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3001 DFFNEGX1_23/a_17_6# OAI21X1_17/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3002 DFFNEGX1_12/a_76_6# BUFX2_17/Y DFFNEGX1_12/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3003 gnd BUFX2_17/Y DFFNEGX1_12/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3004 DFFNEGX1_12/a_66_6# DFFNEGX1_12/a_2_6# DFFNEGX1_12/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3005 out_mines[13] DFFNEGX1_12/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3006 DFFNEGX1_12/a_23_6# BUFX2_17/Y DFFNEGX1_12/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3007 DFFNEGX1_12/a_23_6# DFFNEGX1_12/a_2_6# DFFNEGX1_12/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3008 gnd DFFNEGX1_12/a_34_4# DFFNEGX1_12/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3009 vdd DFFNEGX1_12/a_34_4# DFFNEGX1_12/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3010 DFFNEGX1_12/a_61_74# DFFNEGX1_12/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3011 DFFNEGX1_12/a_34_4# DFFNEGX1_12/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3012 DFFNEGX1_12/a_34_4# DFFNEGX1_12/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3013 vdd out_mines[13] DFFNEGX1_12/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3014 gnd out_mines[13] DFFNEGX1_12/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3015 DFFNEGX1_12/a_61_6# DFFNEGX1_12/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3016 DFFNEGX1_12/a_76_84# DFFNEGX1_12/a_2_6# DFFNEGX1_12/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3017 out_mines[13] DFFNEGX1_12/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3018 vdd BUFX2_17/Y DFFNEGX1_12/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3019 DFFNEGX1_12/a_31_6# DFFNEGX1_12/a_2_6# DFFNEGX1_12/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3020 DFFNEGX1_12/a_66_6# BUFX2_17/Y DFFNEGX1_12/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3021 DFFNEGX1_12/a_17_74# OAI21X1_25/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3022 DFFNEGX1_12/a_31_74# BUFX2_17/Y DFFNEGX1_12/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3023 DFFNEGX1_12/a_17_6# OAI21X1_25/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3024 DFFNEGX1_34/a_76_6# BUFX2_15/Y DFFNEGX1_34/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3025 gnd BUFX2_15/Y DFFNEGX1_34/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3026 DFFNEGX1_34/a_66_6# DFFNEGX1_34/a_2_6# DFFNEGX1_34/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3027 out_temp_mine_cnt[3] DFFNEGX1_34/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3028 DFFNEGX1_34/a_23_6# BUFX2_15/Y DFFNEGX1_34/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3029 DFFNEGX1_34/a_23_6# DFFNEGX1_34/a_2_6# DFFNEGX1_34/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3030 gnd DFFNEGX1_34/a_34_4# DFFNEGX1_34/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3031 vdd DFFNEGX1_34/a_34_4# DFFNEGX1_34/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3032 DFFNEGX1_34/a_61_74# DFFNEGX1_34/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3033 DFFNEGX1_34/a_34_4# DFFNEGX1_34/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3034 DFFNEGX1_34/a_34_4# DFFNEGX1_34/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3035 vdd out_temp_mine_cnt[3] DFFNEGX1_34/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3036 gnd out_temp_mine_cnt[3] DFFNEGX1_34/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3037 DFFNEGX1_34/a_61_6# DFFNEGX1_34/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3038 DFFNEGX1_34/a_76_84# DFFNEGX1_34/a_2_6# DFFNEGX1_34/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3039 out_temp_mine_cnt[3] DFFNEGX1_34/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3040 vdd BUFX2_15/Y DFFNEGX1_34/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3041 DFFNEGX1_34/a_31_6# DFFNEGX1_34/a_2_6# DFFNEGX1_34/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3042 DFFNEGX1_34/a_66_6# BUFX2_15/Y DFFNEGX1_34/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3043 DFFNEGX1_34/a_17_74# AND2X2_10/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3044 DFFNEGX1_34/a_31_74# BUFX2_15/Y DFFNEGX1_34/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3045 DFFNEGX1_34/a_17_6# AND2X2_10/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3046 DFFNEGX1_56/a_76_6# BUFX2_13/Y DFFNEGX1_56/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3047 gnd BUFX2_13/Y DFFNEGX1_56/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3048 DFFNEGX1_56/a_66_6# DFFNEGX1_56/a_2_6# DFFNEGX1_56/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3049 out_temp_decoded[10] DFFNEGX1_56/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3050 DFFNEGX1_56/a_23_6# BUFX2_13/Y DFFNEGX1_56/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3051 DFFNEGX1_56/a_23_6# DFFNEGX1_56/a_2_6# DFFNEGX1_56/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3052 gnd DFFNEGX1_56/a_34_4# DFFNEGX1_56/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3053 vdd DFFNEGX1_56/a_34_4# DFFNEGX1_56/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3054 DFFNEGX1_56/a_61_74# DFFNEGX1_56/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3055 DFFNEGX1_56/a_34_4# DFFNEGX1_56/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3056 DFFNEGX1_56/a_34_4# DFFNEGX1_56/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3057 vdd out_temp_decoded[10] DFFNEGX1_56/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3058 gnd out_temp_decoded[10] DFFNEGX1_56/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3059 DFFNEGX1_56/a_61_6# DFFNEGX1_56/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3060 DFFNEGX1_56/a_76_84# DFFNEGX1_56/a_2_6# DFFNEGX1_56/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3061 out_temp_decoded[10] DFFNEGX1_56/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3062 vdd BUFX2_13/Y DFFNEGX1_56/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3063 DFFNEGX1_56/a_31_6# DFFNEGX1_56/a_2_6# DFFNEGX1_56/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3064 DFFNEGX1_56/a_66_6# BUFX2_13/Y DFFNEGX1_56/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3065 DFFNEGX1_56/a_17_74# OAI21X1_92/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3066 DFFNEGX1_56/a_31_74# BUFX2_13/Y DFFNEGX1_56/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3067 DFFNEGX1_56/a_17_6# OAI21X1_92/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3068 DFFNEGX1_45/a_76_6# BUFX2_14/Y DFFNEGX1_45/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3069 gnd BUFX2_14/Y DFFNEGX1_45/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3070 DFFNEGX1_45/a_66_6# DFFNEGX1_45/a_2_6# DFFNEGX1_45/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3071 out_temp_decoded[21] DFFNEGX1_45/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3072 DFFNEGX1_45/a_23_6# BUFX2_14/Y DFFNEGX1_45/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3073 DFFNEGX1_45/a_23_6# DFFNEGX1_45/a_2_6# DFFNEGX1_45/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3074 gnd DFFNEGX1_45/a_34_4# DFFNEGX1_45/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3075 vdd DFFNEGX1_45/a_34_4# DFFNEGX1_45/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3076 DFFNEGX1_45/a_61_74# DFFNEGX1_45/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3077 DFFNEGX1_45/a_34_4# DFFNEGX1_45/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3078 DFFNEGX1_45/a_34_4# DFFNEGX1_45/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3079 vdd out_temp_decoded[21] DFFNEGX1_45/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3080 gnd out_temp_decoded[21] DFFNEGX1_45/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3081 DFFNEGX1_45/a_61_6# DFFNEGX1_45/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3082 DFFNEGX1_45/a_76_84# DFFNEGX1_45/a_2_6# DFFNEGX1_45/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3083 out_temp_decoded[21] DFFNEGX1_45/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3084 vdd BUFX2_14/Y DFFNEGX1_45/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3085 DFFNEGX1_45/a_31_6# DFFNEGX1_45/a_2_6# DFFNEGX1_45/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3086 DFFNEGX1_45/a_66_6# BUFX2_14/Y DFFNEGX1_45/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3087 DFFNEGX1_45/a_17_74# OAI21X1_103/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3088 DFFNEGX1_45/a_31_74# BUFX2_14/Y DFFNEGX1_45/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3089 DFFNEGX1_45/a_17_6# OAI21X1_103/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3090 DFFNEGX1_67/a_76_6# BUFX2_12/Y DFFNEGX1_67/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3091 gnd BUFX2_12/Y DFFNEGX1_67/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3092 DFFNEGX1_67/a_66_6# DFFNEGX1_67/a_2_6# DFFNEGX1_67/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3093 out_temp_cleared[24] DFFNEGX1_67/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3094 DFFNEGX1_67/a_23_6# BUFX2_12/Y DFFNEGX1_67/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3095 DFFNEGX1_67/a_23_6# DFFNEGX1_67/a_2_6# DFFNEGX1_67/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3096 gnd DFFNEGX1_67/a_34_4# DFFNEGX1_67/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3097 vdd DFFNEGX1_67/a_34_4# DFFNEGX1_67/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3098 DFFNEGX1_67/a_61_74# DFFNEGX1_67/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3099 DFFNEGX1_67/a_34_4# DFFNEGX1_67/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3100 DFFNEGX1_67/a_34_4# DFFNEGX1_67/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3101 vdd out_temp_cleared[24] DFFNEGX1_67/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3102 gnd out_temp_cleared[24] DFFNEGX1_67/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3103 DFFNEGX1_67/a_61_6# DFFNEGX1_67/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3104 DFFNEGX1_67/a_76_84# DFFNEGX1_67/a_2_6# DFFNEGX1_67/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3105 out_temp_cleared[24] DFFNEGX1_67/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3106 vdd BUFX2_12/Y DFFNEGX1_67/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3107 DFFNEGX1_67/a_31_6# DFFNEGX1_67/a_2_6# DFFNEGX1_67/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3108 DFFNEGX1_67/a_66_6# BUFX2_12/Y DFFNEGX1_67/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3109 DFFNEGX1_67/a_17_74# OAI22X1_4/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3110 DFFNEGX1_67/a_31_74# BUFX2_12/Y DFFNEGX1_67/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3111 DFFNEGX1_67/a_17_6# OAI22X1_4/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3112 DFFNEGX1_78/a_76_6# BUFX2_12/Y DFFNEGX1_78/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3113 gnd BUFX2_12/Y DFFNEGX1_78/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3114 DFFNEGX1_78/a_66_6# DFFNEGX1_78/a_2_6# DFFNEGX1_78/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3115 out_temp_cleared[13] DFFNEGX1_78/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3116 DFFNEGX1_78/a_23_6# BUFX2_12/Y DFFNEGX1_78/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3117 DFFNEGX1_78/a_23_6# DFFNEGX1_78/a_2_6# DFFNEGX1_78/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3118 gnd DFFNEGX1_78/a_34_4# DFFNEGX1_78/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3119 vdd DFFNEGX1_78/a_34_4# DFFNEGX1_78/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3120 DFFNEGX1_78/a_61_74# DFFNEGX1_78/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3121 DFFNEGX1_78/a_34_4# DFFNEGX1_78/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3122 DFFNEGX1_78/a_34_4# DFFNEGX1_78/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3123 vdd out_temp_cleared[13] DFFNEGX1_78/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3124 gnd out_temp_cleared[13] DFFNEGX1_78/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3125 DFFNEGX1_78/a_61_6# DFFNEGX1_78/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3126 DFFNEGX1_78/a_76_84# DFFNEGX1_78/a_2_6# DFFNEGX1_78/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3127 out_temp_cleared[13] DFFNEGX1_78/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3128 vdd BUFX2_12/Y DFFNEGX1_78/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3129 DFFNEGX1_78/a_31_6# DFFNEGX1_78/a_2_6# DFFNEGX1_78/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3130 DFFNEGX1_78/a_66_6# BUFX2_12/Y DFFNEGX1_78/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3131 DFFNEGX1_78/a_17_74# OAI22X1_15/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3132 DFFNEGX1_78/a_31_74# BUFX2_12/Y DFFNEGX1_78/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3133 DFFNEGX1_78/a_17_6# OAI22X1_15/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3134 DFFNEGX1_89/a_76_6# BUFX2_11/Y DFFNEGX1_89/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3135 gnd BUFX2_11/Y DFFNEGX1_89/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3136 DFFNEGX1_89/a_66_6# DFFNEGX1_89/a_2_6# DFFNEGX1_89/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3137 out_temp_cleared[2] DFFNEGX1_89/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3138 DFFNEGX1_89/a_23_6# BUFX2_11/Y DFFNEGX1_89/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3139 DFFNEGX1_89/a_23_6# DFFNEGX1_89/a_2_6# DFFNEGX1_89/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3140 gnd DFFNEGX1_89/a_34_4# DFFNEGX1_89/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3141 vdd DFFNEGX1_89/a_34_4# DFFNEGX1_89/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3142 DFFNEGX1_89/a_61_74# DFFNEGX1_89/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3143 DFFNEGX1_89/a_34_4# DFFNEGX1_89/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3144 DFFNEGX1_89/a_34_4# DFFNEGX1_89/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3145 vdd out_temp_cleared[2] DFFNEGX1_89/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3146 gnd out_temp_cleared[2] DFFNEGX1_89/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3147 DFFNEGX1_89/a_61_6# DFFNEGX1_89/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3148 DFFNEGX1_89/a_76_84# DFFNEGX1_89/a_2_6# DFFNEGX1_89/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3149 out_temp_cleared[2] DFFNEGX1_89/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3150 vdd BUFX2_11/Y DFFNEGX1_89/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3151 DFFNEGX1_89/a_31_6# DFFNEGX1_89/a_2_6# DFFNEGX1_89/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3152 DFFNEGX1_89/a_66_6# BUFX2_11/Y DFFNEGX1_89/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3153 DFFNEGX1_89/a_17_74# OAI22X1_26/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3154 DFFNEGX1_89/a_31_74# BUFX2_11/Y DFFNEGX1_89/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3155 DFFNEGX1_89/a_17_6# OAI22X1_26/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3156 gnd in_incr[0] XOR2X1_10/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3157 NOR2X1_0/B XOR2X1_10/a_2_6# XOR2X1_10/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3158 XOR2X1_10/a_13_43# NOR2X1_8/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3159 XOR2X1_10/a_18_54# XOR2X1_10/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3160 XOR2X1_10/a_35_6# in_incr[0] NOR2X1_0/B Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3161 XOR2X1_10/a_18_6# XOR2X1_10/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3162 vdd in_incr[0] XOR2X1_10/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3163 vdd NOR2X1_8/Y XOR2X1_10/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3164 NOR2X1_0/B in_incr[0] XOR2X1_10/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3165 XOR2X1_10/a_35_54# XOR2X1_10/a_2_6# NOR2X1_0/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3166 XOR2X1_10/a_13_43# NOR2X1_8/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3167 gnd NOR2X1_8/Y XOR2X1_10/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3168 gnd XOR2X1_22/Y XOR2X1_21/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3169 INVX2_49/A XOR2X1_21/a_2_6# XOR2X1_21/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3170 XOR2X1_21/a_13_43# INVX2_40/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3171 XOR2X1_21/a_18_54# XOR2X1_21/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3172 XOR2X1_21/a_35_6# XOR2X1_22/Y INVX2_49/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3173 XOR2X1_21/a_18_6# XOR2X1_21/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3174 vdd XOR2X1_22/Y XOR2X1_21/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3175 vdd INVX2_40/Y XOR2X1_21/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3176 INVX2_49/A XOR2X1_22/Y XOR2X1_21/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3177 XOR2X1_21/a_35_54# XOR2X1_21/a_2_6# INVX2_49/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3178 XOR2X1_21/a_13_43# INVX2_40/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3179 gnd INVX2_40/Y XOR2X1_21/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3180 DFFNEGX1_102/a_76_6# BUFX2_10/Y DFFNEGX1_102/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3181 gnd BUFX2_10/Y DFFNEGX1_102/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3182 DFFNEGX1_102/a_66_6# DFFNEGX1_102/a_2_6# DFFNEGX1_102/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3183 out_global_score[8] DFFNEGX1_102/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3184 DFFNEGX1_102/a_23_6# BUFX2_10/Y DFFNEGX1_102/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3185 DFFNEGX1_102/a_23_6# DFFNEGX1_102/a_2_6# DFFNEGX1_102/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3186 gnd DFFNEGX1_102/a_34_4# DFFNEGX1_102/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3187 vdd DFFNEGX1_102/a_34_4# DFFNEGX1_102/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3188 DFFNEGX1_102/a_61_74# DFFNEGX1_102/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3189 DFFNEGX1_102/a_34_4# DFFNEGX1_102/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3190 DFFNEGX1_102/a_34_4# DFFNEGX1_102/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3191 vdd out_global_score[8] DFFNEGX1_102/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3192 gnd out_global_score[8] DFFNEGX1_102/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3193 DFFNEGX1_102/a_61_6# DFFNEGX1_102/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3194 DFFNEGX1_102/a_76_84# DFFNEGX1_102/a_2_6# DFFNEGX1_102/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3195 out_global_score[8] DFFNEGX1_102/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3196 vdd BUFX2_10/Y DFFNEGX1_102/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3197 DFFNEGX1_102/a_31_6# DFFNEGX1_102/a_2_6# DFFNEGX1_102/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3198 DFFNEGX1_102/a_66_6# BUFX2_10/Y DFFNEGX1_102/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3199 DFFNEGX1_102/a_17_74# INVX2_208/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3200 DFFNEGX1_102/a_31_74# BUFX2_10/Y DFFNEGX1_102/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3201 DFFNEGX1_102/a_17_6# INVX2_208/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3202 NOR2X1_40/B OAI21X1_1/A vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=26u as=100p ps=50u
M3203 NAND3X1_0/a_9_6# OAI21X1_1/A gnd Gnd nfet w=30 l=2
+  ad=45p pd=33u as=0.15n ps=70u
M3204 NOR2X1_40/B out_temp_data_in[2] vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=59.999996p ps=26u
M3205 NOR2X1_40/B out_temp_data_in[2] NAND3X1_0/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=45p ps=33u
M3206 vdd INVX2_30/Y NOR2X1_40/B vdd pfet w=20 l=2
+  ad=59.999996p pd=26u as=59.999996p ps=26u
M3207 NAND3X1_0/a_14_6# INVX2_30/Y NAND3X1_0/a_9_6# Gnd nfet w=30 l=2
+  ad=45p pd=33u as=45p ps=33u
M3208 DFFNEGX1_113/a_76_6# BUFX2_9/Y DFFNEGX1_113/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3209 gnd BUFX2_9/Y DFFNEGX1_113/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3210 DFFNEGX1_113/a_66_6# DFFNEGX1_113/a_2_6# DFFNEGX1_113/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3211 out_global_score[19] DFFNEGX1_113/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3212 DFFNEGX1_113/a_23_6# BUFX2_9/Y DFFNEGX1_113/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3213 DFFNEGX1_113/a_23_6# DFFNEGX1_113/a_2_6# DFFNEGX1_113/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3214 gnd DFFNEGX1_113/a_34_4# DFFNEGX1_113/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3215 vdd DFFNEGX1_113/a_34_4# DFFNEGX1_113/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3216 DFFNEGX1_113/a_61_74# DFFNEGX1_113/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3217 DFFNEGX1_113/a_34_4# DFFNEGX1_113/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3218 DFFNEGX1_113/a_34_4# DFFNEGX1_113/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3219 vdd out_global_score[19] DFFNEGX1_113/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3220 gnd out_global_score[19] DFFNEGX1_113/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3221 DFFNEGX1_113/a_61_6# DFFNEGX1_113/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3222 DFFNEGX1_113/a_76_84# DFFNEGX1_113/a_2_6# DFFNEGX1_113/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3223 out_global_score[19] DFFNEGX1_113/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3224 vdd BUFX2_9/Y DFFNEGX1_113/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3225 DFFNEGX1_113/a_31_6# DFFNEGX1_113/a_2_6# DFFNEGX1_113/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3226 DFFNEGX1_113/a_66_6# BUFX2_9/Y DFFNEGX1_113/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3227 DFFNEGX1_113/a_17_74# INVX2_197/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3228 DFFNEGX1_113/a_31_74# BUFX2_9/Y DFFNEGX1_113/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3229 DFFNEGX1_113/a_17_6# INVX2_197/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3230 DFFNEGX1_135/a_76_6# BUFX2_5/Y DFFNEGX1_135/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3231 gnd BUFX2_5/Y DFFNEGX1_135/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3232 DFFNEGX1_135/a_66_6# DFFNEGX1_135/a_2_6# DFFNEGX1_135/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3233 INVX2_120/A DFFNEGX1_135/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3234 DFFNEGX1_135/a_23_6# BUFX2_5/Y DFFNEGX1_135/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3235 DFFNEGX1_135/a_23_6# DFFNEGX1_135/a_2_6# DFFNEGX1_135/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3236 gnd DFFNEGX1_135/a_34_4# DFFNEGX1_135/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3237 vdd DFFNEGX1_135/a_34_4# DFFNEGX1_135/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3238 DFFNEGX1_135/a_61_74# DFFNEGX1_135/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3239 DFFNEGX1_135/a_34_4# DFFNEGX1_135/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3240 DFFNEGX1_135/a_34_4# DFFNEGX1_135/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3241 vdd INVX2_120/A DFFNEGX1_135/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3242 gnd INVX2_120/A DFFNEGX1_135/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3243 DFFNEGX1_135/a_61_6# DFFNEGX1_135/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3244 DFFNEGX1_135/a_76_84# DFFNEGX1_135/a_2_6# DFFNEGX1_135/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3245 INVX2_120/A DFFNEGX1_135/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3246 vdd BUFX2_5/Y DFFNEGX1_135/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3247 DFFNEGX1_135/a_31_6# DFFNEGX1_135/a_2_6# DFFNEGX1_135/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3248 DFFNEGX1_135/a_66_6# BUFX2_5/Y DFFNEGX1_135/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3249 DFFNEGX1_135/a_17_74# NOR2X1_119/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3250 DFFNEGX1_135/a_31_74# BUFX2_5/Y DFFNEGX1_135/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3251 DFFNEGX1_135/a_17_6# NOR2X1_119/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3252 DFFNEGX1_124/a_76_6# BUFX2_5/Y DFFNEGX1_124/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3253 gnd BUFX2_5/Y DFFNEGX1_124/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3254 DFFNEGX1_124/a_66_6# DFFNEGX1_124/a_2_6# DFFNEGX1_124/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3255 out_global_score[30] DFFNEGX1_124/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3256 DFFNEGX1_124/a_23_6# BUFX2_5/Y DFFNEGX1_124/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3257 DFFNEGX1_124/a_23_6# DFFNEGX1_124/a_2_6# DFFNEGX1_124/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3258 gnd DFFNEGX1_124/a_34_4# DFFNEGX1_124/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3259 vdd DFFNEGX1_124/a_34_4# DFFNEGX1_124/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3260 DFFNEGX1_124/a_61_74# DFFNEGX1_124/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3261 DFFNEGX1_124/a_34_4# DFFNEGX1_124/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3262 DFFNEGX1_124/a_34_4# DFFNEGX1_124/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3263 vdd out_global_score[30] DFFNEGX1_124/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3264 gnd out_global_score[30] DFFNEGX1_124/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3265 DFFNEGX1_124/a_61_6# DFFNEGX1_124/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3266 DFFNEGX1_124/a_76_84# DFFNEGX1_124/a_2_6# DFFNEGX1_124/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3267 out_global_score[30] DFFNEGX1_124/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3268 vdd BUFX2_5/Y DFFNEGX1_124/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3269 DFFNEGX1_124/a_31_6# DFFNEGX1_124/a_2_6# DFFNEGX1_124/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3270 DFFNEGX1_124/a_66_6# BUFX2_5/Y DFFNEGX1_124/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3271 DFFNEGX1_124/a_17_74# INVX2_186/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3272 DFFNEGX1_124/a_31_74# BUFX2_5/Y DFFNEGX1_124/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3273 DFFNEGX1_124/a_17_6# INVX2_186/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3274 gnd out_global_score[28] AOI22X1_5/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M3275 INVX2_188/A INVX2_257/Y AOI22X1_5/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3276 AOI22X1_5/a_11_6# HAX1_2/YS gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3277 AOI22X1_5/a_2_54# INVX2_257/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M3278 AOI22X1_5/a_28_6# INVX2_255/Y INVX2_188/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3279 vdd HAX1_2/YS AOI22X1_5/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3280 INVX2_188/A INVX2_255/Y AOI22X1_5/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M3281 AOI22X1_5/a_2_54# out_global_score[28] INVX2_188/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3282 gnd AOI21X1_16/Y OAI21X1_140/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M3283 vdd XOR2X1_11/Y OAI21X1_140/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M3284 OAI21X1_140/Y XOR2X1_11/Y OAI21X1_140/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3285 OAI21X1_140/Y AOI21X1_15/Y OAI21X1_140/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3286 OAI21X1_140/a_9_54# AOI21X1_16/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3287 OAI21X1_140/a_2_6# AOI21X1_15/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3288 gnd OAI22X1_82/Y OAI21X1_151/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M3289 vdd INVX2_35/Y AOI21X1_18/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M3290 AOI21X1_18/B INVX2_35/Y OAI21X1_151/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3291 AOI21X1_18/B OAI22X1_81/Y OAI21X1_151/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3292 OAI21X1_151/a_9_54# OAI22X1_82/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3293 OAI21X1_151/a_2_6# OAI22X1_81/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3294 gnd in_place OAI21X1_162/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M3295 vdd INVX2_125/Y AOI21X1_26/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M3296 AOI21X1_26/A INVX2_125/Y OAI21X1_162/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3297 AOI21X1_26/A out_state_main[2] OAI21X1_162/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3298 OAI21X1_162/a_9_54# in_place vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3299 OAI21X1_162/a_2_6# out_state_main[2] gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3300 OAI21X1_3/C out_mines[24] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M3301 NAND2X1_15/a_9_6# out_mines[24] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3302 vdd OAI21X1_3/A OAI21X1_3/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3303 OAI21X1_3/C OAI21X1_3/A NAND2X1_15/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3304 OAI21X1_53/C out_temp_index[4] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M3305 NAND2X1_48/a_9_6# out_temp_index[4] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3306 vdd NOR2X1_67/Y OAI21X1_53/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3307 OAI21X1_53/C NOR2X1_67/Y NAND2X1_48/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3308 OAI21X1_39/C out_mines[6] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M3309 NAND2X1_37/a_9_6# out_mines[6] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3310 vdd INVX2_232/Y OAI21X1_39/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3311 OAI21X1_39/C INVX2_232/Y NAND2X1_37/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3312 OAI21X1_21/C out_mines[15] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M3313 NAND2X1_26/a_9_6# out_mines[15] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3314 vdd INVX2_229/Y OAI21X1_21/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3315 OAI21X1_21/C INVX2_229/Y NAND2X1_26/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3316 OAI21X1_62/C out_n_nearby[1] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M3317 NAND2X1_59/a_9_6# out_n_nearby[1] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3318 vdd AOI21X1_2/A OAI21X1_62/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3319 OAI21X1_62/C AOI21X1_2/A NAND2X1_59/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3320 gnd out_global_score[9] AOI22X1_24/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M3321 INVX2_207/A INVX2_258/Y AOI22X1_24/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3322 AOI22X1_24/a_11_6# HAX1_21/YS gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3323 AOI22X1_24/a_2_54# INVX2_258/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M3324 AOI22X1_24/a_28_6# OR2X1_11/B INVX2_207/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3325 vdd HAX1_21/YS AOI22X1_24/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3326 INVX2_207/A OR2X1_11/B AOI22X1_24/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M3327 AOI22X1_24/a_2_54# out_global_score[9] INVX2_207/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3328 gnd out_global_score[20] AOI22X1_13/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M3329 INVX2_196/A INVX2_257/Y AOI22X1_13/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3330 AOI22X1_13/a_11_6# HAX1_10/YS gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3331 AOI22X1_13/a_2_54# INVX2_257/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M3332 AOI22X1_13/a_28_6# INVX2_255/Y INVX2_196/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3333 vdd HAX1_10/YS AOI22X1_13/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3334 INVX2_196/A INVX2_255/Y AOI22X1_13/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M3335 AOI22X1_13/a_2_54# out_global_score[20] INVX2_196/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3336 gnd out_temp_cleared[17] AOI22X1_46/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M3337 NAND3X1_41/B out_mines[16] AOI22X1_46/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3338 AOI22X1_46/a_11_6# out_temp_cleared[16] gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3339 AOI22X1_46/a_2_54# out_mines[16] vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M3340 AOI22X1_46/a_28_6# out_mines[17] NAND3X1_41/B Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3341 vdd out_temp_cleared[16] AOI22X1_46/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3342 NAND3X1_41/B out_mines[17] AOI22X1_46/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M3343 AOI22X1_46/a_2_54# out_temp_cleared[17] NAND3X1_41/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3344 gnd out_temp_decoded[24] AOI22X1_35/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M3345 NAND2X1_63/A out_mines[23] AOI22X1_35/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3346 AOI22X1_35/a_11_6# out_temp_decoded[23] gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3347 AOI22X1_35/a_2_54# out_mines[23] vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M3348 AOI22X1_35/a_28_6# out_mines[24] NAND2X1_63/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3349 vdd out_temp_decoded[23] AOI22X1_35/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3350 NAND2X1_63/A out_mines[24] AOI22X1_35/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M3351 AOI22X1_35/a_2_54# out_temp_decoded[24] NAND2X1_63/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3352 gnd out_temp_data_in[2] AOI22X1_57/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M3353 OAI22X1_37/D OAI21X1_1/B AOI22X1_57/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3354 AOI22X1_57/a_11_6# AOI22X1_57/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3355 AOI22X1_57/a_2_54# OAI21X1_1/B vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M3356 AOI22X1_57/a_28_6# INVX2_42/Y OAI22X1_37/D Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3357 vdd AOI22X1_57/A AOI22X1_57/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3358 OAI22X1_37/D INVX2_42/Y AOI22X1_57/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M3359 AOI22X1_57/a_2_54# out_temp_data_in[2] OAI22X1_37/D vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3360 gnd INVX2_31/Y AOI22X1_68/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M3361 AOI22X1_68/Y out_mines[5] AOI22X1_68/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3362 AOI22X1_68/a_11_6# INVX2_32/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3363 AOI22X1_68/a_2_54# out_mines[5] vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M3364 AOI22X1_68/a_28_6# out_mines[13] AOI22X1_68/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3365 vdd INVX2_32/Y AOI22X1_68/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3366 AOI22X1_68/Y out_mines[13] AOI22X1_68/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M3367 AOI22X1_68/a_2_54# INVX2_31/Y AOI22X1_68/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3368 gnd BUFX2_25/Y OAI22X1_8/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M3369 OAI22X1_8/a_2_6# OR2X1_11/A OAI22X1_8/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M3370 OAI22X1_8/Y INVX2_60/Y OAI22X1_8/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3371 OAI22X1_8/Y INVX2_93/Y OAI22X1_8/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M3372 OAI22X1_8/a_28_54# INVX2_60/Y OAI22X1_8/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3373 OAI22X1_8/a_9_54# BUFX2_25/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3374 OAI22X1_8/a_2_6# INVX2_93/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3375 vdd OR2X1_11/A OAI22X1_8/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3376 INVX2_17/Y out_temp_index[4] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3377 INVX2_17/Y out_temp_index[4] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3378 INVX2_39/Y INVX2_39/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3379 INVX2_39/Y INVX2_39/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3380 INVX2_28/Y out_mines[3] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3381 INVX2_28/Y out_mines[3] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3382 gnd XOR2X1_0/A XOR2X1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3383 XOR2X1_0/Y XOR2X1_0/a_2_6# XOR2X1_0/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3384 XOR2X1_0/a_13_43# XOR2X1_5/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3385 XOR2X1_0/a_18_54# XOR2X1_0/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3386 XOR2X1_0/a_35_6# XOR2X1_0/A XOR2X1_0/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3387 XOR2X1_0/a_18_6# XOR2X1_0/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3388 vdd XOR2X1_0/A XOR2X1_0/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3389 vdd XOR2X1_5/Y XOR2X1_0/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3390 XOR2X1_0/Y XOR2X1_0/A XOR2X1_0/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3391 XOR2X1_0/a_35_54# XOR2X1_0/a_2_6# XOR2X1_0/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3392 XOR2X1_0/a_13_43# XOR2X1_5/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3393 gnd XOR2X1_5/Y XOR2X1_0/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3394 gnd XOR2X1_0/Y MUX2X1_1/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M3395 MUX2X1_1/a_17_50# XOR2X1_5/Y vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3396 MUX2X1_1/Y NOR2X1_7/Y MUX2X1_1/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M3397 MUX2X1_1/a_30_54# MUX2X1_1/a_2_10# MUX2X1_1/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3398 MUX2X1_1/a_17_10# XOR2X1_5/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3399 vdd NOR2X1_7/Y MUX2X1_1/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3400 MUX2X1_1/a_30_10# NOR2X1_7/Y MUX2X1_1/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M3401 gnd NOR2X1_7/Y MUX2X1_1/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M3402 vdd XOR2X1_0/Y MUX2X1_1/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3403 MUX2X1_1/Y MUX2X1_1/a_2_10# MUX2X1_1/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3404 NOR2X1_27/B in_mult[3] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3405 NOR2X1_27/B in_mult[3] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3406 OR2X1_2/A MUX2X1_15/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3407 OR2X1_2/A MUX2X1_15/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3408 HAX1_49/A MUX2X1_26/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3409 HAX1_49/A MUX2X1_26/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3410 NOR2X1_5/A MUX2X1_4/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3411 NOR2X1_5/A MUX2X1_4/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3412 INVX2_184/Y INVX2_184/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3413 INVX2_184/Y INVX2_184/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3414 INVX2_195/Y INVX2_195/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3415 INVX2_195/Y INVX2_195/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3416 DFFNEGX1_13/a_76_6# BUFX2_17/Y DFFNEGX1_13/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3417 gnd BUFX2_17/Y DFFNEGX1_13/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3418 DFFNEGX1_13/a_66_6# DFFNEGX1_13/a_2_6# DFFNEGX1_13/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3419 out_mines[14] DFFNEGX1_13/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3420 DFFNEGX1_13/a_23_6# BUFX2_17/Y DFFNEGX1_13/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3421 DFFNEGX1_13/a_23_6# DFFNEGX1_13/a_2_6# DFFNEGX1_13/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3422 gnd DFFNEGX1_13/a_34_4# DFFNEGX1_13/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3423 vdd DFFNEGX1_13/a_34_4# DFFNEGX1_13/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3424 DFFNEGX1_13/a_61_74# DFFNEGX1_13/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3425 DFFNEGX1_13/a_34_4# DFFNEGX1_13/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3426 DFFNEGX1_13/a_34_4# DFFNEGX1_13/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3427 vdd out_mines[14] DFFNEGX1_13/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3428 gnd out_mines[14] DFFNEGX1_13/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3429 DFFNEGX1_13/a_61_6# DFFNEGX1_13/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3430 DFFNEGX1_13/a_76_84# DFFNEGX1_13/a_2_6# DFFNEGX1_13/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3431 out_mines[14] DFFNEGX1_13/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3432 vdd BUFX2_17/Y DFFNEGX1_13/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3433 DFFNEGX1_13/a_31_6# DFFNEGX1_13/a_2_6# DFFNEGX1_13/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3434 DFFNEGX1_13/a_66_6# BUFX2_17/Y DFFNEGX1_13/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3435 DFFNEGX1_13/a_17_74# OAI21X1_23/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3436 DFFNEGX1_13/a_31_74# BUFX2_17/Y DFFNEGX1_13/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3437 DFFNEGX1_13/a_17_6# OAI21X1_23/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3438 DFFNEGX1_24/a_76_6# BUFX2_16/Y DFFNEGX1_24/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3439 gnd BUFX2_16/Y DFFNEGX1_24/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3440 DFFNEGX1_24/a_66_6# DFFNEGX1_24/a_2_6# DFFNEGX1_24/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3441 out_mines[24] DFFNEGX1_24/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3442 DFFNEGX1_24/a_23_6# BUFX2_16/Y DFFNEGX1_24/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3443 DFFNEGX1_24/a_23_6# DFFNEGX1_24/a_2_6# DFFNEGX1_24/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3444 gnd DFFNEGX1_24/a_34_4# DFFNEGX1_24/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3445 vdd DFFNEGX1_24/a_34_4# DFFNEGX1_24/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3446 DFFNEGX1_24/a_61_74# DFFNEGX1_24/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3447 DFFNEGX1_24/a_34_4# DFFNEGX1_24/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3448 DFFNEGX1_24/a_34_4# DFFNEGX1_24/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3449 vdd out_mines[24] DFFNEGX1_24/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3450 gnd out_mines[24] DFFNEGX1_24/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3451 DFFNEGX1_24/a_61_6# DFFNEGX1_24/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3452 DFFNEGX1_24/a_76_84# DFFNEGX1_24/a_2_6# DFFNEGX1_24/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3453 out_mines[24] DFFNEGX1_24/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3454 vdd BUFX2_16/Y DFFNEGX1_24/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3455 DFFNEGX1_24/a_31_6# DFFNEGX1_24/a_2_6# DFFNEGX1_24/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3456 DFFNEGX1_24/a_66_6# BUFX2_16/Y DFFNEGX1_24/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3457 DFFNEGX1_24/a_17_74# OAI21X1_3/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3458 DFFNEGX1_24/a_31_74# BUFX2_16/Y DFFNEGX1_24/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3459 DFFNEGX1_24/a_17_6# OAI21X1_3/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3460 DFFNEGX1_35/a_76_6# BUFX2_15/Y DFFNEGX1_35/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3461 gnd BUFX2_15/Y DFFNEGX1_35/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3462 DFFNEGX1_35/a_66_6# DFFNEGX1_35/a_2_6# DFFNEGX1_35/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3463 out_temp_mine_cnt[4] DFFNEGX1_35/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3464 DFFNEGX1_35/a_23_6# BUFX2_15/Y DFFNEGX1_35/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3465 DFFNEGX1_35/a_23_6# DFFNEGX1_35/a_2_6# DFFNEGX1_35/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3466 gnd DFFNEGX1_35/a_34_4# DFFNEGX1_35/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3467 vdd DFFNEGX1_35/a_34_4# DFFNEGX1_35/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3468 DFFNEGX1_35/a_61_74# DFFNEGX1_35/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3469 DFFNEGX1_35/a_34_4# DFFNEGX1_35/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3470 DFFNEGX1_35/a_34_4# DFFNEGX1_35/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3471 vdd out_temp_mine_cnt[4] DFFNEGX1_35/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3472 gnd out_temp_mine_cnt[4] DFFNEGX1_35/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3473 DFFNEGX1_35/a_61_6# DFFNEGX1_35/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3474 DFFNEGX1_35/a_76_84# DFFNEGX1_35/a_2_6# DFFNEGX1_35/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3475 out_temp_mine_cnt[4] DFFNEGX1_35/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3476 vdd BUFX2_15/Y DFFNEGX1_35/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3477 DFFNEGX1_35/a_31_6# DFFNEGX1_35/a_2_6# DFFNEGX1_35/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3478 DFFNEGX1_35/a_66_6# BUFX2_15/Y DFFNEGX1_35/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3479 DFFNEGX1_35/a_17_74# AND2X2_9/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3480 DFFNEGX1_35/a_31_74# BUFX2_15/Y DFFNEGX1_35/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3481 DFFNEGX1_35/a_17_6# AND2X2_9/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3482 DFFNEGX1_68/a_76_6# BUFX2_12/Y DFFNEGX1_68/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3483 gnd BUFX2_12/Y DFFNEGX1_68/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3484 DFFNEGX1_68/a_66_6# DFFNEGX1_68/a_2_6# DFFNEGX1_68/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3485 out_temp_cleared[23] DFFNEGX1_68/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3486 DFFNEGX1_68/a_23_6# BUFX2_12/Y DFFNEGX1_68/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3487 DFFNEGX1_68/a_23_6# DFFNEGX1_68/a_2_6# DFFNEGX1_68/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3488 gnd DFFNEGX1_68/a_34_4# DFFNEGX1_68/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3489 vdd DFFNEGX1_68/a_34_4# DFFNEGX1_68/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3490 DFFNEGX1_68/a_61_74# DFFNEGX1_68/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3491 DFFNEGX1_68/a_34_4# DFFNEGX1_68/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3492 DFFNEGX1_68/a_34_4# DFFNEGX1_68/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3493 vdd out_temp_cleared[23] DFFNEGX1_68/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3494 gnd out_temp_cleared[23] DFFNEGX1_68/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3495 DFFNEGX1_68/a_61_6# DFFNEGX1_68/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3496 DFFNEGX1_68/a_76_84# DFFNEGX1_68/a_2_6# DFFNEGX1_68/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3497 out_temp_cleared[23] DFFNEGX1_68/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3498 vdd BUFX2_12/Y DFFNEGX1_68/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3499 DFFNEGX1_68/a_31_6# DFFNEGX1_68/a_2_6# DFFNEGX1_68/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3500 DFFNEGX1_68/a_66_6# BUFX2_12/Y DFFNEGX1_68/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3501 DFFNEGX1_68/a_17_74# OAI22X1_5/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3502 DFFNEGX1_68/a_31_74# BUFX2_12/Y DFFNEGX1_68/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3503 DFFNEGX1_68/a_17_6# OAI22X1_5/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3504 DFFNEGX1_57/a_76_6# BUFX2_13/Y DFFNEGX1_57/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3505 gnd BUFX2_13/Y DFFNEGX1_57/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3506 DFFNEGX1_57/a_66_6# DFFNEGX1_57/a_2_6# DFFNEGX1_57/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3507 out_temp_decoded[9] DFFNEGX1_57/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3508 DFFNEGX1_57/a_23_6# BUFX2_13/Y DFFNEGX1_57/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3509 DFFNEGX1_57/a_23_6# DFFNEGX1_57/a_2_6# DFFNEGX1_57/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3510 gnd DFFNEGX1_57/a_34_4# DFFNEGX1_57/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3511 vdd DFFNEGX1_57/a_34_4# DFFNEGX1_57/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3512 DFFNEGX1_57/a_61_74# DFFNEGX1_57/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3513 DFFNEGX1_57/a_34_4# DFFNEGX1_57/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3514 DFFNEGX1_57/a_34_4# DFFNEGX1_57/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3515 vdd out_temp_decoded[9] DFFNEGX1_57/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3516 gnd out_temp_decoded[9] DFFNEGX1_57/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3517 DFFNEGX1_57/a_61_6# DFFNEGX1_57/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3518 DFFNEGX1_57/a_76_84# DFFNEGX1_57/a_2_6# DFFNEGX1_57/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3519 out_temp_decoded[9] DFFNEGX1_57/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3520 vdd BUFX2_13/Y DFFNEGX1_57/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3521 DFFNEGX1_57/a_31_6# DFFNEGX1_57/a_2_6# DFFNEGX1_57/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3522 DFFNEGX1_57/a_66_6# BUFX2_13/Y DFFNEGX1_57/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3523 DFFNEGX1_57/a_17_74# OAI21X1_91/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3524 DFFNEGX1_57/a_31_74# BUFX2_13/Y DFFNEGX1_57/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3525 DFFNEGX1_57/a_17_6# OAI21X1_91/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3526 DFFNEGX1_46/a_76_6# BUFX2_14/Y DFFNEGX1_46/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3527 gnd BUFX2_14/Y DFFNEGX1_46/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3528 DFFNEGX1_46/a_66_6# DFFNEGX1_46/a_2_6# DFFNEGX1_46/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3529 out_temp_decoded[20] DFFNEGX1_46/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3530 DFFNEGX1_46/a_23_6# BUFX2_14/Y DFFNEGX1_46/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3531 DFFNEGX1_46/a_23_6# DFFNEGX1_46/a_2_6# DFFNEGX1_46/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3532 gnd DFFNEGX1_46/a_34_4# DFFNEGX1_46/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3533 vdd DFFNEGX1_46/a_34_4# DFFNEGX1_46/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3534 DFFNEGX1_46/a_61_74# DFFNEGX1_46/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3535 DFFNEGX1_46/a_34_4# DFFNEGX1_46/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3536 DFFNEGX1_46/a_34_4# DFFNEGX1_46/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3537 vdd out_temp_decoded[20] DFFNEGX1_46/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3538 gnd out_temp_decoded[20] DFFNEGX1_46/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3539 DFFNEGX1_46/a_61_6# DFFNEGX1_46/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3540 DFFNEGX1_46/a_76_84# DFFNEGX1_46/a_2_6# DFFNEGX1_46/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3541 out_temp_decoded[20] DFFNEGX1_46/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3542 vdd BUFX2_14/Y DFFNEGX1_46/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3543 DFFNEGX1_46/a_31_6# DFFNEGX1_46/a_2_6# DFFNEGX1_46/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3544 DFFNEGX1_46/a_66_6# BUFX2_14/Y DFFNEGX1_46/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3545 DFFNEGX1_46/a_17_74# OAI21X1_102/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3546 DFFNEGX1_46/a_31_74# BUFX2_14/Y DFFNEGX1_46/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3547 DFFNEGX1_46/a_17_6# OAI21X1_102/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3548 DFFNEGX1_79/a_76_6# BUFX2_12/Y DFFNEGX1_79/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3549 gnd BUFX2_12/Y DFFNEGX1_79/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3550 DFFNEGX1_79/a_66_6# DFFNEGX1_79/a_2_6# DFFNEGX1_79/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3551 out_temp_cleared[12] DFFNEGX1_79/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3552 DFFNEGX1_79/a_23_6# BUFX2_12/Y DFFNEGX1_79/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3553 DFFNEGX1_79/a_23_6# DFFNEGX1_79/a_2_6# DFFNEGX1_79/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3554 gnd DFFNEGX1_79/a_34_4# DFFNEGX1_79/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3555 vdd DFFNEGX1_79/a_34_4# DFFNEGX1_79/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3556 DFFNEGX1_79/a_61_74# DFFNEGX1_79/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3557 DFFNEGX1_79/a_34_4# DFFNEGX1_79/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3558 DFFNEGX1_79/a_34_4# DFFNEGX1_79/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3559 vdd out_temp_cleared[12] DFFNEGX1_79/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3560 gnd out_temp_cleared[12] DFFNEGX1_79/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3561 DFFNEGX1_79/a_61_6# DFFNEGX1_79/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3562 DFFNEGX1_79/a_76_84# DFFNEGX1_79/a_2_6# DFFNEGX1_79/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3563 out_temp_cleared[12] DFFNEGX1_79/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3564 vdd BUFX2_12/Y DFFNEGX1_79/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3565 DFFNEGX1_79/a_31_6# DFFNEGX1_79/a_2_6# DFFNEGX1_79/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3566 DFFNEGX1_79/a_66_6# BUFX2_12/Y DFFNEGX1_79/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3567 DFFNEGX1_79/a_17_74# OAI22X1_16/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3568 DFFNEGX1_79/a_31_74# BUFX2_12/Y DFFNEGX1_79/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3569 DFFNEGX1_79/a_17_6# OAI22X1_16/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3570 gnd out_temp_data_in[4] XOR2X1_11/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3571 XOR2X1_11/Y XOR2X1_11/a_2_6# XOR2X1_11/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3572 XOR2X1_11/a_13_43# OR2X1_8/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3573 XOR2X1_11/a_18_54# XOR2X1_11/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3574 XOR2X1_11/a_35_6# out_temp_data_in[4] XOR2X1_11/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3575 XOR2X1_11/a_18_6# XOR2X1_11/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3576 vdd out_temp_data_in[4] XOR2X1_11/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3577 vdd OR2X1_8/Y XOR2X1_11/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3578 XOR2X1_11/Y out_temp_data_in[4] XOR2X1_11/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3579 XOR2X1_11/a_35_54# XOR2X1_11/a_2_6# XOR2X1_11/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3580 XOR2X1_11/a_13_43# OR2X1_8/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3581 gnd OR2X1_8/Y XOR2X1_11/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3582 gnd XOR2X1_29/B XOR2X1_22/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3583 XOR2X1_22/Y XOR2X1_22/a_2_6# XOR2X1_22/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3584 XOR2X1_22/a_13_43# INVX2_50/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3585 XOR2X1_22/a_18_54# XOR2X1_22/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3586 XOR2X1_22/a_35_6# XOR2X1_29/B XOR2X1_22/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3587 XOR2X1_22/a_18_6# XOR2X1_22/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3588 vdd XOR2X1_29/B XOR2X1_22/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3589 vdd INVX2_50/A XOR2X1_22/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3590 XOR2X1_22/Y XOR2X1_29/B XOR2X1_22/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3591 XOR2X1_22/a_35_54# XOR2X1_22/a_2_6# XOR2X1_22/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3592 XOR2X1_22/a_13_43# INVX2_50/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3593 gnd INVX2_50/A XOR2X1_22/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3594 NOR2X1_47/B out_temp_data_in[2] vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M3595 NAND3X1_1/a_9_6# out_temp_data_in[2] gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M3596 NOR2X1_47/B out_temp_data_in[4] vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3597 NOR2X1_47/B out_temp_data_in[4] NAND3X1_1/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M3598 vdd OAI21X1_1/A NOR2X1_47/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3599 NAND3X1_1/a_14_6# OAI21X1_1/A NAND3X1_1/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M3600 DFFNEGX1_103/a_76_6# BUFX2_10/Y DFFNEGX1_103/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3601 gnd BUFX2_10/Y DFFNEGX1_103/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3602 DFFNEGX1_103/a_66_6# DFFNEGX1_103/a_2_6# DFFNEGX1_103/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3603 out_global_score[9] DFFNEGX1_103/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3604 DFFNEGX1_103/a_23_6# BUFX2_10/Y DFFNEGX1_103/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3605 DFFNEGX1_103/a_23_6# DFFNEGX1_103/a_2_6# DFFNEGX1_103/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3606 gnd DFFNEGX1_103/a_34_4# DFFNEGX1_103/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3607 vdd DFFNEGX1_103/a_34_4# DFFNEGX1_103/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3608 DFFNEGX1_103/a_61_74# DFFNEGX1_103/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3609 DFFNEGX1_103/a_34_4# DFFNEGX1_103/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3610 DFFNEGX1_103/a_34_4# DFFNEGX1_103/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3611 vdd out_global_score[9] DFFNEGX1_103/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3612 gnd out_global_score[9] DFFNEGX1_103/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3613 DFFNEGX1_103/a_61_6# DFFNEGX1_103/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3614 DFFNEGX1_103/a_76_84# DFFNEGX1_103/a_2_6# DFFNEGX1_103/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3615 out_global_score[9] DFFNEGX1_103/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3616 vdd BUFX2_10/Y DFFNEGX1_103/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3617 DFFNEGX1_103/a_31_6# DFFNEGX1_103/a_2_6# DFFNEGX1_103/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3618 DFFNEGX1_103/a_66_6# BUFX2_10/Y DFFNEGX1_103/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3619 DFFNEGX1_103/a_17_74# INVX2_207/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3620 DFFNEGX1_103/a_31_74# BUFX2_10/Y DFFNEGX1_103/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3621 DFFNEGX1_103/a_17_6# INVX2_207/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3622 DFFNEGX1_114/a_76_6# BUFX2_9/Y DFFNEGX1_114/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3623 gnd BUFX2_9/Y DFFNEGX1_114/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3624 DFFNEGX1_114/a_66_6# DFFNEGX1_114/a_2_6# DFFNEGX1_114/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3625 out_global_score[20] DFFNEGX1_114/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3626 DFFNEGX1_114/a_23_6# BUFX2_9/Y DFFNEGX1_114/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3627 DFFNEGX1_114/a_23_6# DFFNEGX1_114/a_2_6# DFFNEGX1_114/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3628 gnd DFFNEGX1_114/a_34_4# DFFNEGX1_114/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3629 vdd DFFNEGX1_114/a_34_4# DFFNEGX1_114/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3630 DFFNEGX1_114/a_61_74# DFFNEGX1_114/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3631 DFFNEGX1_114/a_34_4# DFFNEGX1_114/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3632 DFFNEGX1_114/a_34_4# DFFNEGX1_114/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3633 vdd out_global_score[20] DFFNEGX1_114/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3634 gnd out_global_score[20] DFFNEGX1_114/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3635 DFFNEGX1_114/a_61_6# DFFNEGX1_114/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3636 DFFNEGX1_114/a_76_84# DFFNEGX1_114/a_2_6# DFFNEGX1_114/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3637 out_global_score[20] DFFNEGX1_114/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3638 vdd BUFX2_9/Y DFFNEGX1_114/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3639 DFFNEGX1_114/a_31_6# DFFNEGX1_114/a_2_6# DFFNEGX1_114/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3640 DFFNEGX1_114/a_66_6# BUFX2_9/Y DFFNEGX1_114/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3641 DFFNEGX1_114/a_17_74# INVX2_196/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3642 DFFNEGX1_114/a_31_74# BUFX2_9/Y DFFNEGX1_114/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3643 DFFNEGX1_114/a_17_6# INVX2_196/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3644 DFFNEGX1_125/a_76_6# BUFX2_5/Y DFFNEGX1_125/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3645 gnd BUFX2_5/Y DFFNEGX1_125/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3646 DFFNEGX1_125/a_66_6# DFFNEGX1_125/a_2_6# DFFNEGX1_125/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3647 out_global_score[31] DFFNEGX1_125/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3648 DFFNEGX1_125/a_23_6# BUFX2_5/Y DFFNEGX1_125/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3649 DFFNEGX1_125/a_23_6# DFFNEGX1_125/a_2_6# DFFNEGX1_125/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3650 gnd DFFNEGX1_125/a_34_4# DFFNEGX1_125/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3651 vdd DFFNEGX1_125/a_34_4# DFFNEGX1_125/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3652 DFFNEGX1_125/a_61_74# DFFNEGX1_125/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3653 DFFNEGX1_125/a_34_4# DFFNEGX1_125/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3654 DFFNEGX1_125/a_34_4# DFFNEGX1_125/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3655 vdd out_global_score[31] DFFNEGX1_125/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3656 gnd out_global_score[31] DFFNEGX1_125/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3657 DFFNEGX1_125/a_61_6# DFFNEGX1_125/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3658 DFFNEGX1_125/a_76_84# DFFNEGX1_125/a_2_6# DFFNEGX1_125/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3659 out_global_score[31] DFFNEGX1_125/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3660 vdd BUFX2_5/Y DFFNEGX1_125/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3661 DFFNEGX1_125/a_31_6# DFFNEGX1_125/a_2_6# DFFNEGX1_125/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3662 DFFNEGX1_125/a_66_6# BUFX2_5/Y DFFNEGX1_125/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3663 DFFNEGX1_125/a_17_74# INVX2_185/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3664 DFFNEGX1_125/a_31_74# BUFX2_5/Y DFFNEGX1_125/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3665 DFFNEGX1_125/a_17_6# INVX2_185/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3666 DFFNEGX1_136/a_76_6# INVX2_259/Y DFFNEGX1_136/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3667 gnd INVX2_259/Y DFFNEGX1_136/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3668 DFFNEGX1_136/a_66_6# DFFNEGX1_136/a_2_6# DFFNEGX1_136/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3669 out_state_main[1] DFFNEGX1_136/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3670 DFFNEGX1_136/a_23_6# INVX2_259/Y DFFNEGX1_136/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3671 DFFNEGX1_136/a_23_6# DFFNEGX1_136/a_2_6# DFFNEGX1_136/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3672 gnd DFFNEGX1_136/a_34_4# DFFNEGX1_136/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3673 vdd DFFNEGX1_136/a_34_4# DFFNEGX1_136/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3674 DFFNEGX1_136/a_61_74# DFFNEGX1_136/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3675 DFFNEGX1_136/a_34_4# DFFNEGX1_136/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3676 DFFNEGX1_136/a_34_4# DFFNEGX1_136/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3677 vdd out_state_main[1] DFFNEGX1_136/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3678 gnd out_state_main[1] DFFNEGX1_136/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3679 DFFNEGX1_136/a_61_6# DFFNEGX1_136/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3680 DFFNEGX1_136/a_76_84# DFFNEGX1_136/a_2_6# DFFNEGX1_136/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3681 out_state_main[1] DFFNEGX1_136/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3682 vdd INVX2_259/Y DFFNEGX1_136/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3683 DFFNEGX1_136/a_31_6# DFFNEGX1_136/a_2_6# DFFNEGX1_136/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3684 DFFNEGX1_136/a_66_6# INVX2_259/Y DFFNEGX1_136/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3685 DFFNEGX1_136/a_17_74# INVX2_120/A vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3686 DFFNEGX1_136/a_31_74# INVX2_259/Y DFFNEGX1_136/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3687 DFFNEGX1_136/a_17_6# INVX2_120/A gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3688 gnd OAI22X1_52/Y OAI21X1_130/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M3689 vdd INVX2_52/A OAI21X1_130/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M3690 OAI21X1_130/Y INVX2_52/A OAI21X1_130/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3691 OAI21X1_130/Y OAI22X1_51/Y OAI21X1_130/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3692 OAI21X1_130/a_9_54# OAI22X1_52/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3693 OAI21X1_130/a_2_6# OAI22X1_51/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3694 gnd OAI22X1_66/Y OAI21X1_141/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M3695 vdd INVX2_38/Y AOI21X1_15/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M3696 AOI21X1_15/B INVX2_38/Y OAI21X1_141/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3697 AOI21X1_15/B OAI22X1_65/Y OAI21X1_141/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3698 OAI21X1_141/a_9_54# OAI22X1_66/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3699 OAI21X1_141/a_2_6# OAI22X1_65/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3700 gnd out_global_score[27] AOI22X1_6/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M3701 INVX2_189/A INVX2_258/Y AOI22X1_6/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3702 AOI22X1_6/a_11_6# HAX1_3/YS gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3703 AOI22X1_6/a_2_54# INVX2_258/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M3704 AOI22X1_6/a_28_6# INVX2_255/Y INVX2_189/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3705 vdd HAX1_3/YS AOI22X1_6/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3706 INVX2_189/A INVX2_255/Y AOI22X1_6/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M3707 AOI22X1_6/a_2_54# out_global_score[27] INVX2_189/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3708 gnd OAI22X1_84/Y OAI21X1_152/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M3709 vdd XOR2X1_4/Y AOI21X1_18/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M3710 AOI21X1_18/A XOR2X1_4/Y OAI21X1_152/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3711 AOI21X1_18/A OAI22X1_83/Y OAI21X1_152/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3712 OAI21X1_152/a_9_54# OAI22X1_84/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3713 OAI21X1_152/a_2_6# OAI22X1_83/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3714 OAI21X1_5/C out_mines[23] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M3715 NAND2X1_16/a_9_6# out_mines[23] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3716 vdd OAI21X1_5/A OAI21X1_5/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3717 OAI21X1_5/C OAI21X1_5/A NAND2X1_16/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3718 OAI21X1_54/C out_temp_index[3] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M3719 NAND2X1_49/a_9_6# out_temp_index[3] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3720 vdd NOR2X1_67/Y OAI21X1_54/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3721 OAI21X1_54/C NOR2X1_67/Y NAND2X1_49/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3722 OAI21X1_8/A NAND3X1_7/C vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M3723 NAND2X1_38/a_9_6# NAND3X1_7/C gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3724 vdd NOR2X1_66/Y OAI21X1_8/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3725 OAI21X1_8/A NOR2X1_66/Y NAND2X1_38/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3726 OAI21X1_23/C out_mines[14] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M3727 NAND2X1_27/a_9_6# out_mines[14] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3728 vdd INVX2_230/Y OAI21X1_23/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3729 OAI21X1_23/C INVX2_230/Y NAND2X1_27/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3730 gnd out_global_score[19] AOI22X1_14/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M3731 INVX2_197/A INVX2_257/Y AOI22X1_14/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3732 AOI22X1_14/a_11_6# HAX1_11/YS gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3733 AOI22X1_14/a_2_54# INVX2_257/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M3734 AOI22X1_14/a_28_6# INVX2_255/Y INVX2_197/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3735 vdd HAX1_11/YS AOI22X1_14/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3736 INVX2_197/A INVX2_255/Y AOI22X1_14/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M3737 AOI22X1_14/a_2_54# out_global_score[19] INVX2_197/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3738 gnd out_global_score[8] AOI22X1_25/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M3739 INVX2_208/A INVX2_258/Y AOI22X1_25/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3740 AOI22X1_25/a_11_6# HAX1_22/YS gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3741 AOI22X1_25/a_2_54# INVX2_258/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M3742 AOI22X1_25/a_28_6# OR2X1_11/B INVX2_208/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3743 vdd HAX1_22/YS AOI22X1_25/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3744 INVX2_208/A OR2X1_11/B AOI22X1_25/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M3745 AOI22X1_25/a_2_54# out_global_score[8] INVX2_208/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3746 gnd out_temp_decoded[7] AOI22X1_36/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M3747 OAI21X1_66/C out_mines[6] AOI22X1_36/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3748 AOI22X1_36/a_11_6# out_temp_decoded[6] gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3749 AOI22X1_36/a_2_54# out_mines[6] vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M3750 AOI22X1_36/a_28_6# out_mines[7] OAI21X1_66/C Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3751 vdd out_temp_decoded[6] AOI22X1_36/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3752 OAI21X1_66/C out_mines[7] AOI22X1_36/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M3753 AOI22X1_36/a_2_54# out_temp_decoded[7] OAI21X1_66/C vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3754 gnd NOR2X1_95/Y AOI22X1_47/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M3755 NAND3X1_41/A INVX2_14/Y AOI22X1_47/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3756 AOI22X1_47/a_11_6# NOR2X1_96/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3757 AOI22X1_47/a_2_54# INVX2_14/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M3758 AOI22X1_47/a_28_6# INVX2_12/Y NAND3X1_41/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3759 vdd NOR2X1_96/Y AOI22X1_47/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3760 NAND3X1_41/A INVX2_12/Y AOI22X1_47/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M3761 AOI22X1_47/a_2_54# NOR2X1_95/Y NAND3X1_41/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3762 gnd INVX2_31/Y AOI22X1_58/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M3763 OAI22X1_40/D out_mines[10] AOI22X1_58/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3764 AOI22X1_58/a_11_6# INVX2_32/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3765 AOI22X1_58/a_2_54# out_mines[10] vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M3766 AOI22X1_58/a_28_6# out_mines[18] OAI22X1_40/D Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3767 vdd INVX2_32/Y AOI22X1_58/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3768 OAI22X1_40/D out_mines[18] AOI22X1_58/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M3769 AOI22X1_58/a_2_54# INVX2_31/Y OAI22X1_40/D vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3770 gnd NOR2X1_113/Y AOI22X1_69/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M3771 AND2X2_16/A AOI22X1_69/B AOI22X1_69/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3772 AOI22X1_69/a_11_6# NOR2X1_114/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3773 AOI22X1_69/a_2_54# AOI22X1_69/B vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M3774 AOI22X1_69/a_28_6# AOI21X1_8/B AND2X2_16/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3775 vdd NOR2X1_114/Y AOI22X1_69/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3776 AND2X2_16/A AOI21X1_8/B AOI22X1_69/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M3777 AOI22X1_69/a_2_54# NOR2X1_113/Y AND2X2_16/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3778 gnd BUFX2_25/Y OAI22X1_9/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M3779 OAI22X1_9/a_2_6# OR2X1_11/A OAI22X1_9/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M3780 OAI22X1_9/Y INVX2_61/Y OAI22X1_9/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3781 OAI22X1_9/Y INVX2_94/Y OAI22X1_9/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M3782 OAI22X1_9/a_28_54# INVX2_61/Y OAI22X1_9/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3783 OAI22X1_9/a_9_54# BUFX2_25/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3784 OAI22X1_9/a_2_6# INVX2_94/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3785 vdd OR2X1_11/A OAI22X1_9/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3786 INVX2_18/Y out_mines[23] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3787 INVX2_18/Y out_mines[23] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3788 INVX2_29/Y out_temp_mine_cnt[0] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3789 INVX2_29/Y out_temp_mine_cnt[0] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3790 gnd XOR2X1_1/A XOR2X1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3791 XOR2X1_1/Y XOR2X1_1/a_2_6# XOR2X1_1/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3792 XOR2X1_1/a_13_43# out_temp_mine_cnt[4] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3793 XOR2X1_1/a_18_54# XOR2X1_1/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3794 XOR2X1_1/a_35_6# XOR2X1_1/A XOR2X1_1/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3795 XOR2X1_1/a_18_6# XOR2X1_1/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3796 vdd XOR2X1_1/A XOR2X1_1/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3797 vdd out_temp_mine_cnt[4] XOR2X1_1/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3798 XOR2X1_1/Y XOR2X1_1/A XOR2X1_1/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3799 XOR2X1_1/a_35_54# XOR2X1_1/a_2_6# XOR2X1_1/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3800 XOR2X1_1/a_13_43# out_temp_mine_cnt[4] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3801 gnd out_temp_mine_cnt[4] XOR2X1_1/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3802 gnd MUX2X1_2/A MUX2X1_2/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M3803 MUX2X1_2/a_17_50# XOR2X1_6/Y vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3804 MUX2X1_2/Y NOR2X1_7/Y MUX2X1_2/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M3805 MUX2X1_2/a_30_54# MUX2X1_2/a_2_10# MUX2X1_2/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3806 MUX2X1_2/a_17_10# XOR2X1_6/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3807 vdd NOR2X1_7/Y MUX2X1_2/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3808 MUX2X1_2/a_30_10# NOR2X1_7/Y MUX2X1_2/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M3809 gnd NOR2X1_7/Y MUX2X1_2/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M3810 vdd MUX2X1_2/A MUX2X1_2/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3811 MUX2X1_2/Y MUX2X1_2/a_2_10# MUX2X1_2/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3812 MUX2X1_19/A FAX1_1/YS gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3813 MUX2X1_19/A FAX1_1/YS vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3814 INVX2_130/Y out_start gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3815 INVX2_130/Y out_start vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3816 HAX1_45/A MUX2X1_16/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3817 HAX1_45/A MUX2X1_16/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3818 OR2X1_4/A MUX2X1_5/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3819 OR2X1_4/A MUX2X1_5/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3820 MUX2X1_32/B XNOR2X1_1/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3821 MUX2X1_32/B XNOR2X1_1/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3822 INVX2_196/Y INVX2_196/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3823 INVX2_196/Y INVX2_196/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3824 INVX2_185/Y INVX2_185/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3825 INVX2_185/Y INVX2_185/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3826 DFFNEGX1_25/a_76_6# BUFX2_16/Y DFFNEGX1_25/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3827 gnd BUFX2_16/Y DFFNEGX1_25/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3828 DFFNEGX1_25/a_66_6# DFFNEGX1_25/a_2_6# DFFNEGX1_25/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3829 out_mines[19] DFFNEGX1_25/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3830 DFFNEGX1_25/a_23_6# BUFX2_16/Y DFFNEGX1_25/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3831 DFFNEGX1_25/a_23_6# DFFNEGX1_25/a_2_6# DFFNEGX1_25/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3832 gnd DFFNEGX1_25/a_34_4# DFFNEGX1_25/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3833 vdd DFFNEGX1_25/a_34_4# DFFNEGX1_25/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3834 DFFNEGX1_25/a_61_74# DFFNEGX1_25/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3835 DFFNEGX1_25/a_34_4# DFFNEGX1_25/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3836 DFFNEGX1_25/a_34_4# DFFNEGX1_25/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3837 vdd out_mines[19] DFFNEGX1_25/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3838 gnd out_mines[19] DFFNEGX1_25/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3839 DFFNEGX1_25/a_61_6# DFFNEGX1_25/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3840 DFFNEGX1_25/a_76_84# DFFNEGX1_25/a_2_6# DFFNEGX1_25/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3841 out_mines[19] DFFNEGX1_25/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3842 vdd BUFX2_16/Y DFFNEGX1_25/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3843 DFFNEGX1_25/a_31_6# DFFNEGX1_25/a_2_6# DFFNEGX1_25/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3844 DFFNEGX1_25/a_66_6# BUFX2_16/Y DFFNEGX1_25/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3845 DFFNEGX1_25/a_17_74# OAI21X1_13/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3846 DFFNEGX1_25/a_31_74# BUFX2_16/Y DFFNEGX1_25/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3847 DFFNEGX1_25/a_17_6# OAI21X1_13/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3848 DFFNEGX1_14/a_76_6# BUFX2_16/Y DFFNEGX1_14/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3849 gnd BUFX2_16/Y DFFNEGX1_14/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3850 DFFNEGX1_14/a_66_6# DFFNEGX1_14/a_2_6# DFFNEGX1_14/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3851 out_mines[12] DFFNEGX1_14/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3852 DFFNEGX1_14/a_23_6# BUFX2_16/Y DFFNEGX1_14/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3853 DFFNEGX1_14/a_23_6# DFFNEGX1_14/a_2_6# DFFNEGX1_14/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3854 gnd DFFNEGX1_14/a_34_4# DFFNEGX1_14/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3855 vdd DFFNEGX1_14/a_34_4# DFFNEGX1_14/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3856 DFFNEGX1_14/a_61_74# DFFNEGX1_14/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3857 DFFNEGX1_14/a_34_4# DFFNEGX1_14/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3858 DFFNEGX1_14/a_34_4# DFFNEGX1_14/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3859 vdd out_mines[12] DFFNEGX1_14/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3860 gnd out_mines[12] DFFNEGX1_14/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3861 DFFNEGX1_14/a_61_6# DFFNEGX1_14/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3862 DFFNEGX1_14/a_76_84# DFFNEGX1_14/a_2_6# DFFNEGX1_14/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3863 out_mines[12] DFFNEGX1_14/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3864 vdd BUFX2_16/Y DFFNEGX1_14/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3865 DFFNEGX1_14/a_31_6# DFFNEGX1_14/a_2_6# DFFNEGX1_14/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3866 DFFNEGX1_14/a_66_6# BUFX2_16/Y DFFNEGX1_14/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3867 DFFNEGX1_14/a_17_74# OAI21X1_27/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3868 DFFNEGX1_14/a_31_74# BUFX2_16/Y DFFNEGX1_14/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3869 DFFNEGX1_14/a_17_6# OAI21X1_27/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3870 DFFNEGX1_58/a_76_6# BUFX2_13/Y DFFNEGX1_58/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3871 gnd BUFX2_13/Y DFFNEGX1_58/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3872 DFFNEGX1_58/a_66_6# DFFNEGX1_58/a_2_6# DFFNEGX1_58/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3873 out_temp_decoded[8] DFFNEGX1_58/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3874 DFFNEGX1_58/a_23_6# BUFX2_13/Y DFFNEGX1_58/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3875 DFFNEGX1_58/a_23_6# DFFNEGX1_58/a_2_6# DFFNEGX1_58/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3876 gnd DFFNEGX1_58/a_34_4# DFFNEGX1_58/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3877 vdd DFFNEGX1_58/a_34_4# DFFNEGX1_58/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3878 DFFNEGX1_58/a_61_74# DFFNEGX1_58/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3879 DFFNEGX1_58/a_34_4# DFFNEGX1_58/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3880 DFFNEGX1_58/a_34_4# DFFNEGX1_58/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3881 vdd out_temp_decoded[8] DFFNEGX1_58/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3882 gnd out_temp_decoded[8] DFFNEGX1_58/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3883 DFFNEGX1_58/a_61_6# DFFNEGX1_58/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3884 DFFNEGX1_58/a_76_84# DFFNEGX1_58/a_2_6# DFFNEGX1_58/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3885 out_temp_decoded[8] DFFNEGX1_58/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3886 vdd BUFX2_13/Y DFFNEGX1_58/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3887 DFFNEGX1_58/a_31_6# DFFNEGX1_58/a_2_6# DFFNEGX1_58/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3888 DFFNEGX1_58/a_66_6# BUFX2_13/Y DFFNEGX1_58/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3889 DFFNEGX1_58/a_17_74# OAI21X1_90/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3890 DFFNEGX1_58/a_31_74# BUFX2_13/Y DFFNEGX1_58/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3891 DFFNEGX1_58/a_17_6# OAI21X1_90/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3892 DFFNEGX1_47/a_76_6# BUFX2_14/Y DFFNEGX1_47/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3893 gnd BUFX2_14/Y DFFNEGX1_47/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3894 DFFNEGX1_47/a_66_6# DFFNEGX1_47/a_2_6# DFFNEGX1_47/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3895 out_temp_decoded[19] DFFNEGX1_47/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3896 DFFNEGX1_47/a_23_6# BUFX2_14/Y DFFNEGX1_47/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3897 DFFNEGX1_47/a_23_6# DFFNEGX1_47/a_2_6# DFFNEGX1_47/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3898 gnd DFFNEGX1_47/a_34_4# DFFNEGX1_47/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3899 vdd DFFNEGX1_47/a_34_4# DFFNEGX1_47/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3900 DFFNEGX1_47/a_61_74# DFFNEGX1_47/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3901 DFFNEGX1_47/a_34_4# DFFNEGX1_47/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3902 DFFNEGX1_47/a_34_4# DFFNEGX1_47/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3903 vdd out_temp_decoded[19] DFFNEGX1_47/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3904 gnd out_temp_decoded[19] DFFNEGX1_47/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3905 DFFNEGX1_47/a_61_6# DFFNEGX1_47/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3906 DFFNEGX1_47/a_76_84# DFFNEGX1_47/a_2_6# DFFNEGX1_47/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3907 out_temp_decoded[19] DFFNEGX1_47/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3908 vdd BUFX2_14/Y DFFNEGX1_47/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3909 DFFNEGX1_47/a_31_6# DFFNEGX1_47/a_2_6# DFFNEGX1_47/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3910 DFFNEGX1_47/a_66_6# BUFX2_14/Y DFFNEGX1_47/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3911 DFFNEGX1_47/a_17_74# OAI21X1_101/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3912 DFFNEGX1_47/a_31_74# BUFX2_14/Y DFFNEGX1_47/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3913 DFFNEGX1_47/a_17_6# OAI21X1_101/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3914 DFFNEGX1_36/a_76_6# INVX2_259/Y DFFNEGX1_36/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3915 gnd INVX2_259/Y DFFNEGX1_36/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3916 DFFNEGX1_36/a_66_6# DFFNEGX1_36/a_2_6# DFFNEGX1_36/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3917 out_place_done DFFNEGX1_36/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3918 DFFNEGX1_36/a_23_6# INVX2_259/Y DFFNEGX1_36/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3919 DFFNEGX1_36/a_23_6# DFFNEGX1_36/a_2_6# DFFNEGX1_36/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3920 gnd DFFNEGX1_36/a_34_4# DFFNEGX1_36/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3921 vdd DFFNEGX1_36/a_34_4# DFFNEGX1_36/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3922 DFFNEGX1_36/a_61_74# DFFNEGX1_36/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3923 DFFNEGX1_36/a_34_4# DFFNEGX1_36/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3924 DFFNEGX1_36/a_34_4# DFFNEGX1_36/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3925 vdd out_place_done DFFNEGX1_36/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3926 gnd out_place_done DFFNEGX1_36/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3927 DFFNEGX1_36/a_61_6# DFFNEGX1_36/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3928 DFFNEGX1_36/a_76_84# DFFNEGX1_36/a_2_6# DFFNEGX1_36/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3929 out_place_done DFFNEGX1_36/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3930 vdd INVX2_259/Y DFFNEGX1_36/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3931 DFFNEGX1_36/a_31_6# DFFNEGX1_36/a_2_6# DFFNEGX1_36/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3932 DFFNEGX1_36/a_66_6# INVX2_259/Y DFFNEGX1_36/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3933 DFFNEGX1_36/a_17_74# NAND2X1_14/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3934 DFFNEGX1_36/a_31_74# INVX2_259/Y DFFNEGX1_36/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3935 DFFNEGX1_36/a_17_6# NAND2X1_14/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3936 DFFNEGX1_69/a_76_6# BUFX2_12/Y DFFNEGX1_69/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3937 gnd BUFX2_12/Y DFFNEGX1_69/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3938 DFFNEGX1_69/a_66_6# DFFNEGX1_69/a_2_6# DFFNEGX1_69/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3939 out_temp_cleared[22] DFFNEGX1_69/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3940 DFFNEGX1_69/a_23_6# BUFX2_12/Y DFFNEGX1_69/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3941 DFFNEGX1_69/a_23_6# DFFNEGX1_69/a_2_6# DFFNEGX1_69/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3942 gnd DFFNEGX1_69/a_34_4# DFFNEGX1_69/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3943 vdd DFFNEGX1_69/a_34_4# DFFNEGX1_69/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3944 DFFNEGX1_69/a_61_74# DFFNEGX1_69/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3945 DFFNEGX1_69/a_34_4# DFFNEGX1_69/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3946 DFFNEGX1_69/a_34_4# DFFNEGX1_69/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3947 vdd out_temp_cleared[22] DFFNEGX1_69/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3948 gnd out_temp_cleared[22] DFFNEGX1_69/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3949 DFFNEGX1_69/a_61_6# DFFNEGX1_69/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3950 DFFNEGX1_69/a_76_84# DFFNEGX1_69/a_2_6# DFFNEGX1_69/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M3951 out_temp_cleared[22] DFFNEGX1_69/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3952 vdd BUFX2_12/Y DFFNEGX1_69/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3953 DFFNEGX1_69/a_31_6# DFFNEGX1_69/a_2_6# DFFNEGX1_69/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3954 DFFNEGX1_69/a_66_6# BUFX2_12/Y DFFNEGX1_69/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3955 DFFNEGX1_69/a_17_74# OAI22X1_6/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3956 DFFNEGX1_69/a_31_74# BUFX2_12/Y DFFNEGX1_69/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3957 DFFNEGX1_69/a_17_6# OAI22X1_6/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M3958 gnd out_temp_data_in[4] XOR2X1_12/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3959 XOR2X1_12/Y XOR2X1_12/a_2_6# XOR2X1_12/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3960 XOR2X1_12/a_13_43# OR2X1_10/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3961 XOR2X1_12/a_18_54# XOR2X1_12/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3962 XOR2X1_12/a_35_6# out_temp_data_in[4] XOR2X1_12/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3963 XOR2X1_12/a_18_6# XOR2X1_12/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3964 vdd out_temp_data_in[4] XOR2X1_12/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3965 vdd OR2X1_10/Y XOR2X1_12/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3966 XOR2X1_12/Y out_temp_data_in[4] XOR2X1_12/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3967 XOR2X1_12/a_35_54# XOR2X1_12/a_2_6# XOR2X1_12/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3968 XOR2X1_12/a_13_43# OR2X1_10/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3969 gnd OR2X1_10/Y XOR2X1_12/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3970 gnd XOR2X1_23/A XOR2X1_23/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3971 XOR2X1_23/Y XOR2X1_23/a_2_6# XOR2X1_23/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M3972 XOR2X1_23/a_13_43# XOR2X1_23/B gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3973 XOR2X1_23/a_18_54# XOR2X1_23/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M3974 XOR2X1_23/a_35_6# XOR2X1_23/A XOR2X1_23/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3975 XOR2X1_23/a_18_6# XOR2X1_23/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3976 vdd XOR2X1_23/A XOR2X1_23/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M3977 vdd XOR2X1_23/B XOR2X1_23/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M3978 XOR2X1_23/Y XOR2X1_23/A XOR2X1_23/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M3979 XOR2X1_23/a_35_54# XOR2X1_23/a_2_6# XOR2X1_23/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M3980 XOR2X1_23/a_13_43# XOR2X1_23/B vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M3981 gnd XOR2X1_23/B XOR2X1_23/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3982 NOR2X1_52/B OAI21X1_1/B vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M3983 NAND3X1_2/a_9_6# OAI21X1_1/B gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M3984 NOR2X1_52/B out_temp_data_in[4] vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3985 NOR2X1_52/B out_temp_data_in[4] NAND3X1_2/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M3986 vdd OAI21X1_1/A NOR2X1_52/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M3987 NAND3X1_2/a_14_6# OAI21X1_1/A NAND3X1_2/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M3988 DFFNEGX1_104/a_76_6# BUFX2_10/Y DFFNEGX1_104/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M3989 gnd BUFX2_10/Y DFFNEGX1_104/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M3990 DFFNEGX1_104/a_66_6# DFFNEGX1_104/a_2_6# DFFNEGX1_104/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3991 out_global_score[10] DFFNEGX1_104/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3992 DFFNEGX1_104/a_23_6# BUFX2_10/Y DFFNEGX1_104/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M3993 DFFNEGX1_104/a_23_6# DFFNEGX1_104/a_2_6# DFFNEGX1_104/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M3994 gnd DFFNEGX1_104/a_34_4# DFFNEGX1_104/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M3995 vdd DFFNEGX1_104/a_34_4# DFFNEGX1_104/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M3996 DFFNEGX1_104/a_61_74# DFFNEGX1_104/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M3997 DFFNEGX1_104/a_34_4# DFFNEGX1_104/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M3998 DFFNEGX1_104/a_34_4# DFFNEGX1_104/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M3999 vdd out_global_score[10] DFFNEGX1_104/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4000 gnd out_global_score[10] DFFNEGX1_104/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4001 DFFNEGX1_104/a_61_6# DFFNEGX1_104/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4002 DFFNEGX1_104/a_76_84# DFFNEGX1_104/a_2_6# DFFNEGX1_104/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M4003 out_global_score[10] DFFNEGX1_104/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4004 vdd BUFX2_10/Y DFFNEGX1_104/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4005 DFFNEGX1_104/a_31_6# DFFNEGX1_104/a_2_6# DFFNEGX1_104/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4006 DFFNEGX1_104/a_66_6# BUFX2_10/Y DFFNEGX1_104/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4007 DFFNEGX1_104/a_17_74# INVX2_206/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4008 DFFNEGX1_104/a_31_74# BUFX2_10/Y DFFNEGX1_104/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4009 DFFNEGX1_104/a_17_6# INVX2_206/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4010 DFFNEGX1_115/a_76_6# BUFX2_9/Y DFFNEGX1_115/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M4011 gnd BUFX2_9/Y DFFNEGX1_115/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4012 DFFNEGX1_115/a_66_6# DFFNEGX1_115/a_2_6# DFFNEGX1_115/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4013 out_global_score[21] DFFNEGX1_115/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4014 DFFNEGX1_115/a_23_6# BUFX2_9/Y DFFNEGX1_115/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M4015 DFFNEGX1_115/a_23_6# DFFNEGX1_115/a_2_6# DFFNEGX1_115/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M4016 gnd DFFNEGX1_115/a_34_4# DFFNEGX1_115/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4017 vdd DFFNEGX1_115/a_34_4# DFFNEGX1_115/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M4018 DFFNEGX1_115/a_61_74# DFFNEGX1_115/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4019 DFFNEGX1_115/a_34_4# DFFNEGX1_115/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4020 DFFNEGX1_115/a_34_4# DFFNEGX1_115/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4021 vdd out_global_score[21] DFFNEGX1_115/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4022 gnd out_global_score[21] DFFNEGX1_115/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4023 DFFNEGX1_115/a_61_6# DFFNEGX1_115/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4024 DFFNEGX1_115/a_76_84# DFFNEGX1_115/a_2_6# DFFNEGX1_115/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M4025 out_global_score[21] DFFNEGX1_115/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4026 vdd BUFX2_9/Y DFFNEGX1_115/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4027 DFFNEGX1_115/a_31_6# DFFNEGX1_115/a_2_6# DFFNEGX1_115/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4028 DFFNEGX1_115/a_66_6# BUFX2_9/Y DFFNEGX1_115/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4029 DFFNEGX1_115/a_17_74# INVX2_195/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4030 DFFNEGX1_115/a_31_74# BUFX2_9/Y DFFNEGX1_115/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4031 DFFNEGX1_115/a_17_6# INVX2_195/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4032 DFFNEGX1_126/a_76_6# BUFX2_5/Y DFFNEGX1_126/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M4033 gnd BUFX2_5/Y DFFNEGX1_126/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4034 DFFNEGX1_126/a_66_6# DFFNEGX1_126/a_2_6# DFFNEGX1_126/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4035 out_n_nearby[1] DFFNEGX1_126/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4036 DFFNEGX1_126/a_23_6# BUFX2_5/Y DFFNEGX1_126/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M4037 DFFNEGX1_126/a_23_6# DFFNEGX1_126/a_2_6# DFFNEGX1_126/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M4038 gnd DFFNEGX1_126/a_34_4# DFFNEGX1_126/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4039 vdd DFFNEGX1_126/a_34_4# DFFNEGX1_126/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M4040 DFFNEGX1_126/a_61_74# DFFNEGX1_126/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4041 DFFNEGX1_126/a_34_4# DFFNEGX1_126/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4042 DFFNEGX1_126/a_34_4# DFFNEGX1_126/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4043 vdd out_n_nearby[1] DFFNEGX1_126/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4044 gnd out_n_nearby[1] DFFNEGX1_126/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4045 DFFNEGX1_126/a_61_6# DFFNEGX1_126/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4046 DFFNEGX1_126/a_76_84# DFFNEGX1_126/a_2_6# DFFNEGX1_126/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M4047 out_n_nearby[1] DFFNEGX1_126/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4048 vdd BUFX2_5/Y DFFNEGX1_126/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4049 DFFNEGX1_126/a_31_6# DFFNEGX1_126/a_2_6# DFFNEGX1_126/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4050 DFFNEGX1_126/a_66_6# BUFX2_5/Y DFFNEGX1_126/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4051 DFFNEGX1_126/a_17_74# OAI21X1_62/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4052 DFFNEGX1_126/a_31_74# BUFX2_5/Y DFFNEGX1_126/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4053 DFFNEGX1_126/a_17_6# OAI21X1_62/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4054 DFFNEGX1_137/a_76_6# BUFX2_5/Y DFFNEGX1_137/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M4055 gnd BUFX2_5/Y DFFNEGX1_137/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4056 DFFNEGX1_137/a_66_6# DFFNEGX1_137/a_2_6# DFFNEGX1_137/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4057 INVX2_127/A DFFNEGX1_137/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4058 DFFNEGX1_137/a_23_6# BUFX2_5/Y DFFNEGX1_137/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M4059 DFFNEGX1_137/a_23_6# DFFNEGX1_137/a_2_6# DFFNEGX1_137/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M4060 gnd DFFNEGX1_137/a_34_4# DFFNEGX1_137/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4061 vdd DFFNEGX1_137/a_34_4# DFFNEGX1_137/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M4062 DFFNEGX1_137/a_61_74# DFFNEGX1_137/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4063 DFFNEGX1_137/a_34_4# DFFNEGX1_137/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4064 DFFNEGX1_137/a_34_4# DFFNEGX1_137/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4065 vdd INVX2_127/A DFFNEGX1_137/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4066 gnd INVX2_127/A DFFNEGX1_137/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4067 DFFNEGX1_137/a_61_6# DFFNEGX1_137/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4068 DFFNEGX1_137/a_76_84# DFFNEGX1_137/a_2_6# DFFNEGX1_137/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M4069 INVX2_127/A DFFNEGX1_137/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4070 vdd BUFX2_5/Y DFFNEGX1_137/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4071 DFFNEGX1_137/a_31_6# DFFNEGX1_137/a_2_6# DFFNEGX1_137/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4072 DFFNEGX1_137/a_66_6# BUFX2_5/Y DFFNEGX1_137/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4073 DFFNEGX1_137/a_17_74# AOI21X1_24/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4074 DFFNEGX1_137/a_31_74# BUFX2_5/Y DFFNEGX1_137/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4075 DFFNEGX1_137/a_17_6# AOI21X1_24/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4076 gnd INVX2_19/Y OAI21X1_120/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M4077 vdd AOI22X1_68/Y INVX2_33/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M4078 INVX2_33/A AOI22X1_68/Y OAI21X1_120/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4079 INVX2_33/A NOR2X1_110/B OAI21X1_120/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4080 OAI21X1_120/a_9_54# INVX2_19/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4081 OAI21X1_120/a_2_6# NOR2X1_110/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4082 gnd AOI22X1_73/Y OAI21X1_131/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M4083 vdd OAI21X1_132/Y XOR2X1_29/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M4084 XOR2X1_29/B OAI21X1_132/Y OAI21X1_131/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4085 XOR2X1_29/B XOR2X1_13/Y OAI21X1_131/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4086 OAI21X1_131/a_9_54# AOI22X1_73/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4087 OAI21X1_131/a_2_6# XOR2X1_13/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4088 gnd out_global_score[26] AOI22X1_7/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M4089 INVX2_190/A INVX2_257/Y AOI22X1_7/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M4090 AOI22X1_7/a_11_6# HAX1_4/YS gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4091 AOI22X1_7/a_2_54# INVX2_257/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M4092 AOI22X1_7/a_28_6# INVX2_255/Y INVX2_190/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4093 vdd HAX1_4/YS AOI22X1_7/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4094 INVX2_190/A INVX2_255/Y AOI22X1_7/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M4095 AOI22X1_7/a_2_54# out_global_score[26] INVX2_190/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4096 gnd OAI22X1_86/Y OAI21X1_153/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M4097 vdd INVX2_35/Y OAI21X1_153/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M4098 OAI21X1_153/Y INVX2_35/Y OAI21X1_153/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4099 OAI21X1_153/Y OAI22X1_85/Y OAI21X1_153/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4100 OAI21X1_153/a_9_54# OAI22X1_86/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4101 OAI21X1_153/a_2_6# OAI22X1_85/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4102 gnd OAI22X1_68/Y OAI21X1_142/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M4103 vdd XOR2X1_3/Y AOI21X1_15/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M4104 AOI21X1_15/A XOR2X1_3/Y OAI21X1_142/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4105 AOI21X1_15/A OAI22X1_67/Y OAI21X1_142/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4106 OAI21X1_142/a_9_54# OAI22X1_68/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4107 OAI21X1_142/a_2_6# OAI22X1_67/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4108 OAI21X1_7/C out_mines[22] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M4109 NAND2X1_17/a_9_6# out_mines[22] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4110 vdd OAI21X1_7/A OAI21X1_7/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4111 OAI21X1_7/C OAI21X1_7/A NAND2X1_17/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4112 OAI21X1_41/C out_mines[5] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M4113 NAND2X1_39/a_9_6# out_mines[5] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4114 vdd INVX2_237/Y OAI21X1_41/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4115 OAI21X1_41/C INVX2_237/Y NAND2X1_39/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4116 OAI21X1_25/C out_mines[13] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M4117 NAND2X1_28/a_9_6# out_mines[13] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4118 vdd INVX2_235/Y OAI21X1_25/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4119 OAI21X1_25/C INVX2_235/Y NAND2X1_28/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4120 gnd out_global_score[18] AOI22X1_15/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M4121 INVX2_198/A INVX2_257/Y AOI22X1_15/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M4122 AOI22X1_15/a_11_6# HAX1_12/YS gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4123 AOI22X1_15/a_2_54# INVX2_257/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M4124 AOI22X1_15/a_28_6# OR2X1_11/B INVX2_198/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4125 vdd HAX1_12/YS AOI22X1_15/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4126 INVX2_198/A OR2X1_11/B AOI22X1_15/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M4127 AOI22X1_15/a_2_54# out_global_score[18] INVX2_198/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4128 gnd out_global_score[7] AOI22X1_26/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M4129 INVX2_209/A INVX2_258/Y AOI22X1_26/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M4130 AOI22X1_26/a_11_6# HAX1_23/YS gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4131 AOI22X1_26/a_2_54# INVX2_258/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M4132 AOI22X1_26/a_28_6# OR2X1_11/B INVX2_209/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4133 vdd HAX1_23/YS AOI22X1_26/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4134 INVX2_209/A OR2X1_11/B AOI22X1_26/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M4135 AOI22X1_26/a_2_54# out_global_score[7] INVX2_209/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4136 gnd out_temp_decoded[11] AOI22X1_37/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M4137 OAI21X1_67/C out_mines[10] AOI22X1_37/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M4138 AOI22X1_37/a_11_6# out_temp_decoded[10] gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4139 AOI22X1_37/a_2_54# out_mines[10] vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M4140 AOI22X1_37/a_28_6# out_mines[11] OAI21X1_67/C Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4141 vdd out_temp_decoded[10] AOI22X1_37/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4142 OAI21X1_67/C out_mines[11] AOI22X1_37/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M4143 AOI22X1_37/a_2_54# out_temp_decoded[11] OAI21X1_67/C vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4144 gnd out_temp_cleared[18] AOI22X1_48/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M4145 NAND3X1_44/B INVX2_21/Y AOI22X1_48/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M4146 AOI22X1_48/a_11_6# NOR2X1_99/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4147 AOI22X1_48/a_2_54# INVX2_21/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M4148 AOI22X1_48/a_28_6# out_mines[18] NAND3X1_44/B Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4149 vdd NOR2X1_99/Y AOI22X1_48/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4150 NAND3X1_44/B out_mines[18] AOI22X1_48/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M4151 AOI22X1_48/a_2_54# out_temp_cleared[18] NAND3X1_44/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4152 gnd out_temp_data_in[0] AOI22X1_59/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M4153 AOI22X1_59/Y INVX2_251/Y AOI22X1_59/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M4154 AOI22X1_59/a_11_6# AOI22X1_66/D gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4155 AOI22X1_59/a_2_54# INVX2_251/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M4156 AOI22X1_59/a_28_6# AOI22X1_69/B AOI22X1_59/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4157 vdd AOI22X1_66/D AOI22X1_59/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4158 AOI22X1_59/Y AOI22X1_69/B AOI22X1_59/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M4159 AOI22X1_59/a_2_54# out_temp_data_in[0] AOI22X1_59/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4160 vdd HAX1_40/A HAX1_40/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M4161 HAX1_40/a_41_74# HAX1_40/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M4162 HAX1_40/a_9_6# HAX1_40/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4163 HAX1_40/a_41_74# HAX1_40/B HAX1_40/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M4164 vdd HAX1_40/A HAX1_40/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4165 vdd HAX1_40/a_2_74# HAX1_41/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4166 HAX1_40/a_38_6# HAX1_40/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4167 HAX1_40/YS HAX1_40/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4168 HAX1_40/a_38_6# HAX1_40/A HAX1_40/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4169 HAX1_40/YS HAX1_40/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4170 HAX1_40/a_2_74# HAX1_40/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4171 HAX1_40/a_2_74# HAX1_40/B HAX1_40/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4172 HAX1_40/a_49_54# HAX1_40/B HAX1_40/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4173 gnd HAX1_40/a_2_74# HAX1_41/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M4174 INVX2_19/Y out_mines[21] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4175 INVX2_19/Y out_mines[21] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4176 gnd HAX1_0/YC XOR2X1_2/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4177 XOR2X1_2/Y XOR2X1_2/a_2_6# XOR2X1_2/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M4178 XOR2X1_2/a_13_43# out_global_score[31] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4179 XOR2X1_2/a_18_54# XOR2X1_2/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4180 XOR2X1_2/a_35_6# HAX1_0/YC XOR2X1_2/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4181 XOR2X1_2/a_18_6# XOR2X1_2/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4182 vdd HAX1_0/YC XOR2X1_2/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4183 vdd out_global_score[31] XOR2X1_2/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4184 XOR2X1_2/Y HAX1_0/YC XOR2X1_2/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M4185 XOR2X1_2/a_35_54# XOR2X1_2/a_2_6# XOR2X1_2/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4186 XOR2X1_2/a_13_43# out_global_score[31] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4187 gnd out_global_score[31] XOR2X1_2/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4188 gnd MUX2X1_3/A MUX2X1_3/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M4189 MUX2X1_3/a_17_50# XOR2X1_7/Y vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4190 MUX2X1_3/Y NOR2X1_7/Y MUX2X1_3/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M4191 MUX2X1_3/a_30_54# MUX2X1_3/a_2_10# MUX2X1_3/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4192 MUX2X1_3/a_17_10# XOR2X1_7/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4193 vdd NOR2X1_7/Y MUX2X1_3/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4194 MUX2X1_3/a_30_10# NOR2X1_7/Y MUX2X1_3/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M4195 gnd NOR2X1_7/Y MUX2X1_3/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M4196 vdd MUX2X1_3/A MUX2X1_3/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4197 MUX2X1_3/Y MUX2X1_3/a_2_10# MUX2X1_3/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4198 INVX2_120/Y INVX2_120/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4199 INVX2_120/Y INVX2_120/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4200 INVX2_131/Y out_decode gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4201 INVX2_131/Y out_decode vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4202 HAX1_44/A MUX2X1_17/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4203 HAX1_44/A MUX2X1_17/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4204 HAX1_41/A MUX2X1_6/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4205 HAX1_41/A MUX2X1_6/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4206 NOR2X1_0/A MUX2X1_29/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4207 NOR2X1_0/A MUX2X1_29/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4208 NOR2X1_32/B in_mult[4] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4209 NOR2X1_32/B in_mult[4] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4210 INVX2_197/Y INVX2_197/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4211 INVX2_197/Y INVX2_197/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4212 INVX2_186/Y INVX2_186/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4213 INVX2_186/Y INVX2_186/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4214 DFFNEGX1_15/a_76_6# BUFX2_16/Y DFFNEGX1_15/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M4215 gnd BUFX2_16/Y DFFNEGX1_15/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4216 DFFNEGX1_15/a_66_6# DFFNEGX1_15/a_2_6# DFFNEGX1_15/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4217 out_mines[8] DFFNEGX1_15/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4218 DFFNEGX1_15/a_23_6# BUFX2_16/Y DFFNEGX1_15/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M4219 DFFNEGX1_15/a_23_6# DFFNEGX1_15/a_2_6# DFFNEGX1_15/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M4220 gnd DFFNEGX1_15/a_34_4# DFFNEGX1_15/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4221 vdd DFFNEGX1_15/a_34_4# DFFNEGX1_15/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M4222 DFFNEGX1_15/a_61_74# DFFNEGX1_15/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4223 DFFNEGX1_15/a_34_4# DFFNEGX1_15/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4224 DFFNEGX1_15/a_34_4# DFFNEGX1_15/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4225 vdd out_mines[8] DFFNEGX1_15/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4226 gnd out_mines[8] DFFNEGX1_15/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4227 DFFNEGX1_15/a_61_6# DFFNEGX1_15/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4228 DFFNEGX1_15/a_76_84# DFFNEGX1_15/a_2_6# DFFNEGX1_15/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M4229 out_mines[8] DFFNEGX1_15/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4230 vdd BUFX2_16/Y DFFNEGX1_15/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4231 DFFNEGX1_15/a_31_6# DFFNEGX1_15/a_2_6# DFFNEGX1_15/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4232 DFFNEGX1_15/a_66_6# BUFX2_16/Y DFFNEGX1_15/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4233 DFFNEGX1_15/a_17_74# OAI21X1_35/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4234 DFFNEGX1_15/a_31_74# BUFX2_16/Y DFFNEGX1_15/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4235 DFFNEGX1_15/a_17_6# OAI21X1_35/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4236 DFFNEGX1_26/a_76_6# BUFX2_16/Y DFFNEGX1_26/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M4237 gnd BUFX2_16/Y DFFNEGX1_26/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4238 DFFNEGX1_26/a_66_6# DFFNEGX1_26/a_2_6# DFFNEGX1_26/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4239 out_mines[18] DFFNEGX1_26/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4240 DFFNEGX1_26/a_23_6# BUFX2_16/Y DFFNEGX1_26/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M4241 DFFNEGX1_26/a_23_6# DFFNEGX1_26/a_2_6# DFFNEGX1_26/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M4242 gnd DFFNEGX1_26/a_34_4# DFFNEGX1_26/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4243 vdd DFFNEGX1_26/a_34_4# DFFNEGX1_26/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M4244 DFFNEGX1_26/a_61_74# DFFNEGX1_26/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4245 DFFNEGX1_26/a_34_4# DFFNEGX1_26/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4246 DFFNEGX1_26/a_34_4# DFFNEGX1_26/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4247 vdd out_mines[18] DFFNEGX1_26/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4248 gnd out_mines[18] DFFNEGX1_26/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4249 DFFNEGX1_26/a_61_6# DFFNEGX1_26/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4250 DFFNEGX1_26/a_76_84# DFFNEGX1_26/a_2_6# DFFNEGX1_26/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M4251 out_mines[18] DFFNEGX1_26/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4252 vdd BUFX2_16/Y DFFNEGX1_26/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4253 DFFNEGX1_26/a_31_6# DFFNEGX1_26/a_2_6# DFFNEGX1_26/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4254 DFFNEGX1_26/a_66_6# BUFX2_16/Y DFFNEGX1_26/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4255 DFFNEGX1_26/a_17_74# OAI21X1_15/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4256 DFFNEGX1_26/a_31_74# BUFX2_16/Y DFFNEGX1_26/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4257 DFFNEGX1_26/a_17_6# OAI21X1_15/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4258 DFFNEGX1_59/a_76_6# BUFX2_13/Y DFFNEGX1_59/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M4259 gnd BUFX2_13/Y DFFNEGX1_59/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4260 DFFNEGX1_59/a_66_6# DFFNEGX1_59/a_2_6# DFFNEGX1_59/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4261 out_temp_decoded[7] DFFNEGX1_59/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4262 DFFNEGX1_59/a_23_6# BUFX2_13/Y DFFNEGX1_59/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M4263 DFFNEGX1_59/a_23_6# DFFNEGX1_59/a_2_6# DFFNEGX1_59/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M4264 gnd DFFNEGX1_59/a_34_4# DFFNEGX1_59/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4265 vdd DFFNEGX1_59/a_34_4# DFFNEGX1_59/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M4266 DFFNEGX1_59/a_61_74# DFFNEGX1_59/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4267 DFFNEGX1_59/a_34_4# DFFNEGX1_59/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4268 DFFNEGX1_59/a_34_4# DFFNEGX1_59/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4269 vdd out_temp_decoded[7] DFFNEGX1_59/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4270 gnd out_temp_decoded[7] DFFNEGX1_59/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4271 DFFNEGX1_59/a_61_6# DFFNEGX1_59/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4272 DFFNEGX1_59/a_76_84# DFFNEGX1_59/a_2_6# DFFNEGX1_59/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M4273 out_temp_decoded[7] DFFNEGX1_59/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4274 vdd BUFX2_13/Y DFFNEGX1_59/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4275 DFFNEGX1_59/a_31_6# DFFNEGX1_59/a_2_6# DFFNEGX1_59/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4276 DFFNEGX1_59/a_66_6# BUFX2_13/Y DFFNEGX1_59/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4277 DFFNEGX1_59/a_17_74# OAI21X1_89/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4278 DFFNEGX1_59/a_31_74# BUFX2_13/Y DFFNEGX1_59/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4279 DFFNEGX1_59/a_17_6# OAI21X1_89/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4280 DFFNEGX1_48/a_76_6# BUFX2_14/Y DFFNEGX1_48/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M4281 gnd BUFX2_14/Y DFFNEGX1_48/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4282 DFFNEGX1_48/a_66_6# DFFNEGX1_48/a_2_6# DFFNEGX1_48/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4283 out_temp_decoded[18] DFFNEGX1_48/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4284 DFFNEGX1_48/a_23_6# BUFX2_14/Y DFFNEGX1_48/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M4285 DFFNEGX1_48/a_23_6# DFFNEGX1_48/a_2_6# DFFNEGX1_48/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M4286 gnd DFFNEGX1_48/a_34_4# DFFNEGX1_48/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4287 vdd DFFNEGX1_48/a_34_4# DFFNEGX1_48/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M4288 DFFNEGX1_48/a_61_74# DFFNEGX1_48/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4289 DFFNEGX1_48/a_34_4# DFFNEGX1_48/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4290 DFFNEGX1_48/a_34_4# DFFNEGX1_48/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4291 vdd out_temp_decoded[18] DFFNEGX1_48/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4292 gnd out_temp_decoded[18] DFFNEGX1_48/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4293 DFFNEGX1_48/a_61_6# DFFNEGX1_48/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4294 DFFNEGX1_48/a_76_84# DFFNEGX1_48/a_2_6# DFFNEGX1_48/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M4295 out_temp_decoded[18] DFFNEGX1_48/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4296 vdd BUFX2_14/Y DFFNEGX1_48/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4297 DFFNEGX1_48/a_31_6# DFFNEGX1_48/a_2_6# DFFNEGX1_48/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4298 DFFNEGX1_48/a_66_6# BUFX2_14/Y DFFNEGX1_48/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4299 DFFNEGX1_48/a_17_74# OAI21X1_100/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4300 DFFNEGX1_48/a_31_74# BUFX2_14/Y DFFNEGX1_48/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4301 DFFNEGX1_48/a_17_6# OAI21X1_100/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4302 DFFNEGX1_37/a_76_6# BUFX2_15/Y DFFNEGX1_37/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M4303 gnd BUFX2_15/Y DFFNEGX1_37/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4304 DFFNEGX1_37/a_66_6# DFFNEGX1_37/a_2_6# DFFNEGX1_37/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4305 out_temp_data_in[4] DFFNEGX1_37/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4306 DFFNEGX1_37/a_23_6# BUFX2_15/Y DFFNEGX1_37/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M4307 DFFNEGX1_37/a_23_6# DFFNEGX1_37/a_2_6# DFFNEGX1_37/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M4308 gnd DFFNEGX1_37/a_34_4# DFFNEGX1_37/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4309 vdd DFFNEGX1_37/a_34_4# DFFNEGX1_37/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M4310 DFFNEGX1_37/a_61_74# DFFNEGX1_37/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4311 DFFNEGX1_37/a_34_4# DFFNEGX1_37/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4312 DFFNEGX1_37/a_34_4# DFFNEGX1_37/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4313 vdd out_temp_data_in[4] DFFNEGX1_37/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4314 gnd out_temp_data_in[4] DFFNEGX1_37/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4315 DFFNEGX1_37/a_61_6# DFFNEGX1_37/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4316 DFFNEGX1_37/a_76_84# DFFNEGX1_37/a_2_6# DFFNEGX1_37/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M4317 out_temp_data_in[4] DFFNEGX1_37/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4318 vdd BUFX2_15/Y DFFNEGX1_37/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4319 DFFNEGX1_37/a_31_6# DFFNEGX1_37/a_2_6# DFFNEGX1_37/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4320 DFFNEGX1_37/a_66_6# BUFX2_15/Y DFFNEGX1_37/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4321 DFFNEGX1_37/a_17_74# OAI21X1_111/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4322 DFFNEGX1_37/a_31_74# BUFX2_15/Y DFFNEGX1_37/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4323 DFFNEGX1_37/a_17_6# OAI21X1_111/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4324 gnd out_temp_data_in[4] XOR2X1_13/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4325 XOR2X1_13/Y XOR2X1_13/a_2_6# XOR2X1_13/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M4326 XOR2X1_13/a_13_43# OR2X1_7/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4327 XOR2X1_13/a_18_54# XOR2X1_13/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4328 XOR2X1_13/a_35_6# out_temp_data_in[4] XOR2X1_13/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4329 XOR2X1_13/a_18_6# XOR2X1_13/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4330 vdd out_temp_data_in[4] XOR2X1_13/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4331 vdd OR2X1_7/Y XOR2X1_13/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4332 XOR2X1_13/Y out_temp_data_in[4] XOR2X1_13/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M4333 XOR2X1_13/a_35_54# XOR2X1_13/a_2_6# XOR2X1_13/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4334 XOR2X1_13/a_13_43# OR2X1_7/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4335 gnd OR2X1_7/Y XOR2X1_13/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4336 gnd XOR2X1_24/A XOR2X1_24/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4337 XOR2X1_24/Y XOR2X1_24/a_2_6# XOR2X1_24/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M4338 XOR2X1_24/a_13_43# XOR2X1_25/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4339 XOR2X1_24/a_18_54# XOR2X1_24/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4340 XOR2X1_24/a_35_6# XOR2X1_24/A XOR2X1_24/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4341 XOR2X1_24/a_18_6# XOR2X1_24/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4342 vdd XOR2X1_24/A XOR2X1_24/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4343 vdd XOR2X1_25/Y XOR2X1_24/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4344 XOR2X1_24/Y XOR2X1_24/A XOR2X1_24/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M4345 XOR2X1_24/a_35_54# XOR2X1_24/a_2_6# XOR2X1_24/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4346 XOR2X1_24/a_13_43# XOR2X1_25/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4347 gnd XOR2X1_25/Y XOR2X1_24/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4348 NOR2X1_56/B out_temp_data_in[3] vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M4349 NAND3X1_3/a_9_6# out_temp_data_in[3] gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M4350 NOR2X1_56/B out_temp_data_in[2] vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4351 NOR2X1_56/B out_temp_data_in[2] NAND3X1_3/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M4352 vdd INVX2_30/Y NOR2X1_56/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4353 NAND3X1_3/a_14_6# INVX2_30/Y NAND3X1_3/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M4354 DFFNEGX1_105/a_76_6# BUFX2_10/Y DFFNEGX1_105/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M4355 gnd BUFX2_10/Y DFFNEGX1_105/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4356 DFFNEGX1_105/a_66_6# DFFNEGX1_105/a_2_6# DFFNEGX1_105/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4357 out_global_score[11] DFFNEGX1_105/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4358 DFFNEGX1_105/a_23_6# BUFX2_10/Y DFFNEGX1_105/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M4359 DFFNEGX1_105/a_23_6# DFFNEGX1_105/a_2_6# DFFNEGX1_105/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M4360 gnd DFFNEGX1_105/a_34_4# DFFNEGX1_105/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4361 vdd DFFNEGX1_105/a_34_4# DFFNEGX1_105/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M4362 DFFNEGX1_105/a_61_74# DFFNEGX1_105/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4363 DFFNEGX1_105/a_34_4# DFFNEGX1_105/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4364 DFFNEGX1_105/a_34_4# DFFNEGX1_105/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4365 vdd out_global_score[11] DFFNEGX1_105/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4366 gnd out_global_score[11] DFFNEGX1_105/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4367 DFFNEGX1_105/a_61_6# DFFNEGX1_105/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4368 DFFNEGX1_105/a_76_84# DFFNEGX1_105/a_2_6# DFFNEGX1_105/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M4369 out_global_score[11] DFFNEGX1_105/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4370 vdd BUFX2_10/Y DFFNEGX1_105/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4371 DFFNEGX1_105/a_31_6# DFFNEGX1_105/a_2_6# DFFNEGX1_105/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4372 DFFNEGX1_105/a_66_6# BUFX2_10/Y DFFNEGX1_105/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4373 DFFNEGX1_105/a_17_74# INVX2_205/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4374 DFFNEGX1_105/a_31_74# BUFX2_10/Y DFFNEGX1_105/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4375 DFFNEGX1_105/a_17_6# INVX2_205/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4376 DFFNEGX1_116/a_76_6# BUFX2_9/Y DFFNEGX1_116/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M4377 gnd BUFX2_9/Y DFFNEGX1_116/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4378 DFFNEGX1_116/a_66_6# DFFNEGX1_116/a_2_6# DFFNEGX1_116/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4379 out_global_score[22] DFFNEGX1_116/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4380 DFFNEGX1_116/a_23_6# BUFX2_9/Y DFFNEGX1_116/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M4381 DFFNEGX1_116/a_23_6# DFFNEGX1_116/a_2_6# DFFNEGX1_116/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M4382 gnd DFFNEGX1_116/a_34_4# DFFNEGX1_116/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4383 vdd DFFNEGX1_116/a_34_4# DFFNEGX1_116/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M4384 DFFNEGX1_116/a_61_74# DFFNEGX1_116/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4385 DFFNEGX1_116/a_34_4# DFFNEGX1_116/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4386 DFFNEGX1_116/a_34_4# DFFNEGX1_116/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4387 vdd out_global_score[22] DFFNEGX1_116/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4388 gnd out_global_score[22] DFFNEGX1_116/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4389 DFFNEGX1_116/a_61_6# DFFNEGX1_116/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4390 DFFNEGX1_116/a_76_84# DFFNEGX1_116/a_2_6# DFFNEGX1_116/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M4391 out_global_score[22] DFFNEGX1_116/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4392 vdd BUFX2_9/Y DFFNEGX1_116/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4393 DFFNEGX1_116/a_31_6# DFFNEGX1_116/a_2_6# DFFNEGX1_116/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4394 DFFNEGX1_116/a_66_6# BUFX2_9/Y DFFNEGX1_116/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4395 DFFNEGX1_116/a_17_74# INVX2_194/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4396 DFFNEGX1_116/a_31_74# BUFX2_9/Y DFFNEGX1_116/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4397 DFFNEGX1_116/a_17_6# INVX2_194/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4398 DFFNEGX1_138/a_76_6# INVX2_259/Y DFFNEGX1_138/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M4399 gnd INVX2_259/Y DFFNEGX1_138/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4400 DFFNEGX1_138/a_66_6# DFFNEGX1_138/a_2_6# DFFNEGX1_138/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4401 out_load DFFNEGX1_138/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4402 DFFNEGX1_138/a_23_6# INVX2_259/Y DFFNEGX1_138/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M4403 DFFNEGX1_138/a_23_6# DFFNEGX1_138/a_2_6# DFFNEGX1_138/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M4404 gnd DFFNEGX1_138/a_34_4# DFFNEGX1_138/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4405 vdd DFFNEGX1_138/a_34_4# DFFNEGX1_138/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M4406 DFFNEGX1_138/a_61_74# DFFNEGX1_138/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4407 DFFNEGX1_138/a_34_4# DFFNEGX1_138/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4408 DFFNEGX1_138/a_34_4# DFFNEGX1_138/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4409 vdd out_load DFFNEGX1_138/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4410 gnd out_load DFFNEGX1_138/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4411 DFFNEGX1_138/a_61_6# DFFNEGX1_138/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4412 DFFNEGX1_138/a_76_84# DFFNEGX1_138/a_2_6# DFFNEGX1_138/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M4413 out_load DFFNEGX1_138/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4414 vdd INVX2_259/Y DFFNEGX1_138/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4415 DFFNEGX1_138/a_31_6# DFFNEGX1_138/a_2_6# DFFNEGX1_138/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4416 DFFNEGX1_138/a_66_6# INVX2_259/Y DFFNEGX1_138/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4417 DFFNEGX1_138/a_17_74# NOR2X1_124/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4418 DFFNEGX1_138/a_31_74# INVX2_259/Y DFFNEGX1_138/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4419 DFFNEGX1_138/a_17_6# NOR2X1_124/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4420 DFFNEGX1_127/a_76_6# BUFX2_5/Y DFFNEGX1_127/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M4421 gnd BUFX2_5/Y DFFNEGX1_127/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4422 DFFNEGX1_127/a_66_6# DFFNEGX1_127/a_2_6# DFFNEGX1_127/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4423 out_n_nearby[0] DFFNEGX1_127/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4424 DFFNEGX1_127/a_23_6# BUFX2_5/Y DFFNEGX1_127/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M4425 DFFNEGX1_127/a_23_6# DFFNEGX1_127/a_2_6# DFFNEGX1_127/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M4426 gnd DFFNEGX1_127/a_34_4# DFFNEGX1_127/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4427 vdd DFFNEGX1_127/a_34_4# DFFNEGX1_127/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M4428 DFFNEGX1_127/a_61_74# DFFNEGX1_127/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4429 DFFNEGX1_127/a_34_4# DFFNEGX1_127/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4430 DFFNEGX1_127/a_34_4# DFFNEGX1_127/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4431 vdd out_n_nearby[0] DFFNEGX1_127/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4432 gnd out_n_nearby[0] DFFNEGX1_127/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4433 DFFNEGX1_127/a_61_6# DFFNEGX1_127/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4434 DFFNEGX1_127/a_76_84# DFFNEGX1_127/a_2_6# DFFNEGX1_127/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M4435 out_n_nearby[0] DFFNEGX1_127/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4436 vdd BUFX2_5/Y DFFNEGX1_127/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4437 DFFNEGX1_127/a_31_6# DFFNEGX1_127/a_2_6# DFFNEGX1_127/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4438 DFFNEGX1_127/a_66_6# BUFX2_5/Y DFFNEGX1_127/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4439 DFFNEGX1_127/a_17_74# OAI21X1_60/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4440 DFFNEGX1_127/a_31_74# BUFX2_5/Y DFFNEGX1_127/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4441 DFFNEGX1_127/a_17_6# OAI21X1_60/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4442 gnd OAI21X1_1/A OAI21X1_110/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M4443 vdd NAND2X1_99/Y OAI21X1_110/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M4444 OAI21X1_110/Y NAND2X1_99/Y OAI21X1_110/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4445 OAI21X1_110/Y INVX2_217/Y OAI21X1_110/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4446 OAI21X1_110/a_9_54# OAI21X1_1/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4447 OAI21X1_110/a_2_6# INVX2_217/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4448 gnd INVX2_23/Y OAI21X1_121/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M4449 vdd AOI22X1_70/Y AOI21X1_8/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M4450 AOI21X1_8/B AOI22X1_70/Y OAI21X1_121/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4451 AOI21X1_8/B NOR2X1_110/B OAI21X1_121/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4452 OAI21X1_121/a_9_54# INVX2_23/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4453 OAI21X1_121/a_2_6# NOR2X1_110/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4454 gnd OAI22X1_70/Y OAI21X1_143/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M4455 vdd INVX2_38/Y AOI21X1_16/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M4456 AOI21X1_16/B INVX2_38/Y OAI21X1_143/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4457 AOI21X1_16/B OAI22X1_69/Y OAI21X1_143/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4458 OAI21X1_143/a_9_54# OAI22X1_70/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4459 OAI21X1_143/a_2_6# OAI22X1_69/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4460 gnd out_global_score[25] AOI22X1_8/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M4461 INVX2_191/A INVX2_257/Y AOI22X1_8/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M4462 AOI22X1_8/a_11_6# HAX1_5/YS gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4463 AOI22X1_8/a_2_54# INVX2_257/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M4464 AOI22X1_8/a_28_6# INVX2_255/Y INVX2_191/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4465 vdd HAX1_5/YS AOI22X1_8/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4466 INVX2_191/A INVX2_255/Y AOI22X1_8/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M4467 AOI22X1_8/a_2_54# out_global_score[25] INVX2_191/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4468 gnd OAI22X1_88/Y OAI21X1_154/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M4469 vdd XOR2X1_4/Y OAI21X1_154/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M4470 OAI21X1_154/Y XOR2X1_4/Y OAI21X1_154/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4471 OAI21X1_154/Y OAI22X1_87/Y OAI21X1_154/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4472 OAI21X1_154/a_9_54# OAI22X1_88/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4473 OAI21X1_154/a_2_6# OAI22X1_87/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4474 gnd AOI21X1_14/Y OAI21X1_132/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M4475 vdd XOR2X1_13/Y OAI21X1_132/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M4476 OAI21X1_132/Y XOR2X1_13/Y OAI21X1_132/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4477 OAI21X1_132/Y AOI21X1_13/Y OAI21X1_132/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4478 OAI21X1_132/a_9_54# AOI21X1_14/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4479 OAI21X1_132/a_2_6# AOI21X1_13/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4480 OAI21X1_9/C out_mines[21] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M4481 NAND2X1_18/a_9_6# out_mines[21] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4482 vdd OAI21X1_9/A OAI21X1_9/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4483 OAI21X1_9/C OAI21X1_9/A NAND2X1_18/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4484 OAI21X1_27/C out_mines[12] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M4485 NAND2X1_29/a_9_6# out_mines[12] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4486 vdd INVX2_236/Y OAI21X1_27/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4487 OAI21X1_27/C INVX2_236/Y NAND2X1_29/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4488 gnd out_global_score[17] AOI22X1_16/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M4489 INVX2_199/A INVX2_257/Y AOI22X1_16/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M4490 AOI22X1_16/a_11_6# HAX1_13/YS gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4491 AOI22X1_16/a_2_54# INVX2_257/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M4492 AOI22X1_16/a_28_6# OR2X1_11/B INVX2_199/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4493 vdd HAX1_13/YS AOI22X1_16/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4494 INVX2_199/A OR2X1_11/B AOI22X1_16/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M4495 AOI22X1_16/a_2_54# out_global_score[17] INVX2_199/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4496 gnd out_global_score[6] AOI22X1_27/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M4497 INVX2_210/A INVX2_258/Y AOI22X1_27/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M4498 AOI22X1_27/a_11_6# HAX1_24/YS gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4499 AOI22X1_27/a_2_54# INVX2_258/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M4500 AOI22X1_27/a_28_6# OR2X1_11/B INVX2_210/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4501 vdd HAX1_24/YS AOI22X1_27/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4502 INVX2_210/A OR2X1_11/B AOI22X1_27/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M4503 AOI22X1_27/a_2_54# out_global_score[6] INVX2_210/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4504 gnd out_temp_decoded[19] AOI22X1_38/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M4505 OAI21X1_68/C out_mines[18] AOI22X1_38/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M4506 AOI22X1_38/a_11_6# out_temp_decoded[18] gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4507 AOI22X1_38/a_2_54# out_mines[18] vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M4508 AOI22X1_38/a_28_6# out_mines[19] OAI21X1_68/C Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4509 vdd out_temp_decoded[18] AOI22X1_38/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4510 OAI21X1_68/C out_mines[19] AOI22X1_38/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M4511 AOI22X1_38/a_2_54# out_temp_decoded[19] OAI21X1_68/C vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4512 gnd out_temp_cleared[20] AOI22X1_49/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M4513 NAND3X1_44/A out_mines[19] AOI22X1_49/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M4514 AOI22X1_49/a_11_6# out_temp_cleared[19] gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4515 AOI22X1_49/a_2_54# out_mines[19] vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M4516 AOI22X1_49/a_28_6# out_mines[20] NAND3X1_44/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4517 vdd out_temp_cleared[19] AOI22X1_49/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4518 NAND3X1_44/A out_mines[20] AOI22X1_49/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M4519 AOI22X1_49/a_2_54# out_temp_cleared[20] NAND3X1_44/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4520 vdd HAX1_41/A HAX1_41/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M4521 HAX1_41/a_41_74# HAX1_41/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M4522 HAX1_41/a_9_6# HAX1_41/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4523 HAX1_41/a_41_74# HAX1_41/B HAX1_41/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M4524 vdd HAX1_41/A HAX1_41/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4525 vdd HAX1_41/a_2_74# OR2X1_4/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4526 HAX1_41/a_38_6# HAX1_41/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4527 HAX1_41/YS HAX1_41/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4528 HAX1_41/a_38_6# HAX1_41/A HAX1_41/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4529 HAX1_41/YS HAX1_41/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4530 HAX1_41/a_2_74# HAX1_41/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4531 HAX1_41/a_2_74# HAX1_41/B HAX1_41/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4532 HAX1_41/a_49_54# HAX1_41/B HAX1_41/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4533 gnd HAX1_41/a_2_74# OR2X1_4/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M4534 vdd HAX1_30/A HAX1_30/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M4535 HAX1_30/a_41_74# HAX1_30/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M4536 HAX1_30/a_9_6# HAX1_30/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4537 HAX1_30/a_41_74# HAX1_30/B HAX1_30/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M4538 vdd HAX1_30/A HAX1_30/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4539 vdd HAX1_30/a_2_74# FAX1_10/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4540 HAX1_30/a_38_6# HAX1_30/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4541 FAX1_3/A HAX1_30/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4542 HAX1_30/a_38_6# HAX1_30/A HAX1_30/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4543 FAX1_3/A HAX1_30/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4544 HAX1_30/a_2_74# HAX1_30/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4545 HAX1_30/a_2_74# HAX1_30/B HAX1_30/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4546 HAX1_30/a_49_54# HAX1_30/B HAX1_30/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4547 gnd HAX1_30/a_2_74# FAX1_10/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M4548 gnd OAI21X1_0/A OAI21X1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M4549 vdd OAI21X1_0/C INVX2_52/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M4550 INVX2_52/A OAI21X1_0/C OAI21X1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4551 INVX2_52/A OAI21X1_1/B OAI21X1_0/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4552 OAI21X1_0/a_9_54# OAI21X1_0/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4553 OAI21X1_0/a_2_6# OAI21X1_1/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4554 gnd OR2X1_9/Y XOR2X1_3/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4555 XOR2X1_3/Y XOR2X1_3/a_2_6# XOR2X1_3/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M4556 XOR2X1_3/a_13_43# out_temp_data_in[2] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4557 XOR2X1_3/a_18_54# XOR2X1_3/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4558 XOR2X1_3/a_35_6# OR2X1_9/Y XOR2X1_3/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4559 XOR2X1_3/a_18_6# XOR2X1_3/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4560 vdd OR2X1_9/Y XOR2X1_3/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4561 vdd out_temp_data_in[2] XOR2X1_3/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4562 XOR2X1_3/Y OR2X1_9/Y XOR2X1_3/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M4563 XOR2X1_3/a_35_54# XOR2X1_3/a_2_6# XOR2X1_3/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4564 XOR2X1_3/a_13_43# out_temp_data_in[2] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4565 gnd out_temp_data_in[2] XOR2X1_3/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4566 gnd MUX2X1_4/A MUX2X1_4/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M4567 MUX2X1_4/a_17_50# XOR2X1_8/Y vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4568 MUX2X1_4/Y NOR2X1_7/Y MUX2X1_4/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M4569 MUX2X1_4/a_30_54# MUX2X1_4/a_2_10# MUX2X1_4/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4570 MUX2X1_4/a_17_10# XOR2X1_8/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4571 vdd NOR2X1_7/Y MUX2X1_4/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4572 MUX2X1_4/a_30_10# NOR2X1_7/Y MUX2X1_4/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M4573 gnd NOR2X1_7/Y MUX2X1_4/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M4574 vdd MUX2X1_4/A MUX2X1_4/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4575 MUX2X1_4/Y MUX2X1_4/a_2_10# MUX2X1_4/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4576 INVX2_121/Y INVX2_121/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4577 INVX2_121/Y INVX2_121/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4578 INVX2_132/Y out_alu gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4579 INVX2_132/Y out_alu vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4580 OAI22X1_2/D out_temp_cleared[3] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4581 OAI22X1_2/D out_temp_cleared[3] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4582 MUX2X1_22/B XNOR2X1_5/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4583 MUX2X1_22/B XNOR2X1_5/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4584 MUX2X1_14/A FAX1_0/YS gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4585 MUX2X1_14/A FAX1_0/YS vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4586 NOR2X1_4/A MUX2X1_9/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4587 NOR2X1_4/A MUX2X1_9/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4588 INVX2_198/Y INVX2_198/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4589 INVX2_198/Y INVX2_198/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4590 HAX1_48/A MUX2X1_27/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4591 HAX1_48/A MUX2X1_27/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4592 INVX2_187/Y INVX2_187/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4593 INVX2_187/Y INVX2_187/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4594 DFFNEGX1_16/a_76_6# BUFX2_16/Y DFFNEGX1_16/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M4595 gnd BUFX2_16/Y DFFNEGX1_16/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4596 DFFNEGX1_16/a_66_6# DFFNEGX1_16/a_2_6# DFFNEGX1_16/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4597 out_mines[9] DFFNEGX1_16/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4598 DFFNEGX1_16/a_23_6# BUFX2_16/Y DFFNEGX1_16/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M4599 DFFNEGX1_16/a_23_6# DFFNEGX1_16/a_2_6# DFFNEGX1_16/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M4600 gnd DFFNEGX1_16/a_34_4# DFFNEGX1_16/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4601 vdd DFFNEGX1_16/a_34_4# DFFNEGX1_16/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M4602 DFFNEGX1_16/a_61_74# DFFNEGX1_16/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4603 DFFNEGX1_16/a_34_4# DFFNEGX1_16/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4604 DFFNEGX1_16/a_34_4# DFFNEGX1_16/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4605 vdd out_mines[9] DFFNEGX1_16/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4606 gnd out_mines[9] DFFNEGX1_16/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4607 DFFNEGX1_16/a_61_6# DFFNEGX1_16/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4608 DFFNEGX1_16/a_76_84# DFFNEGX1_16/a_2_6# DFFNEGX1_16/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M4609 out_mines[9] DFFNEGX1_16/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4610 vdd BUFX2_16/Y DFFNEGX1_16/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4611 DFFNEGX1_16/a_31_6# DFFNEGX1_16/a_2_6# DFFNEGX1_16/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4612 DFFNEGX1_16/a_66_6# BUFX2_16/Y DFFNEGX1_16/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4613 DFFNEGX1_16/a_17_74# OAI21X1_33/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4614 DFFNEGX1_16/a_31_74# BUFX2_16/Y DFFNEGX1_16/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4615 DFFNEGX1_16/a_17_6# OAI21X1_33/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4616 DFFNEGX1_27/a_76_6# BUFX2_15/Y DFFNEGX1_27/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M4617 gnd BUFX2_15/Y DFFNEGX1_27/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4618 DFFNEGX1_27/a_66_6# DFFNEGX1_27/a_2_6# DFFNEGX1_27/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4619 out_mines[11] DFFNEGX1_27/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4620 DFFNEGX1_27/a_23_6# BUFX2_15/Y DFFNEGX1_27/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M4621 DFFNEGX1_27/a_23_6# DFFNEGX1_27/a_2_6# DFFNEGX1_27/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M4622 gnd DFFNEGX1_27/a_34_4# DFFNEGX1_27/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4623 vdd DFFNEGX1_27/a_34_4# DFFNEGX1_27/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M4624 DFFNEGX1_27/a_61_74# DFFNEGX1_27/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4625 DFFNEGX1_27/a_34_4# DFFNEGX1_27/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4626 DFFNEGX1_27/a_34_4# DFFNEGX1_27/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4627 vdd out_mines[11] DFFNEGX1_27/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4628 gnd out_mines[11] DFFNEGX1_27/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4629 DFFNEGX1_27/a_61_6# DFFNEGX1_27/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4630 DFFNEGX1_27/a_76_84# DFFNEGX1_27/a_2_6# DFFNEGX1_27/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M4631 out_mines[11] DFFNEGX1_27/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4632 vdd BUFX2_15/Y DFFNEGX1_27/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4633 DFFNEGX1_27/a_31_6# DFFNEGX1_27/a_2_6# DFFNEGX1_27/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4634 DFFNEGX1_27/a_66_6# BUFX2_15/Y DFFNEGX1_27/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4635 DFFNEGX1_27/a_17_74# OAI21X1_29/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4636 DFFNEGX1_27/a_31_74# BUFX2_15/Y DFFNEGX1_27/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4637 DFFNEGX1_27/a_17_6# OAI21X1_29/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4638 DFFNEGX1_49/a_76_6# BUFX2_14/Y DFFNEGX1_49/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M4639 gnd BUFX2_14/Y DFFNEGX1_49/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4640 DFFNEGX1_49/a_66_6# DFFNEGX1_49/a_2_6# DFFNEGX1_49/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4641 out_temp_decoded[17] DFFNEGX1_49/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4642 DFFNEGX1_49/a_23_6# BUFX2_14/Y DFFNEGX1_49/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M4643 DFFNEGX1_49/a_23_6# DFFNEGX1_49/a_2_6# DFFNEGX1_49/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M4644 gnd DFFNEGX1_49/a_34_4# DFFNEGX1_49/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4645 vdd DFFNEGX1_49/a_34_4# DFFNEGX1_49/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M4646 DFFNEGX1_49/a_61_74# DFFNEGX1_49/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4647 DFFNEGX1_49/a_34_4# DFFNEGX1_49/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4648 DFFNEGX1_49/a_34_4# DFFNEGX1_49/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4649 vdd out_temp_decoded[17] DFFNEGX1_49/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4650 gnd out_temp_decoded[17] DFFNEGX1_49/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4651 DFFNEGX1_49/a_61_6# DFFNEGX1_49/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4652 DFFNEGX1_49/a_76_84# DFFNEGX1_49/a_2_6# DFFNEGX1_49/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M4653 out_temp_decoded[17] DFFNEGX1_49/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4654 vdd BUFX2_14/Y DFFNEGX1_49/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4655 DFFNEGX1_49/a_31_6# DFFNEGX1_49/a_2_6# DFFNEGX1_49/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4656 DFFNEGX1_49/a_66_6# BUFX2_14/Y DFFNEGX1_49/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4657 DFFNEGX1_49/a_17_74# OAI21X1_99/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4658 DFFNEGX1_49/a_31_74# BUFX2_14/Y DFFNEGX1_49/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4659 DFFNEGX1_49/a_17_6# OAI21X1_99/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4660 DFFNEGX1_38/a_76_6# BUFX2_15/Y DFFNEGX1_38/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M4661 gnd BUFX2_15/Y DFFNEGX1_38/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4662 DFFNEGX1_38/a_66_6# DFFNEGX1_38/a_2_6# DFFNEGX1_38/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4663 out_temp_data_in[3] DFFNEGX1_38/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4664 DFFNEGX1_38/a_23_6# BUFX2_15/Y DFFNEGX1_38/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M4665 DFFNEGX1_38/a_23_6# DFFNEGX1_38/a_2_6# DFFNEGX1_38/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M4666 gnd DFFNEGX1_38/a_34_4# DFFNEGX1_38/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4667 vdd DFFNEGX1_38/a_34_4# DFFNEGX1_38/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M4668 DFFNEGX1_38/a_61_74# DFFNEGX1_38/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4669 DFFNEGX1_38/a_34_4# DFFNEGX1_38/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4670 DFFNEGX1_38/a_34_4# DFFNEGX1_38/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4671 vdd out_temp_data_in[3] DFFNEGX1_38/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4672 gnd out_temp_data_in[3] DFFNEGX1_38/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4673 DFFNEGX1_38/a_61_6# DFFNEGX1_38/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4674 DFFNEGX1_38/a_76_84# DFFNEGX1_38/a_2_6# DFFNEGX1_38/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M4675 out_temp_data_in[3] DFFNEGX1_38/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4676 vdd BUFX2_15/Y DFFNEGX1_38/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4677 DFFNEGX1_38/a_31_6# DFFNEGX1_38/a_2_6# DFFNEGX1_38/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4678 DFFNEGX1_38/a_66_6# BUFX2_15/Y DFFNEGX1_38/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4679 DFFNEGX1_38/a_17_74# OAI21X1_110/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4680 DFFNEGX1_38/a_31_74# BUFX2_15/Y DFFNEGX1_38/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4681 DFFNEGX1_38/a_17_6# OAI21X1_110/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4682 gnd out_temp_mine_cnt[2] XOR2X1_14/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4683 XOR2X1_14/Y XOR2X1_14/a_2_6# XOR2X1_14/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M4684 XOR2X1_14/a_13_43# in_n_mines[2] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4685 XOR2X1_14/a_18_54# XOR2X1_14/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4686 XOR2X1_14/a_35_6# out_temp_mine_cnt[2] XOR2X1_14/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4687 XOR2X1_14/a_18_6# XOR2X1_14/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4688 vdd out_temp_mine_cnt[2] XOR2X1_14/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4689 vdd in_n_mines[2] XOR2X1_14/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4690 XOR2X1_14/Y out_temp_mine_cnt[2] XOR2X1_14/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M4691 XOR2X1_14/a_35_54# XOR2X1_14/a_2_6# XOR2X1_14/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4692 XOR2X1_14/a_13_43# in_n_mines[2] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4693 gnd in_n_mines[2] XOR2X1_14/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4694 gnd XOR2X1_26/Y XOR2X1_25/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4695 XOR2X1_25/Y XOR2X1_25/a_2_6# XOR2X1_25/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M4696 XOR2X1_25/a_13_43# XOR2X1_25/B gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4697 XOR2X1_25/a_18_54# XOR2X1_25/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4698 XOR2X1_25/a_35_6# XOR2X1_26/Y XOR2X1_25/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4699 XOR2X1_25/a_18_6# XOR2X1_25/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4700 vdd XOR2X1_26/Y XOR2X1_25/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4701 vdd XOR2X1_25/B XOR2X1_25/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4702 XOR2X1_25/Y XOR2X1_26/Y XOR2X1_25/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M4703 XOR2X1_25/a_35_54# XOR2X1_25/a_2_6# XOR2X1_25/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4704 XOR2X1_25/a_13_43# XOR2X1_25/B vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4705 gnd XOR2X1_25/B XOR2X1_25/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4706 NOR2X1_58/A OAI21X1_1/B vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M4707 NAND3X1_4/a_9_6# OAI21X1_1/B gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M4708 NOR2X1_58/A out_temp_data_in[3] vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4709 NOR2X1_58/A out_temp_data_in[3] NAND3X1_4/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M4710 vdd INVX2_30/Y NOR2X1_58/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4711 NAND3X1_4/a_14_6# INVX2_30/Y NAND3X1_4/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M4712 DFFNEGX1_106/a_76_6# BUFX2_9/Y DFFNEGX1_106/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M4713 gnd BUFX2_9/Y DFFNEGX1_106/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4714 DFFNEGX1_106/a_66_6# DFFNEGX1_106/a_2_6# DFFNEGX1_106/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4715 out_global_score[12] DFFNEGX1_106/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4716 DFFNEGX1_106/a_23_6# BUFX2_9/Y DFFNEGX1_106/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M4717 DFFNEGX1_106/a_23_6# DFFNEGX1_106/a_2_6# DFFNEGX1_106/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M4718 gnd DFFNEGX1_106/a_34_4# DFFNEGX1_106/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4719 vdd DFFNEGX1_106/a_34_4# DFFNEGX1_106/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M4720 DFFNEGX1_106/a_61_74# DFFNEGX1_106/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4721 DFFNEGX1_106/a_34_4# DFFNEGX1_106/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4722 DFFNEGX1_106/a_34_4# DFFNEGX1_106/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4723 vdd out_global_score[12] DFFNEGX1_106/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4724 gnd out_global_score[12] DFFNEGX1_106/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4725 DFFNEGX1_106/a_61_6# DFFNEGX1_106/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4726 DFFNEGX1_106/a_76_84# DFFNEGX1_106/a_2_6# DFFNEGX1_106/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M4727 out_global_score[12] DFFNEGX1_106/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4728 vdd BUFX2_9/Y DFFNEGX1_106/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4729 DFFNEGX1_106/a_31_6# DFFNEGX1_106/a_2_6# DFFNEGX1_106/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4730 DFFNEGX1_106/a_66_6# BUFX2_9/Y DFFNEGX1_106/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4731 DFFNEGX1_106/a_17_74# INVX2_204/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4732 DFFNEGX1_106/a_31_74# BUFX2_9/Y DFFNEGX1_106/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4733 DFFNEGX1_106/a_17_6# INVX2_204/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4734 DFFNEGX1_117/a_76_6# BUFX2_9/Y DFFNEGX1_117/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M4735 gnd BUFX2_9/Y DFFNEGX1_117/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4736 DFFNEGX1_117/a_66_6# DFFNEGX1_117/a_2_6# DFFNEGX1_117/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4737 out_global_score[23] DFFNEGX1_117/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4738 DFFNEGX1_117/a_23_6# BUFX2_9/Y DFFNEGX1_117/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M4739 DFFNEGX1_117/a_23_6# DFFNEGX1_117/a_2_6# DFFNEGX1_117/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M4740 gnd DFFNEGX1_117/a_34_4# DFFNEGX1_117/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4741 vdd DFFNEGX1_117/a_34_4# DFFNEGX1_117/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M4742 DFFNEGX1_117/a_61_74# DFFNEGX1_117/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4743 DFFNEGX1_117/a_34_4# DFFNEGX1_117/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4744 DFFNEGX1_117/a_34_4# DFFNEGX1_117/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4745 vdd out_global_score[23] DFFNEGX1_117/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4746 gnd out_global_score[23] DFFNEGX1_117/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4747 DFFNEGX1_117/a_61_6# DFFNEGX1_117/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4748 DFFNEGX1_117/a_76_84# DFFNEGX1_117/a_2_6# DFFNEGX1_117/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M4749 out_global_score[23] DFFNEGX1_117/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4750 vdd BUFX2_9/Y DFFNEGX1_117/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4751 DFFNEGX1_117/a_31_6# DFFNEGX1_117/a_2_6# DFFNEGX1_117/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4752 DFFNEGX1_117/a_66_6# BUFX2_9/Y DFFNEGX1_117/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4753 DFFNEGX1_117/a_17_74# INVX2_193/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4754 DFFNEGX1_117/a_31_74# BUFX2_9/Y DFFNEGX1_117/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4755 DFFNEGX1_117/a_17_6# INVX2_193/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4756 DFFNEGX1_139/a_76_6# INVX2_259/Y DFFNEGX1_139/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M4757 gnd INVX2_259/Y DFFNEGX1_139/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4758 DFFNEGX1_139/a_66_6# DFFNEGX1_139/a_2_6# DFFNEGX1_139/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4759 out_start DFFNEGX1_139/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4760 DFFNEGX1_139/a_23_6# INVX2_259/Y DFFNEGX1_139/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M4761 DFFNEGX1_139/a_23_6# DFFNEGX1_139/a_2_6# DFFNEGX1_139/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M4762 gnd DFFNEGX1_139/a_34_4# DFFNEGX1_139/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4763 vdd DFFNEGX1_139/a_34_4# DFFNEGX1_139/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M4764 DFFNEGX1_139/a_61_74# DFFNEGX1_139/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4765 DFFNEGX1_139/a_34_4# DFFNEGX1_139/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4766 DFFNEGX1_139/a_34_4# DFFNEGX1_139/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4767 vdd out_start DFFNEGX1_139/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4768 gnd out_start DFFNEGX1_139/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4769 DFFNEGX1_139/a_61_6# DFFNEGX1_139/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4770 DFFNEGX1_139/a_76_84# DFFNEGX1_139/a_2_6# DFFNEGX1_139/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M4771 out_start DFFNEGX1_139/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4772 vdd INVX2_259/Y DFFNEGX1_139/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4773 DFFNEGX1_139/a_31_6# DFFNEGX1_139/a_2_6# DFFNEGX1_139/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4774 DFFNEGX1_139/a_66_6# INVX2_259/Y DFFNEGX1_139/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4775 DFFNEGX1_139/a_17_74# OAI21X1_159/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4776 DFFNEGX1_139/a_31_74# INVX2_259/Y DFFNEGX1_139/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4777 DFFNEGX1_139/a_17_6# OAI21X1_159/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4778 DFFNEGX1_128/a_76_6# INVX2_259/Y DFFNEGX1_128/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M4779 gnd INVX2_259/Y DFFNEGX1_128/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4780 DFFNEGX1_128/a_66_6# DFFNEGX1_128/a_2_6# DFFNEGX1_128/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4781 out_display_done DFFNEGX1_128/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4782 DFFNEGX1_128/a_23_6# INVX2_259/Y DFFNEGX1_128/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M4783 DFFNEGX1_128/a_23_6# DFFNEGX1_128/a_2_6# DFFNEGX1_128/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M4784 gnd DFFNEGX1_128/a_34_4# DFFNEGX1_128/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4785 vdd DFFNEGX1_128/a_34_4# DFFNEGX1_128/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M4786 DFFNEGX1_128/a_61_74# DFFNEGX1_128/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4787 DFFNEGX1_128/a_34_4# DFFNEGX1_128/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4788 DFFNEGX1_128/a_34_4# DFFNEGX1_128/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4789 vdd out_display_done DFFNEGX1_128/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4790 gnd out_display_done DFFNEGX1_128/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4791 DFFNEGX1_128/a_61_6# DFFNEGX1_128/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4792 DFFNEGX1_128/a_76_84# DFFNEGX1_128/a_2_6# DFFNEGX1_128/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M4793 out_display_done DFFNEGX1_128/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4794 vdd INVX2_259/Y DFFNEGX1_128/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4795 DFFNEGX1_128/a_31_6# DFFNEGX1_128/a_2_6# DFFNEGX1_128/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4796 DFFNEGX1_128/a_66_6# INVX2_259/Y DFFNEGX1_128/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4797 DFFNEGX1_128/a_17_74# OAI21X1_59/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4798 DFFNEGX1_128/a_31_74# INVX2_259/Y DFFNEGX1_128/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4799 DFFNEGX1_128/a_17_6# OAI21X1_59/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4800 gnd INVX2_63/Y OAI21X1_100/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M4801 vdd NAND2X1_87/Y OAI21X1_100/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M4802 OAI21X1_100/Y NAND2X1_87/Y OAI21X1_100/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4803 OAI21X1_100/Y BUFX2_23/Y OAI21X1_100/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4804 OAI21X1_100/a_9_54# INVX2_63/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4805 OAI21X1_100/a_2_6# BUFX2_23/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4806 gnd INVX2_18/Y OAI21X1_122/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M4807 vdd AOI22X1_71/Y AOI22X1_69/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M4808 AOI22X1_69/B AOI22X1_71/Y OAI21X1_122/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4809 AOI22X1_69/B NOR2X1_110/B OAI21X1_122/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4810 OAI21X1_122/a_9_54# INVX2_18/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4811 OAI21X1_122/a_2_6# NOR2X1_110/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4812 gnd INVX2_30/Y OAI21X1_111/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M4813 vdd OAI21X1_111/C OAI21X1_111/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M4814 OAI21X1_111/Y OAI21X1_111/C OAI21X1_111/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4815 OAI21X1_111/Y INVX2_217/Y OAI21X1_111/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4816 OAI21X1_111/a_9_54# INVX2_30/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4817 OAI21X1_111/a_2_6# INVX2_217/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4818 gnd out_global_score[24] AOI22X1_9/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M4819 INVX2_192/A INVX2_257/Y AOI22X1_9/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M4820 AOI22X1_9/a_11_6# HAX1_6/YS gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4821 AOI22X1_9/a_2_54# INVX2_257/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M4822 AOI22X1_9/a_28_6# INVX2_255/Y INVX2_192/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4823 vdd HAX1_6/YS AOI22X1_9/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4824 INVX2_192/A INVX2_255/Y AOI22X1_9/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M4825 AOI22X1_9/a_2_54# out_global_score[24] INVX2_192/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4826 gnd OAI22X1_72/Y OAI21X1_144/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M4827 vdd XOR2X1_3/Y AOI21X1_16/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M4828 AOI21X1_16/A XOR2X1_3/Y OAI21X1_144/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4829 AOI21X1_16/A OAI22X1_71/Y OAI21X1_144/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4830 OAI21X1_144/a_9_54# OAI22X1_72/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4831 OAI21X1_144/a_2_6# OAI22X1_71/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4832 gnd INVX2_117/Y OAI21X1_155/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M4833 vdd NAND3X1_49/Y OAI21X1_155/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M4834 OAI21X1_155/Y NAND3X1_49/Y OAI21X1_155/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4835 OAI21X1_155/Y OAI21X1_156/Y OAI21X1_155/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4836 OAI21X1_155/a_9_54# INVX2_117/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4837 OAI21X1_155/a_2_6# OAI21X1_156/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4838 gnd OAI22X1_54/Y OAI21X1_133/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M4839 vdd out_temp_data_in[2] AOI21X1_13/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M4840 AOI21X1_13/B out_temp_data_in[2] OAI21X1_133/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4841 AOI21X1_13/B OAI22X1_53/Y OAI21X1_133/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4842 OAI21X1_133/a_9_54# OAI22X1_54/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4843 OAI21X1_133/a_2_6# OAI22X1_53/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4844 OAI21X1_11/C out_mines[20] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M4845 NAND2X1_19/a_9_6# out_mines[20] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4846 vdd INVX2_234/Y OAI21X1_11/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4847 OAI21X1_11/C INVX2_234/Y NAND2X1_19/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4848 gnd out_global_score[16] AOI22X1_17/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M4849 INVX2_200/A INVX2_257/Y AOI22X1_17/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M4850 AOI22X1_17/a_11_6# HAX1_14/YS gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4851 AOI22X1_17/a_2_54# INVX2_257/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M4852 AOI22X1_17/a_28_6# OR2X1_11/B INVX2_200/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4853 vdd HAX1_14/YS AOI22X1_17/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4854 INVX2_200/A OR2X1_11/B AOI22X1_17/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M4855 AOI22X1_17/a_2_54# out_global_score[16] INVX2_200/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4856 gnd out_global_score[5] AOI22X1_28/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M4857 INVX2_211/A INVX2_258/Y AOI22X1_28/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M4858 AOI22X1_28/a_11_6# HAX1_25/YS gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4859 AOI22X1_28/a_2_54# INVX2_258/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M4860 AOI22X1_28/a_28_6# INVX2_255/Y INVX2_211/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4861 vdd HAX1_25/YS AOI22X1_28/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4862 INVX2_211/A INVX2_255/Y AOI22X1_28/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M4863 AOI22X1_28/a_2_54# out_global_score[5] INVX2_211/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4864 gnd out_temp_decoded[16] AOI22X1_39/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M4865 OAI21X1_69/C out_mines[15] AOI22X1_39/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M4866 AOI22X1_39/a_11_6# out_temp_decoded[15] gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4867 AOI22X1_39/a_2_54# out_mines[15] vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M4868 AOI22X1_39/a_28_6# out_mines[16] OAI21X1_69/C Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4869 vdd out_temp_decoded[15] AOI22X1_39/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4870 OAI21X1_69/C out_mines[16] AOI22X1_39/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M4871 AOI22X1_39/a_2_54# out_temp_decoded[16] OAI21X1_69/C vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4872 vdd out_global_score[10] HAX1_20/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M4873 HAX1_20/a_41_74# HAX1_20/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M4874 HAX1_20/a_9_6# out_global_score[10] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4875 HAX1_20/a_41_74# HAX1_20/B HAX1_20/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M4876 vdd out_global_score[10] HAX1_20/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4877 vdd HAX1_20/a_2_74# HAX1_19/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4878 HAX1_20/a_38_6# HAX1_20/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4879 HAX1_20/YS HAX1_20/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4880 HAX1_20/a_38_6# out_global_score[10] HAX1_20/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4881 HAX1_20/YS HAX1_20/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4882 HAX1_20/a_2_74# HAX1_20/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4883 HAX1_20/a_2_74# HAX1_20/B HAX1_20/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4884 HAX1_20/a_49_54# HAX1_20/B HAX1_20/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4885 gnd HAX1_20/a_2_74# HAX1_19/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M4886 vdd HAX1_42/A HAX1_42/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M4887 HAX1_42/a_41_74# HAX1_42/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M4888 HAX1_42/a_9_6# HAX1_42/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4889 HAX1_42/a_41_74# HAX1_42/B HAX1_42/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M4890 vdd HAX1_42/A HAX1_42/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4891 vdd HAX1_42/a_2_74# HAX1_43/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4892 HAX1_42/a_38_6# HAX1_42/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4893 HAX1_42/YS HAX1_42/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4894 HAX1_42/a_38_6# HAX1_42/A HAX1_42/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4895 HAX1_42/YS HAX1_42/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4896 HAX1_42/a_2_74# HAX1_42/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4897 HAX1_42/a_2_74# HAX1_42/B HAX1_42/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4898 HAX1_42/a_49_54# HAX1_42/B HAX1_42/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4899 gnd HAX1_42/a_2_74# HAX1_43/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M4900 vdd HAX1_31/A HAX1_31/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M4901 HAX1_31/a_41_74# HAX1_31/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M4902 HAX1_31/a_9_6# HAX1_31/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4903 HAX1_31/a_41_74# HAX1_31/B HAX1_31/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M4904 vdd HAX1_31/A HAX1_31/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4905 vdd HAX1_31/a_2_74# FAX1_12/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4906 HAX1_31/a_38_6# HAX1_31/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4907 FAX1_14/A HAX1_31/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4908 HAX1_31/a_38_6# HAX1_31/A HAX1_31/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4909 FAX1_14/A HAX1_31/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4910 HAX1_31/a_2_74# HAX1_31/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4911 HAX1_31/a_2_74# HAX1_31/B HAX1_31/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4912 HAX1_31/a_49_54# HAX1_31/B HAX1_31/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4913 gnd HAX1_31/a_2_74# FAX1_12/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M4914 gnd OAI21X1_1/A OAI21X1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M4915 vdd OAI21X1_2/Y AND2X2_6/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M4916 AND2X2_6/B OAI21X1_2/Y OAI21X1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4917 AND2X2_6/B OAI21X1_1/B OAI21X1_1/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4918 OAI21X1_1/a_9_54# OAI21X1_1/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4919 OAI21X1_1/a_2_6# OAI21X1_1/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4920 gnd out_mines[5] OAI22X1_80/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M4921 OAI22X1_80/a_2_6# out_mines[4] OAI22X1_80/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M4922 OAI22X1_80/Y OAI22X1_88/D OAI22X1_80/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4923 OAI22X1_80/Y OAI22X1_88/B OAI22X1_80/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M4924 OAI22X1_80/a_28_54# OAI22X1_88/D OAI22X1_80/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4925 OAI22X1_80/a_9_54# out_mines[5] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4926 OAI22X1_80/a_2_6# OAI22X1_88/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4927 vdd out_mines[4] OAI22X1_80/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4928 gnd out_temp_data_in[1] XOR2X1_4/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4929 XOR2X1_4/Y XOR2X1_4/a_2_6# XOR2X1_4/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M4930 XOR2X1_4/a_13_43# out_temp_data_in[2] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4931 XOR2X1_4/a_18_54# XOR2X1_4/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4932 XOR2X1_4/a_35_6# out_temp_data_in[1] XOR2X1_4/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4933 XOR2X1_4/a_18_6# XOR2X1_4/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4934 vdd out_temp_data_in[1] XOR2X1_4/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4935 vdd out_temp_data_in[2] XOR2X1_4/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M4936 XOR2X1_4/Y out_temp_data_in[1] XOR2X1_4/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M4937 XOR2X1_4/a_35_54# XOR2X1_4/a_2_6# XOR2X1_4/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4938 XOR2X1_4/a_13_43# out_temp_data_in[2] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4939 gnd out_temp_data_in[2] XOR2X1_4/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4940 gnd MUX2X1_5/A MUX2X1_5/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M4941 MUX2X1_5/a_17_50# HAX1_39/A vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4942 MUX2X1_5/Y OR2X1_5/Y MUX2X1_5/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M4943 MUX2X1_5/a_30_54# MUX2X1_5/a_2_10# MUX2X1_5/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M4944 MUX2X1_5/a_17_10# HAX1_39/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4945 vdd OR2X1_5/Y MUX2X1_5/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4946 MUX2X1_5/a_30_10# OR2X1_5/Y MUX2X1_5/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M4947 gnd OR2X1_5/Y MUX2X1_5/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M4948 vdd MUX2X1_5/A MUX2X1_5/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M4949 MUX2X1_5/Y MUX2X1_5/a_2_10# MUX2X1_5/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4950 INVX2_100/Y out_temp_cleared[13] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4951 INVX2_100/Y out_temp_cleared[13] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4952 INVX2_111/Y out_temp_cleared[2] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4953 INVX2_111/Y out_temp_cleared[2] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4954 INVX2_122/Y INVX2_122/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4955 INVX2_122/Y INVX2_122/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4956 NOR2X1_2/A MUX2X1_19/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4957 NOR2X1_2/A MUX2X1_19/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4958 HAX1_40/A MUX2X1_7/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4959 HAX1_40/A MUX2X1_7/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4960 MUX2X1_9/A XOR2X1_9/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4961 MUX2X1_9/A XOR2X1_9/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4962 INVX2_133/Y INVX2_133/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4963 INVX2_133/Y INVX2_133/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4964 INVX2_199/Y INVX2_199/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4965 INVX2_199/Y INVX2_199/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4966 NOR2X1_64/B OAI21X1_4/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4967 NOR2X1_64/B OAI21X1_4/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4968 INVX2_188/Y INVX2_188/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4969 INVX2_188/Y INVX2_188/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4970 DFFNEGX1_17/a_76_6# BUFX2_16/Y DFFNEGX1_17/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M4971 gnd BUFX2_16/Y DFFNEGX1_17/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4972 DFFNEGX1_17/a_66_6# DFFNEGX1_17/a_2_6# DFFNEGX1_17/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4973 out_temp_index[4] DFFNEGX1_17/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4974 DFFNEGX1_17/a_23_6# BUFX2_16/Y DFFNEGX1_17/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M4975 DFFNEGX1_17/a_23_6# DFFNEGX1_17/a_2_6# DFFNEGX1_17/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M4976 gnd DFFNEGX1_17/a_34_4# DFFNEGX1_17/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4977 vdd DFFNEGX1_17/a_34_4# DFFNEGX1_17/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M4978 DFFNEGX1_17/a_61_74# DFFNEGX1_17/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M4979 DFFNEGX1_17/a_34_4# DFFNEGX1_17/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4980 DFFNEGX1_17/a_34_4# DFFNEGX1_17/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M4981 vdd out_temp_index[4] DFFNEGX1_17/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4982 gnd out_temp_index[4] DFFNEGX1_17/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4983 DFFNEGX1_17/a_61_6# DFFNEGX1_17/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4984 DFFNEGX1_17/a_76_84# DFFNEGX1_17/a_2_6# DFFNEGX1_17/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M4985 out_temp_index[4] DFFNEGX1_17/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M4986 vdd BUFX2_16/Y DFFNEGX1_17/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M4987 DFFNEGX1_17/a_31_6# DFFNEGX1_17/a_2_6# DFFNEGX1_17/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4988 DFFNEGX1_17/a_66_6# BUFX2_16/Y DFFNEGX1_17/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4989 DFFNEGX1_17/a_17_74# OAI21X1_53/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4990 DFFNEGX1_17/a_31_74# BUFX2_16/Y DFFNEGX1_17/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M4991 DFFNEGX1_17/a_17_6# OAI21X1_53/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M4992 DFFNEGX1_28/a_76_6# BUFX2_15/Y DFFNEGX1_28/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M4993 gnd BUFX2_15/Y DFFNEGX1_28/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M4994 DFFNEGX1_28/a_66_6# DFFNEGX1_28/a_2_6# DFFNEGX1_28/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4995 out_mines[10] DFFNEGX1_28/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M4996 DFFNEGX1_28/a_23_6# BUFX2_15/Y DFFNEGX1_28/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M4997 DFFNEGX1_28/a_23_6# DFFNEGX1_28/a_2_6# DFFNEGX1_28/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M4998 gnd DFFNEGX1_28/a_34_4# DFFNEGX1_28/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M4999 vdd DFFNEGX1_28/a_34_4# DFFNEGX1_28/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M5000 DFFNEGX1_28/a_61_74# DFFNEGX1_28/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5001 DFFNEGX1_28/a_34_4# DFFNEGX1_28/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5002 DFFNEGX1_28/a_34_4# DFFNEGX1_28/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M5003 vdd out_mines[10] DFFNEGX1_28/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5004 gnd out_mines[10] DFFNEGX1_28/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5005 DFFNEGX1_28/a_61_6# DFFNEGX1_28/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5006 DFFNEGX1_28/a_76_84# DFFNEGX1_28/a_2_6# DFFNEGX1_28/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M5007 out_mines[10] DFFNEGX1_28/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5008 vdd BUFX2_15/Y DFFNEGX1_28/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M5009 DFFNEGX1_28/a_31_6# DFFNEGX1_28/a_2_6# DFFNEGX1_28/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5010 DFFNEGX1_28/a_66_6# BUFX2_15/Y DFFNEGX1_28/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5011 DFFNEGX1_28/a_17_74# OAI21X1_31/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5012 DFFNEGX1_28/a_31_74# BUFX2_15/Y DFFNEGX1_28/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5013 DFFNEGX1_28/a_17_6# OAI21X1_31/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5014 DFFNEGX1_39/a_76_6# BUFX2_15/Y DFFNEGX1_39/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M5015 gnd BUFX2_15/Y DFFNEGX1_39/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5016 DFFNEGX1_39/a_66_6# DFFNEGX1_39/a_2_6# DFFNEGX1_39/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5017 out_temp_data_in[2] DFFNEGX1_39/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5018 DFFNEGX1_39/a_23_6# BUFX2_15/Y DFFNEGX1_39/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M5019 DFFNEGX1_39/a_23_6# DFFNEGX1_39/a_2_6# DFFNEGX1_39/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M5020 gnd DFFNEGX1_39/a_34_4# DFFNEGX1_39/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5021 vdd DFFNEGX1_39/a_34_4# DFFNEGX1_39/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M5022 DFFNEGX1_39/a_61_74# DFFNEGX1_39/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5023 DFFNEGX1_39/a_34_4# DFFNEGX1_39/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5024 DFFNEGX1_39/a_34_4# DFFNEGX1_39/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M5025 vdd out_temp_data_in[2] DFFNEGX1_39/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5026 gnd out_temp_data_in[2] DFFNEGX1_39/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5027 DFFNEGX1_39/a_61_6# DFFNEGX1_39/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5028 DFFNEGX1_39/a_76_84# DFFNEGX1_39/a_2_6# DFFNEGX1_39/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M5029 out_temp_data_in[2] DFFNEGX1_39/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5030 vdd BUFX2_15/Y DFFNEGX1_39/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M5031 DFFNEGX1_39/a_31_6# DFFNEGX1_39/a_2_6# DFFNEGX1_39/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5032 DFFNEGX1_39/a_66_6# BUFX2_15/Y DFFNEGX1_39/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5033 DFFNEGX1_39/a_17_74# OAI21X1_109/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5034 DFFNEGX1_39/a_31_74# BUFX2_15/Y DFFNEGX1_39/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5035 DFFNEGX1_39/a_17_6# OAI21X1_109/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5036 gnd out_temp_mine_cnt[4] XOR2X1_15/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5037 XOR2X1_15/Y XOR2X1_15/a_2_6# XOR2X1_15/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M5038 XOR2X1_15/a_13_43# in_n_mines[4] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5039 XOR2X1_15/a_18_54# XOR2X1_15/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M5040 XOR2X1_15/a_35_6# out_temp_mine_cnt[4] XOR2X1_15/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5041 XOR2X1_15/a_18_6# XOR2X1_15/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5042 vdd out_temp_mine_cnt[4] XOR2X1_15/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M5043 vdd in_n_mines[4] XOR2X1_15/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5044 XOR2X1_15/Y out_temp_mine_cnt[4] XOR2X1_15/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M5045 XOR2X1_15/a_35_54# XOR2X1_15/a_2_6# XOR2X1_15/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5046 XOR2X1_15/a_13_43# in_n_mines[4] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5047 gnd in_n_mines[4] XOR2X1_15/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5048 gnd INVX2_45/A XOR2X1_26/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5049 XOR2X1_26/Y XOR2X1_26/a_2_6# XOR2X1_26/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M5050 XOR2X1_26/a_13_43# INVX2_50/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5051 XOR2X1_26/a_18_54# XOR2X1_26/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M5052 XOR2X1_26/a_35_6# INVX2_45/A XOR2X1_26/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5053 XOR2X1_26/a_18_6# XOR2X1_26/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5054 vdd INVX2_45/A XOR2X1_26/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M5055 vdd INVX2_50/Y XOR2X1_26/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5056 XOR2X1_26/Y INVX2_45/A XOR2X1_26/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M5057 XOR2X1_26/a_35_54# XOR2X1_26/a_2_6# XOR2X1_26/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5058 XOR2X1_26/a_13_43# INVX2_50/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5059 gnd INVX2_50/Y XOR2X1_26/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5060 NOR2X1_59/B OAI21X1_1/A vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M5061 NAND3X1_5/a_9_6# OAI21X1_1/A gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M5062 NOR2X1_59/B OAI21X1_1/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5063 NOR2X1_59/B OAI21X1_1/B NAND3X1_5/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M5064 vdd INVX2_30/Y NOR2X1_59/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5065 NAND3X1_5/a_14_6# INVX2_30/Y NAND3X1_5/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M5066 DFFNEGX1_107/a_76_6# BUFX2_9/Y DFFNEGX1_107/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M5067 gnd BUFX2_9/Y DFFNEGX1_107/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5068 DFFNEGX1_107/a_66_6# DFFNEGX1_107/a_2_6# DFFNEGX1_107/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5069 out_global_score[13] DFFNEGX1_107/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5070 DFFNEGX1_107/a_23_6# BUFX2_9/Y DFFNEGX1_107/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M5071 DFFNEGX1_107/a_23_6# DFFNEGX1_107/a_2_6# DFFNEGX1_107/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M5072 gnd DFFNEGX1_107/a_34_4# DFFNEGX1_107/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5073 vdd DFFNEGX1_107/a_34_4# DFFNEGX1_107/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M5074 DFFNEGX1_107/a_61_74# DFFNEGX1_107/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5075 DFFNEGX1_107/a_34_4# DFFNEGX1_107/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5076 DFFNEGX1_107/a_34_4# DFFNEGX1_107/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M5077 vdd out_global_score[13] DFFNEGX1_107/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5078 gnd out_global_score[13] DFFNEGX1_107/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5079 DFFNEGX1_107/a_61_6# DFFNEGX1_107/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5080 DFFNEGX1_107/a_76_84# DFFNEGX1_107/a_2_6# DFFNEGX1_107/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M5081 out_global_score[13] DFFNEGX1_107/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5082 vdd BUFX2_9/Y DFFNEGX1_107/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M5083 DFFNEGX1_107/a_31_6# DFFNEGX1_107/a_2_6# DFFNEGX1_107/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5084 DFFNEGX1_107/a_66_6# BUFX2_9/Y DFFNEGX1_107/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5085 DFFNEGX1_107/a_17_74# INVX2_203/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5086 DFFNEGX1_107/a_31_74# BUFX2_9/Y DFFNEGX1_107/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5087 DFFNEGX1_107/a_17_6# INVX2_203/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5088 DFFNEGX1_118/a_76_6# BUFX2_9/Y DFFNEGX1_118/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M5089 gnd BUFX2_9/Y DFFNEGX1_118/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5090 DFFNEGX1_118/a_66_6# DFFNEGX1_118/a_2_6# DFFNEGX1_118/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5091 out_global_score[24] DFFNEGX1_118/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5092 DFFNEGX1_118/a_23_6# BUFX2_9/Y DFFNEGX1_118/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M5093 DFFNEGX1_118/a_23_6# DFFNEGX1_118/a_2_6# DFFNEGX1_118/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M5094 gnd DFFNEGX1_118/a_34_4# DFFNEGX1_118/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5095 vdd DFFNEGX1_118/a_34_4# DFFNEGX1_118/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M5096 DFFNEGX1_118/a_61_74# DFFNEGX1_118/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5097 DFFNEGX1_118/a_34_4# DFFNEGX1_118/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5098 DFFNEGX1_118/a_34_4# DFFNEGX1_118/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M5099 vdd out_global_score[24] DFFNEGX1_118/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5100 gnd out_global_score[24] DFFNEGX1_118/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5101 DFFNEGX1_118/a_61_6# DFFNEGX1_118/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5102 DFFNEGX1_118/a_76_84# DFFNEGX1_118/a_2_6# DFFNEGX1_118/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M5103 out_global_score[24] DFFNEGX1_118/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5104 vdd BUFX2_9/Y DFFNEGX1_118/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M5105 DFFNEGX1_118/a_31_6# DFFNEGX1_118/a_2_6# DFFNEGX1_118/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5106 DFFNEGX1_118/a_66_6# BUFX2_9/Y DFFNEGX1_118/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5107 DFFNEGX1_118/a_17_74# INVX2_192/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5108 DFFNEGX1_118/a_31_74# BUFX2_9/Y DFFNEGX1_118/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5109 DFFNEGX1_118/a_17_6# INVX2_192/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5110 DFFNEGX1_129/a_76_6# INVX2_259/Y DFFNEGX1_129/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M5111 gnd INVX2_259/Y DFFNEGX1_129/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5112 DFFNEGX1_129/a_66_6# DFFNEGX1_129/a_2_6# DFFNEGX1_129/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5113 out_alu_done DFFNEGX1_129/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5114 DFFNEGX1_129/a_23_6# INVX2_259/Y DFFNEGX1_129/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M5115 DFFNEGX1_129/a_23_6# DFFNEGX1_129/a_2_6# DFFNEGX1_129/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M5116 gnd DFFNEGX1_129/a_34_4# DFFNEGX1_129/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5117 vdd DFFNEGX1_129/a_34_4# DFFNEGX1_129/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M5118 DFFNEGX1_129/a_61_74# DFFNEGX1_129/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5119 DFFNEGX1_129/a_34_4# DFFNEGX1_129/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5120 DFFNEGX1_129/a_34_4# DFFNEGX1_129/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M5121 vdd out_alu_done DFFNEGX1_129/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5122 gnd out_alu_done DFFNEGX1_129/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5123 DFFNEGX1_129/a_61_6# DFFNEGX1_129/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5124 DFFNEGX1_129/a_76_84# DFFNEGX1_129/a_2_6# DFFNEGX1_129/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M5125 out_alu_done DFFNEGX1_129/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5126 vdd INVX2_259/Y DFFNEGX1_129/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M5127 DFFNEGX1_129/a_31_6# DFFNEGX1_129/a_2_6# DFFNEGX1_129/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5128 DFFNEGX1_129/a_66_6# INVX2_259/Y DFFNEGX1_129/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5129 DFFNEGX1_129/a_17_74# OAI21X1_58/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5130 DFFNEGX1_129/a_31_74# INVX2_259/Y DFFNEGX1_129/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5131 DFFNEGX1_129/a_17_6# OAI21X1_58/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5132 gnd INVX2_61/Y OAI21X1_101/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M5133 vdd NAND2X1_88/Y OAI21X1_101/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M5134 OAI21X1_101/Y NAND2X1_88/Y OAI21X1_101/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5135 OAI21X1_101/Y BUFX2_23/Y OAI21X1_101/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5136 OAI21X1_101/a_9_54# INVX2_61/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5137 OAI21X1_101/a_2_6# BUFX2_23/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5138 gnd INVX2_19/Y OAI21X1_112/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M5139 vdd AOI22X1_55/Y AOI22X1_54/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M5140 AOI22X1_54/B AOI22X1_55/Y OAI21X1_112/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5141 AOI22X1_54/B OAI22X1_38/C OAI21X1_112/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5142 OAI21X1_112/a_9_54# INVX2_19/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5143 OAI21X1_112/a_2_6# OAI22X1_38/C gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5144 gnd OAI22X1_74/Y OAI21X1_145/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M5145 vdd INVX2_38/Y OAI21X1_145/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M5146 OAI21X1_145/Y INVX2_38/Y OAI21X1_145/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5147 OAI21X1_145/Y OAI22X1_73/Y OAI21X1_145/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5148 OAI21X1_145/a_9_54# OAI22X1_74/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5149 OAI21X1_145/a_2_6# OAI22X1_73/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5150 gnd INVX2_120/A OAI21X1_156/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M5151 vdd out_display OAI21X1_156/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M5152 OAI21X1_156/Y out_display OAI21X1_156/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5153 OAI21X1_156/Y INVX2_121/A OAI21X1_156/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5154 OAI21X1_156/a_9_54# INVX2_120/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5155 OAI21X1_156/a_2_6# INVX2_121/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5156 gnd OAI22X1_56/Y OAI21X1_134/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M5157 vdd OAI21X1_1/B AOI21X1_13/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M5158 AOI21X1_13/A OAI21X1_1/B OAI21X1_134/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5159 AOI21X1_13/A OAI22X1_55/Y OAI21X1_134/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5160 OAI21X1_134/a_9_54# OAI22X1_56/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5161 OAI21X1_134/a_2_6# OAI22X1_55/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5162 gnd AOI22X1_72/Y OAI21X1_123/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M5163 vdd OAI21X1_124/Y XOR2X1_25/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M5164 XOR2X1_25/B OAI21X1_124/Y OAI21X1_123/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5165 XOR2X1_25/B XNOR2X1_21/Y OAI21X1_123/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5166 OAI21X1_123/a_9_54# AOI22X1_72/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5167 OAI21X1_123/a_2_6# XNOR2X1_21/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5168 gnd out_global_score[15] AOI22X1_18/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M5169 INVX2_201/A INVX2_257/Y AOI22X1_18/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M5170 AOI22X1_18/a_11_6# HAX1_15/YS gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5171 AOI22X1_18/a_2_54# INVX2_257/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M5172 AOI22X1_18/a_28_6# OR2X1_11/B INVX2_201/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5173 vdd HAX1_15/YS AOI22X1_18/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5174 INVX2_201/A OR2X1_11/B AOI22X1_18/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M5175 AOI22X1_18/a_2_54# out_global_score[15] INVX2_201/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5176 gnd out_global_score[4] AOI22X1_29/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M5177 INVX2_212/A INVX2_258/Y AOI22X1_29/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M5178 AOI22X1_29/a_11_6# HAX1_26/YS gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5179 AOI22X1_29/a_2_54# INVX2_258/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M5180 AOI22X1_29/a_28_6# OR2X1_11/B INVX2_212/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5181 vdd HAX1_26/YS AOI22X1_29/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5182 INVX2_212/A OR2X1_11/B AOI22X1_29/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M5183 AOI22X1_29/a_2_54# out_global_score[4] INVX2_212/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5184 vdd out_global_score[9] HAX1_21/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M5185 HAX1_21/a_41_74# HAX1_21/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M5186 HAX1_21/a_9_6# out_global_score[9] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5187 HAX1_21/a_41_74# HAX1_21/B HAX1_21/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M5188 vdd out_global_score[9] HAX1_21/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5189 vdd HAX1_21/a_2_74# HAX1_20/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5190 HAX1_21/a_38_6# HAX1_21/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5191 HAX1_21/YS HAX1_21/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5192 HAX1_21/a_38_6# out_global_score[9] HAX1_21/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5193 HAX1_21/YS HAX1_21/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M5194 HAX1_21/a_2_74# HAX1_21/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5195 HAX1_21/a_2_74# HAX1_21/B HAX1_21/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5196 HAX1_21/a_49_54# HAX1_21/B HAX1_21/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5197 gnd HAX1_21/a_2_74# HAX1_20/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M5198 vdd HAX1_32/A HAX1_32/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M5199 HAX1_32/a_41_74# HAX1_32/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M5200 HAX1_32/a_9_6# HAX1_32/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5201 HAX1_32/a_41_74# HAX1_32/B HAX1_32/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M5202 vdd HAX1_32/A HAX1_32/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5203 vdd HAX1_32/a_2_74# FAX1_15/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5204 HAX1_32/a_38_6# HAX1_32/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5205 FAX1_16/B HAX1_32/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5206 HAX1_32/a_38_6# HAX1_32/A HAX1_32/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5207 FAX1_16/B HAX1_32/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M5208 HAX1_32/a_2_74# HAX1_32/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5209 HAX1_32/a_2_74# HAX1_32/B HAX1_32/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5210 HAX1_32/a_49_54# HAX1_32/B HAX1_32/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5211 gnd HAX1_32/a_2_74# FAX1_15/C Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M5212 vdd out_global_score[20] HAX1_10/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M5213 HAX1_10/a_41_74# HAX1_10/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M5214 HAX1_10/a_9_6# out_global_score[20] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5215 HAX1_10/a_41_74# HAX1_10/B HAX1_10/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M5216 vdd out_global_score[20] HAX1_10/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5217 vdd HAX1_10/a_2_74# HAX1_9/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5218 HAX1_10/a_38_6# HAX1_10/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5219 HAX1_10/YS HAX1_10/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5220 HAX1_10/a_38_6# out_global_score[20] HAX1_10/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5221 HAX1_10/YS HAX1_10/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M5222 HAX1_10/a_2_74# HAX1_10/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5223 HAX1_10/a_2_74# HAX1_10/B HAX1_10/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5224 HAX1_10/a_49_54# HAX1_10/B HAX1_10/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5225 gnd HAX1_10/a_2_74# HAX1_9/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M5226 vdd HAX1_43/A HAX1_43/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M5227 HAX1_43/a_41_74# HAX1_43/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M5228 HAX1_43/a_9_6# HAX1_43/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5229 HAX1_43/a_41_74# HAX1_43/B HAX1_43/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M5230 vdd HAX1_43/A HAX1_43/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5231 vdd HAX1_43/a_2_74# OR2X1_3/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5232 HAX1_43/a_38_6# HAX1_43/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5233 HAX1_43/YS HAX1_43/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5234 HAX1_43/a_38_6# HAX1_43/A HAX1_43/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5235 HAX1_43/YS HAX1_43/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M5236 HAX1_43/a_2_74# HAX1_43/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5237 HAX1_43/a_2_74# HAX1_43/B HAX1_43/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5238 HAX1_43/a_49_54# HAX1_43/B HAX1_43/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5239 gnd HAX1_43/a_2_74# OR2X1_3/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M5240 gnd out_temp_data_in[0] OAI21X1_2/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M5241 vdd out_temp_data_in[3] OAI21X1_2/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M5242 OAI21X1_2/Y out_temp_data_in[3] OAI21X1_2/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5243 OAI21X1_2/Y out_temp_data_in[1] OAI21X1_2/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5244 OAI21X1_2/a_9_54# out_temp_data_in[0] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5245 OAI21X1_2/a_2_6# out_temp_data_in[1] gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5246 gnd out_mines[9] OAI22X1_70/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M5247 OAI22X1_70/a_2_6# out_mines[8] OAI22X1_70/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M5248 OAI22X1_70/Y OAI22X1_76/D OAI22X1_70/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5249 OAI22X1_70/Y OAI22X1_76/B OAI22X1_70/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M5250 OAI22X1_70/a_28_54# OAI22X1_76/D OAI22X1_70/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M5251 OAI22X1_70/a_9_54# out_mines[9] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5252 OAI22X1_70/a_2_6# OAI22X1_76/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5253 vdd out_mines[8] OAI22X1_70/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5254 gnd out_mines[11] OAI22X1_81/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M5255 OAI22X1_81/a_2_6# out_mines[10] OAI22X1_81/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M5256 OAI22X1_81/Y OAI22X1_87/D OAI22X1_81/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5257 OAI22X1_81/Y OAI22X1_87/B OAI22X1_81/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M5258 OAI22X1_81/a_28_54# OAI22X1_87/D OAI22X1_81/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M5259 OAI22X1_81/a_9_54# out_mines[11] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5260 OAI22X1_81/a_2_6# OAI22X1_87/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5261 vdd out_mines[10] OAI22X1_81/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5262 DFFNEGX1_0/a_76_6# INVX2_259/Y DFFNEGX1_0/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M5263 gnd INVX2_259/Y DFFNEGX1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5264 DFFNEGX1_0/a_66_6# DFFNEGX1_0/a_2_6# DFFNEGX1_0/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5265 INVX2_0/A DFFNEGX1_0/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5266 DFFNEGX1_0/a_23_6# INVX2_259/Y DFFNEGX1_0/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M5267 DFFNEGX1_0/a_23_6# DFFNEGX1_0/a_2_6# DFFNEGX1_0/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M5268 gnd DFFNEGX1_0/a_34_4# DFFNEGX1_0/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5269 vdd DFFNEGX1_0/a_34_4# DFFNEGX1_0/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M5270 DFFNEGX1_0/a_61_74# DFFNEGX1_0/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5271 DFFNEGX1_0/a_34_4# DFFNEGX1_0/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5272 DFFNEGX1_0/a_34_4# DFFNEGX1_0/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M5273 vdd INVX2_0/A DFFNEGX1_0/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5274 gnd INVX2_0/A DFFNEGX1_0/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5275 DFFNEGX1_0/a_61_6# DFFNEGX1_0/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5276 DFFNEGX1_0/a_76_84# DFFNEGX1_0/a_2_6# DFFNEGX1_0/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M5277 INVX2_0/A DFFNEGX1_0/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5278 vdd INVX2_259/Y DFFNEGX1_0/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M5279 DFFNEGX1_0/a_31_6# DFFNEGX1_0/a_2_6# DFFNEGX1_0/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5280 DFFNEGX1_0/a_66_6# INVX2_259/Y DFFNEGX1_0/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5281 DFFNEGX1_0/a_17_74# OAI21X1_57/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5282 DFFNEGX1_0/a_31_74# INVX2_259/Y DFFNEGX1_0/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5283 DFFNEGX1_0/a_17_6# OAI21X1_57/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5284 gnd XOR2X1_5/A XOR2X1_5/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5285 XOR2X1_5/Y XOR2X1_5/a_2_6# XOR2X1_5/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M5286 XOR2X1_5/a_13_43# FAX1_4/YC gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5287 XOR2X1_5/a_18_54# XOR2X1_5/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M5288 XOR2X1_5/a_35_6# XOR2X1_5/A XOR2X1_5/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5289 XOR2X1_5/a_18_6# XOR2X1_5/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5290 vdd XOR2X1_5/A XOR2X1_5/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M5291 vdd FAX1_4/YC XOR2X1_5/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5292 XOR2X1_5/Y XOR2X1_5/A XOR2X1_5/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M5293 XOR2X1_5/a_35_54# XOR2X1_5/a_2_6# XOR2X1_5/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5294 XOR2X1_5/a_13_43# FAX1_4/YC vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5295 gnd FAX1_4/YC XOR2X1_5/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5296 gnd MUX2X1_6/A MUX2X1_6/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M5297 MUX2X1_6/a_17_50# HAX1_38/A vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M5298 MUX2X1_6/Y OR2X1_5/Y MUX2X1_6/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M5299 MUX2X1_6/a_30_54# MUX2X1_6/a_2_10# MUX2X1_6/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M5300 MUX2X1_6/a_17_10# HAX1_38/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5301 vdd OR2X1_5/Y MUX2X1_6/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5302 MUX2X1_6/a_30_10# OR2X1_5/Y MUX2X1_6/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M5303 gnd OR2X1_5/Y MUX2X1_6/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M5304 vdd MUX2X1_6/A MUX2X1_6/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5305 MUX2X1_6/Y MUX2X1_6/a_2_10# MUX2X1_6/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5306 INVX2_101/Y out_temp_cleared[12] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5307 INVX2_101/Y out_temp_cleared[12] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5308 OAI22X1_3/B out_temp_cleared[1] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5309 OAI22X1_3/B out_temp_cleared[1] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5310 INVX2_123/Y INVX2_123/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5311 INVX2_123/Y INVX2_123/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5312 MUX2X1_12/B MUX2X1_8/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5313 MUX2X1_12/B MUX2X1_8/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5314 MUX2X1_4/A XOR2X1_8/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5315 MUX2X1_4/A XOR2X1_8/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5316 NOR2X1_9/A in_mult[0] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5317 NOR2X1_9/A in_mult[0] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5318 OR2X1_1/A MUX2X1_20/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5319 OR2X1_1/A MUX2X1_20/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5320 NOR2X1_64/A OR2X1_12/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5321 NOR2X1_64/A OR2X1_12/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5322 INVX2_189/Y INVX2_189/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5323 INVX2_189/Y INVX2_189/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5324 DFFNEGX1_18/a_76_6# BUFX2_16/Y DFFNEGX1_18/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M5325 gnd BUFX2_16/Y DFFNEGX1_18/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5326 DFFNEGX1_18/a_66_6# DFFNEGX1_18/a_2_6# DFFNEGX1_18/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5327 out_mines[23] DFFNEGX1_18/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5328 DFFNEGX1_18/a_23_6# BUFX2_16/Y DFFNEGX1_18/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M5329 DFFNEGX1_18/a_23_6# DFFNEGX1_18/a_2_6# DFFNEGX1_18/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M5330 gnd DFFNEGX1_18/a_34_4# DFFNEGX1_18/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5331 vdd DFFNEGX1_18/a_34_4# DFFNEGX1_18/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M5332 DFFNEGX1_18/a_61_74# DFFNEGX1_18/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5333 DFFNEGX1_18/a_34_4# DFFNEGX1_18/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5334 DFFNEGX1_18/a_34_4# DFFNEGX1_18/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M5335 vdd out_mines[23] DFFNEGX1_18/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5336 gnd out_mines[23] DFFNEGX1_18/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5337 DFFNEGX1_18/a_61_6# DFFNEGX1_18/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5338 DFFNEGX1_18/a_76_84# DFFNEGX1_18/a_2_6# DFFNEGX1_18/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M5339 out_mines[23] DFFNEGX1_18/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5340 vdd BUFX2_16/Y DFFNEGX1_18/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M5341 DFFNEGX1_18/a_31_6# DFFNEGX1_18/a_2_6# DFFNEGX1_18/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5342 DFFNEGX1_18/a_66_6# BUFX2_16/Y DFFNEGX1_18/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5343 DFFNEGX1_18/a_17_74# OAI21X1_5/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5344 DFFNEGX1_18/a_31_74# BUFX2_16/Y DFFNEGX1_18/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5345 DFFNEGX1_18/a_17_6# OAI21X1_5/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5346 DFFNEGX1_29/a_76_6# BUFX2_15/Y DFFNEGX1_29/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M5347 gnd BUFX2_15/Y DFFNEGX1_29/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5348 DFFNEGX1_29/a_66_6# DFFNEGX1_29/a_2_6# DFFNEGX1_29/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5349 out_mines[3] DFFNEGX1_29/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5350 DFFNEGX1_29/a_23_6# BUFX2_15/Y DFFNEGX1_29/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M5351 DFFNEGX1_29/a_23_6# DFFNEGX1_29/a_2_6# DFFNEGX1_29/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M5352 gnd DFFNEGX1_29/a_34_4# DFFNEGX1_29/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5353 vdd DFFNEGX1_29/a_34_4# DFFNEGX1_29/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M5354 DFFNEGX1_29/a_61_74# DFFNEGX1_29/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5355 DFFNEGX1_29/a_34_4# DFFNEGX1_29/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5356 DFFNEGX1_29/a_34_4# DFFNEGX1_29/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M5357 vdd out_mines[3] DFFNEGX1_29/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5358 gnd out_mines[3] DFFNEGX1_29/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5359 DFFNEGX1_29/a_61_6# DFFNEGX1_29/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5360 DFFNEGX1_29/a_76_84# DFFNEGX1_29/a_2_6# DFFNEGX1_29/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M5361 out_mines[3] DFFNEGX1_29/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5362 vdd BUFX2_15/Y DFFNEGX1_29/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M5363 DFFNEGX1_29/a_31_6# DFFNEGX1_29/a_2_6# DFFNEGX1_29/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5364 DFFNEGX1_29/a_66_6# BUFX2_15/Y DFFNEGX1_29/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5365 DFFNEGX1_29/a_17_74# OAI21X1_45/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5366 DFFNEGX1_29/a_31_74# BUFX2_15/Y DFFNEGX1_29/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5367 DFFNEGX1_29/a_17_6# OAI21X1_45/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5368 gnd XOR2X1_17/Y XOR2X1_16/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5369 XOR2X1_16/Y XOR2X1_16/a_2_6# XOR2X1_16/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M5370 XOR2X1_16/a_13_43# INVX2_45/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5371 XOR2X1_16/a_18_54# XOR2X1_16/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M5372 XOR2X1_16/a_35_6# XOR2X1_17/Y XOR2X1_16/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5373 XOR2X1_16/a_18_6# XOR2X1_16/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5374 vdd XOR2X1_17/Y XOR2X1_16/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M5375 vdd INVX2_45/A XOR2X1_16/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5376 XOR2X1_16/Y XOR2X1_17/Y XOR2X1_16/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M5377 XOR2X1_16/a_35_54# XOR2X1_16/a_2_6# XOR2X1_16/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5378 XOR2X1_16/a_13_43# INVX2_45/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5379 gnd INVX2_45/A XOR2X1_16/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5380 gnd XOR2X1_28/Y XOR2X1_27/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5381 XOR2X1_27/Y XOR2X1_27/a_2_6# XOR2X1_27/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M5382 XOR2X1_27/a_13_43# INVX2_44/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5383 XOR2X1_27/a_18_54# XOR2X1_27/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M5384 XOR2X1_27/a_35_6# XOR2X1_28/Y XOR2X1_27/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5385 XOR2X1_27/a_18_6# XOR2X1_27/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5386 vdd XOR2X1_28/Y XOR2X1_27/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M5387 vdd INVX2_44/A XOR2X1_27/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5388 XOR2X1_27/Y XOR2X1_28/Y XOR2X1_27/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M5389 XOR2X1_27/a_35_54# XOR2X1_27/a_2_6# XOR2X1_27/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5390 XOR2X1_27/a_13_43# INVX2_44/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5391 gnd INVX2_44/A XOR2X1_27/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5392 DFFNEGX1_108/a_76_6# BUFX2_9/Y DFFNEGX1_108/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M5393 gnd BUFX2_9/Y DFFNEGX1_108/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5394 DFFNEGX1_108/a_66_6# DFFNEGX1_108/a_2_6# DFFNEGX1_108/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5395 out_global_score[14] DFFNEGX1_108/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5396 DFFNEGX1_108/a_23_6# BUFX2_9/Y DFFNEGX1_108/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M5397 DFFNEGX1_108/a_23_6# DFFNEGX1_108/a_2_6# DFFNEGX1_108/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M5398 gnd DFFNEGX1_108/a_34_4# DFFNEGX1_108/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5399 vdd DFFNEGX1_108/a_34_4# DFFNEGX1_108/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M5400 DFFNEGX1_108/a_61_74# DFFNEGX1_108/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5401 DFFNEGX1_108/a_34_4# DFFNEGX1_108/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5402 DFFNEGX1_108/a_34_4# DFFNEGX1_108/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M5403 vdd out_global_score[14] DFFNEGX1_108/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5404 gnd out_global_score[14] DFFNEGX1_108/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5405 DFFNEGX1_108/a_61_6# DFFNEGX1_108/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5406 DFFNEGX1_108/a_76_84# DFFNEGX1_108/a_2_6# DFFNEGX1_108/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M5407 out_global_score[14] DFFNEGX1_108/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5408 vdd BUFX2_9/Y DFFNEGX1_108/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M5409 DFFNEGX1_108/a_31_6# DFFNEGX1_108/a_2_6# DFFNEGX1_108/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5410 DFFNEGX1_108/a_66_6# BUFX2_9/Y DFFNEGX1_108/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5411 DFFNEGX1_108/a_17_74# INVX2_202/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5412 DFFNEGX1_108/a_31_74# BUFX2_9/Y DFFNEGX1_108/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5413 DFFNEGX1_108/a_17_6# INVX2_202/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5414 NAND3X1_6/Y out_start vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M5415 NAND3X1_6/a_9_6# out_start gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M5416 NAND3X1_6/Y out_place_done vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5417 NAND3X1_6/Y out_place_done NAND3X1_6/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M5418 vdd AND2X2_8/A NAND3X1_6/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5419 NAND3X1_6/a_14_6# AND2X2_8/A NAND3X1_6/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M5420 DFFNEGX1_119/a_76_6# BUFX2_5/Y DFFNEGX1_119/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M5421 gnd BUFX2_5/Y DFFNEGX1_119/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5422 DFFNEGX1_119/a_66_6# DFFNEGX1_119/a_2_6# DFFNEGX1_119/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5423 out_global_score[25] DFFNEGX1_119/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5424 DFFNEGX1_119/a_23_6# BUFX2_5/Y DFFNEGX1_119/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M5425 DFFNEGX1_119/a_23_6# DFFNEGX1_119/a_2_6# DFFNEGX1_119/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M5426 gnd DFFNEGX1_119/a_34_4# DFFNEGX1_119/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5427 vdd DFFNEGX1_119/a_34_4# DFFNEGX1_119/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M5428 DFFNEGX1_119/a_61_74# DFFNEGX1_119/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5429 DFFNEGX1_119/a_34_4# DFFNEGX1_119/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5430 DFFNEGX1_119/a_34_4# DFFNEGX1_119/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M5431 vdd out_global_score[25] DFFNEGX1_119/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5432 gnd out_global_score[25] DFFNEGX1_119/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5433 DFFNEGX1_119/a_61_6# DFFNEGX1_119/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5434 DFFNEGX1_119/a_76_84# DFFNEGX1_119/a_2_6# DFFNEGX1_119/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M5435 out_global_score[25] DFFNEGX1_119/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5436 vdd BUFX2_5/Y DFFNEGX1_119/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M5437 DFFNEGX1_119/a_31_6# DFFNEGX1_119/a_2_6# DFFNEGX1_119/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5438 DFFNEGX1_119/a_66_6# BUFX2_5/Y DFFNEGX1_119/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5439 DFFNEGX1_119/a_17_74# INVX2_191/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5440 DFFNEGX1_119/a_31_74# BUFX2_5/Y DFFNEGX1_119/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5441 DFFNEGX1_119/a_17_6# INVX2_191/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5442 gnd INVX2_60/Y OAI21X1_102/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M5443 vdd NAND2X1_89/Y OAI21X1_102/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M5444 OAI21X1_102/Y NAND2X1_89/Y OAI21X1_102/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5445 OAI21X1_102/Y BUFX2_23/Y OAI21X1_102/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5446 OAI21X1_102/a_9_54# INVX2_60/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5447 OAI21X1_102/a_2_6# BUFX2_23/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5448 gnd INVX2_33/Y OAI21X1_113/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M5449 vdd OAI21X1_114/Y AOI22X1_57/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M5450 AOI22X1_57/A OAI21X1_114/Y OAI21X1_113/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5451 AOI22X1_57/A INVX2_251/Y OAI21X1_113/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5452 OAI21X1_113/a_9_54# INVX2_33/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5453 OAI21X1_113/a_2_6# INVX2_251/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5454 gnd OAI22X1_76/Y OAI21X1_146/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M5455 vdd XOR2X1_3/Y OAI21X1_146/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M5456 OAI21X1_146/Y XOR2X1_3/Y OAI21X1_146/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5457 OAI21X1_146/Y OAI22X1_75/Y OAI21X1_146/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5458 OAI21X1_146/a_9_54# OAI22X1_76/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5459 OAI21X1_146/a_2_6# OAI22X1_75/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5460 gnd OAI22X1_58/Y OAI21X1_135/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M5461 vdd out_temp_data_in[2] AOI21X1_14/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M5462 AOI21X1_14/B out_temp_data_in[2] OAI21X1_135/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5463 AOI21X1_14/B OAI22X1_57/Y OAI21X1_135/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5464 OAI21X1_135/a_9_54# OAI22X1_58/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5465 OAI21X1_135/a_2_6# OAI22X1_57/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5466 gnd AOI21X1_12/Y OAI21X1_124/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M5467 vdd XNOR2X1_21/Y OAI21X1_124/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M5468 OAI21X1_124/Y XNOR2X1_21/Y OAI21X1_124/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5469 OAI21X1_124/Y AOI21X1_11/Y OAI21X1_124/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5470 OAI21X1_124/a_9_54# AOI21X1_12/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5471 OAI21X1_124/a_2_6# AOI21X1_11/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5472 gnd OAI21X1_157/A OAI21X1_157/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M5473 vdd OR2X1_15/Y OAI21X1_157/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M5474 OAI21X1_157/Y OR2X1_15/Y OAI21X1_157/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5475 OAI21X1_157/Y OAI21X1_157/B OAI21X1_157/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5476 OAI21X1_157/a_9_54# OAI21X1_157/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5477 OAI21X1_157/a_2_6# OAI21X1_157/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5478 vdd in_clka BUFX2_0/a_2_6# vdd pfet w=20 l=2
+  ad=0.11n pd=46u as=100p ps=50u
M5479 gnd in_clka BUFX2_0/a_2_6# Gnd nfet w=10 l=2
+  ad=55p pd=26u as=50p ps=30u
M5480 BUFX2_9/A BUFX2_0/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.11n ps=46u
M5481 BUFX2_9/A BUFX2_0/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=55p ps=26u
M5482 OAI21X1_157/A INVX2_119/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M5483 NAND2X1_130/a_9_6# INVX2_119/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5484 vdd INVX2_117/Y OAI21X1_157/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5485 OAI21X1_157/A INVX2_117/Y NAND2X1_130/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5486 INVX2_0/Y INVX2_0/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5487 INVX2_0/Y INVX2_0/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5488 gnd out_global_score[14] AOI22X1_19/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M5489 INVX2_202/A INVX2_257/Y AOI22X1_19/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M5490 AOI22X1_19/a_11_6# HAX1_16/YS gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5491 AOI22X1_19/a_2_54# INVX2_257/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M5492 AOI22X1_19/a_28_6# OR2X1_11/B INVX2_202/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5493 vdd HAX1_16/YS AOI22X1_19/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5494 INVX2_202/A OR2X1_11/B AOI22X1_19/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M5495 AOI22X1_19/a_2_54# out_global_score[14] INVX2_202/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5496 AOI21X1_0/a_2_54# out_temp_data_in[1] vdd vdd pfet w=40 l=2
+  ad=0.12n pd=46u as=0.12n ps=46u
M5497 AOI21X1_0/a_12_6# out_temp_data_in[0] gnd Gnd nfet w=20 l=2
+  ad=29.999998p pd=23u as=100p ps=50u
M5498 gnd OAI21X1_0/A INVX2_53/A Gnd nfet w=10 l=2
+  ad=50p pd=30u as=55p ps=26u
M5499 vdd out_temp_data_in[0] AOI21X1_0/a_2_54# vdd pfet w=40 l=2
+  ad=0.12n pd=46u as=0.2n ps=90u
M5500 INVX2_53/A OAI21X1_0/A AOI21X1_0/a_2_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=46u
M5501 INVX2_53/A out_temp_data_in[1] AOI21X1_0/a_12_6# Gnd nfet w=20 l=2
+  ad=55p pd=26u as=29.999998p ps=23u
M5502 gnd INVX2_120/Y XNOR2X1_30/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5503 INVX2_121/A INVX2_120/Y XNOR2X1_30/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M5504 XNOR2X1_30/a_12_41# INVX2_119/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5505 XNOR2X1_30/a_18_54# XNOR2X1_30/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M5506 XNOR2X1_30/a_35_6# XNOR2X1_30/a_2_6# INVX2_121/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5507 XNOR2X1_30/a_18_6# XNOR2X1_30/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5508 vdd INVX2_120/Y XNOR2X1_30/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M5509 vdd INVX2_119/A XNOR2X1_30/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5510 INVX2_121/A XNOR2X1_30/a_2_6# XNOR2X1_30/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M5511 XNOR2X1_30/a_35_54# INVX2_120/Y INVX2_121/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5512 XNOR2X1_30/a_12_41# INVX2_119/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5513 gnd INVX2_119/A XNOR2X1_30/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5514 vdd out_global_score[8] HAX1_22/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M5515 HAX1_22/a_41_74# HAX1_22/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M5516 HAX1_22/a_9_6# out_global_score[8] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5517 HAX1_22/a_41_74# HAX1_22/B HAX1_22/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M5518 vdd out_global_score[8] HAX1_22/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5519 vdd HAX1_22/a_2_74# HAX1_21/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5520 HAX1_22/a_38_6# HAX1_22/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5521 HAX1_22/YS HAX1_22/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5522 HAX1_22/a_38_6# out_global_score[8] HAX1_22/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5523 HAX1_22/YS HAX1_22/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M5524 HAX1_22/a_2_74# HAX1_22/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5525 HAX1_22/a_2_74# HAX1_22/B HAX1_22/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5526 HAX1_22/a_49_54# HAX1_22/B HAX1_22/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5527 gnd HAX1_22/a_2_74# HAX1_21/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M5528 vdd out_global_score[19] HAX1_11/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M5529 HAX1_11/a_41_74# HAX1_11/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M5530 HAX1_11/a_9_6# out_global_score[19] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5531 HAX1_11/a_41_74# HAX1_11/B HAX1_11/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M5532 vdd out_global_score[19] HAX1_11/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5533 vdd HAX1_11/a_2_74# HAX1_10/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5534 HAX1_11/a_38_6# HAX1_11/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5535 HAX1_11/YS HAX1_11/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5536 HAX1_11/a_38_6# out_global_score[19] HAX1_11/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5537 HAX1_11/YS HAX1_11/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M5538 HAX1_11/a_2_74# HAX1_11/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5539 HAX1_11/a_2_74# HAX1_11/B HAX1_11/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5540 HAX1_11/a_49_54# HAX1_11/B HAX1_11/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5541 gnd HAX1_11/a_2_74# HAX1_10/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M5542 vdd HAX1_44/A HAX1_44/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M5543 HAX1_44/a_41_74# HAX1_44/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M5544 HAX1_44/a_9_6# HAX1_44/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5545 HAX1_44/a_41_74# HAX1_44/B HAX1_44/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M5546 vdd HAX1_44/A HAX1_44/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5547 vdd HAX1_44/a_2_74# HAX1_45/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5548 HAX1_44/a_38_6# HAX1_44/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5549 HAX1_44/YS HAX1_44/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5550 HAX1_44/a_38_6# HAX1_44/A HAX1_44/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5551 HAX1_44/YS HAX1_44/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M5552 HAX1_44/a_2_74# HAX1_44/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5553 HAX1_44/a_2_74# HAX1_44/B HAX1_44/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5554 HAX1_44/a_49_54# HAX1_44/B HAX1_44/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5555 gnd HAX1_44/a_2_74# HAX1_45/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M5556 vdd HAX1_33/A HAX1_33/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M5557 HAX1_33/a_41_74# HAX1_33/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M5558 HAX1_33/a_9_6# HAX1_33/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5559 HAX1_33/a_41_74# HAX1_33/B HAX1_33/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M5560 vdd HAX1_33/A HAX1_33/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5561 vdd HAX1_33/a_2_74# FAX1_16/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5562 HAX1_33/a_38_6# HAX1_33/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5563 FAX1_9/A HAX1_33/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5564 HAX1_33/a_38_6# HAX1_33/A HAX1_33/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5565 FAX1_9/A HAX1_33/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M5566 HAX1_33/a_2_74# HAX1_33/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5567 HAX1_33/a_2_74# HAX1_33/B HAX1_33/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5568 HAX1_33/a_49_54# HAX1_33/B HAX1_33/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5569 gnd HAX1_33/a_2_74# FAX1_16/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M5570 gnd OAI21X1_3/A OAI21X1_3/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M5571 vdd OAI21X1_3/C OAI21X1_3/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M5572 OAI21X1_3/Y OAI21X1_3/C OAI21X1_3/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5573 OAI21X1_3/Y OAI21X1_9/B OAI21X1_3/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5574 OAI21X1_3/a_9_54# OAI21X1_3/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5575 OAI21X1_3/a_2_6# OAI21X1_9/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5576 gnd out_mines[13] OAI22X1_60/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M5577 OAI22X1_60/a_2_6# out_mines[12] OAI22X1_60/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M5578 OAI22X1_60/Y OAI22X1_64/D OAI22X1_60/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5579 OAI22X1_60/Y OAI22X1_64/B OAI22X1_60/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M5580 OAI22X1_60/a_28_54# OAI22X1_64/D OAI22X1_60/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M5581 OAI22X1_60/a_9_54# out_mines[13] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5582 OAI22X1_60/a_2_6# OAI22X1_64/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5583 vdd out_mines[12] OAI22X1_60/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5584 gnd out_mines[15] OAI22X1_71/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M5585 OAI22X1_71/a_2_6# out_mines[14] OAI22X1_71/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M5586 OAI22X1_71/Y OAI22X1_75/D OAI22X1_71/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5587 OAI22X1_71/Y OAI22X1_75/B OAI22X1_71/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M5588 OAI22X1_71/a_28_54# OAI22X1_75/D OAI22X1_71/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M5589 OAI22X1_71/a_9_54# out_mines[15] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5590 OAI22X1_71/a_2_6# OAI22X1_75/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5591 vdd out_mines[14] OAI22X1_71/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5592 gnd out_mines[9] OAI22X1_82/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M5593 OAI22X1_82/a_2_6# out_mines[8] OAI22X1_82/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M5594 OAI22X1_82/Y OAI22X1_88/D OAI22X1_82/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5595 OAI22X1_82/Y OAI22X1_88/B OAI22X1_82/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M5596 OAI22X1_82/a_28_54# OAI22X1_88/D OAI22X1_82/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M5597 OAI22X1_82/a_9_54# out_mines[9] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5598 OAI22X1_82/a_2_6# OAI22X1_88/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5599 vdd out_mines[8] OAI22X1_82/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5600 DFFNEGX1_1/a_76_6# BUFX2_17/Y DFFNEGX1_1/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M5601 gnd BUFX2_17/Y DFFNEGX1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5602 DFFNEGX1_1/a_66_6# DFFNEGX1_1/a_2_6# DFFNEGX1_1/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5603 out_temp_index[0] DFFNEGX1_1/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5604 DFFNEGX1_1/a_23_6# BUFX2_17/Y DFFNEGX1_1/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M5605 DFFNEGX1_1/a_23_6# DFFNEGX1_1/a_2_6# DFFNEGX1_1/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M5606 gnd DFFNEGX1_1/a_34_4# DFFNEGX1_1/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5607 vdd DFFNEGX1_1/a_34_4# DFFNEGX1_1/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M5608 DFFNEGX1_1/a_61_74# DFFNEGX1_1/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5609 DFFNEGX1_1/a_34_4# DFFNEGX1_1/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5610 DFFNEGX1_1/a_34_4# DFFNEGX1_1/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M5611 vdd out_temp_index[0] DFFNEGX1_1/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5612 gnd out_temp_index[0] DFFNEGX1_1/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5613 DFFNEGX1_1/a_61_6# DFFNEGX1_1/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5614 DFFNEGX1_1/a_76_84# DFFNEGX1_1/a_2_6# DFFNEGX1_1/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M5615 out_temp_index[0] DFFNEGX1_1/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5616 vdd BUFX2_17/Y DFFNEGX1_1/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M5617 DFFNEGX1_1/a_31_6# DFFNEGX1_1/a_2_6# DFFNEGX1_1/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5618 DFFNEGX1_1/a_66_6# BUFX2_17/Y DFFNEGX1_1/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5619 DFFNEGX1_1/a_17_74# OAI21X1_56/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5620 DFFNEGX1_1/a_31_74# BUFX2_17/Y DFFNEGX1_1/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5621 DFFNEGX1_1/a_17_6# OAI21X1_56/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5622 gnd XOR2X1_6/A XOR2X1_6/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5623 XOR2X1_6/Y XOR2X1_6/a_2_6# XOR2X1_6/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M5624 XOR2X1_6/a_13_43# FAX1_4/YS gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5625 XOR2X1_6/a_18_54# XOR2X1_6/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M5626 XOR2X1_6/a_35_6# XOR2X1_6/A XOR2X1_6/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5627 XOR2X1_6/a_18_6# XOR2X1_6/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5628 vdd XOR2X1_6/A XOR2X1_6/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M5629 vdd FAX1_4/YS XOR2X1_6/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5630 XOR2X1_6/Y XOR2X1_6/A XOR2X1_6/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M5631 XOR2X1_6/a_35_54# XOR2X1_6/a_2_6# XOR2X1_6/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5632 XOR2X1_6/a_13_43# FAX1_4/YS vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5633 gnd FAX1_4/YS XOR2X1_6/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5634 gnd MUX2X1_7/A MUX2X1_7/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M5635 MUX2X1_7/a_17_50# MUX2X1_7/B vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M5636 MUX2X1_7/Y OR2X1_5/Y MUX2X1_7/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M5637 MUX2X1_7/a_30_54# MUX2X1_7/a_2_10# MUX2X1_7/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M5638 MUX2X1_7/a_17_10# MUX2X1_7/B gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5639 vdd OR2X1_5/Y MUX2X1_7/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5640 MUX2X1_7/a_30_10# OR2X1_5/Y MUX2X1_7/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M5641 gnd OR2X1_5/Y MUX2X1_7/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M5642 vdd MUX2X1_7/A MUX2X1_7/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5643 MUX2X1_7/Y MUX2X1_7/a_2_10# MUX2X1_7/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5644 INVX2_102/Y out_temp_cleared[11] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5645 INVX2_102/Y out_temp_cleared[11] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5646 OAI22X1_3/D out_temp_cleared[0] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5647 OAI22X1_3/D out_temp_cleared[0] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5648 NAND2X1_6/B XOR2X1_6/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5649 NAND2X1_6/B XOR2X1_6/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5650 MUX2X1_34/A NOR2X1_0/B gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5651 MUX2X1_34/A NOR2X1_0/B vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5652 INVX2_124/Y INVX2_124/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5653 INVX2_124/Y INVX2_124/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5654 HAX1_47/A MUX2X1_21/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5655 HAX1_47/A MUX2X1_21/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5656 OR2X1_3/A MUX2X1_10/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5657 OR2X1_3/A MUX2X1_10/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5658 INVX2_179/Y NOR2X1_64/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5659 INVX2_179/Y NOR2X1_64/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5660 DFFNEGX1_19/a_76_6# BUFX2_16/Y DFFNEGX1_19/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M5661 gnd BUFX2_16/Y DFFNEGX1_19/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5662 DFFNEGX1_19/a_66_6# DFFNEGX1_19/a_2_6# DFFNEGX1_19/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5663 out_mines[21] DFFNEGX1_19/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5664 DFFNEGX1_19/a_23_6# BUFX2_16/Y DFFNEGX1_19/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M5665 DFFNEGX1_19/a_23_6# DFFNEGX1_19/a_2_6# DFFNEGX1_19/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M5666 gnd DFFNEGX1_19/a_34_4# DFFNEGX1_19/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5667 vdd DFFNEGX1_19/a_34_4# DFFNEGX1_19/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M5668 DFFNEGX1_19/a_61_74# DFFNEGX1_19/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5669 DFFNEGX1_19/a_34_4# DFFNEGX1_19/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5670 DFFNEGX1_19/a_34_4# DFFNEGX1_19/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M5671 vdd out_mines[21] DFFNEGX1_19/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5672 gnd out_mines[21] DFFNEGX1_19/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5673 DFFNEGX1_19/a_61_6# DFFNEGX1_19/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5674 DFFNEGX1_19/a_76_84# DFFNEGX1_19/a_2_6# DFFNEGX1_19/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M5675 out_mines[21] DFFNEGX1_19/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5676 vdd BUFX2_16/Y DFFNEGX1_19/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M5677 DFFNEGX1_19/a_31_6# DFFNEGX1_19/a_2_6# DFFNEGX1_19/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5678 DFFNEGX1_19/a_66_6# BUFX2_16/Y DFFNEGX1_19/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5679 DFFNEGX1_19/a_17_74# OAI21X1_9/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5680 DFFNEGX1_19/a_31_74# BUFX2_16/Y DFFNEGX1_19/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5681 DFFNEGX1_19/a_17_6# OAI21X1_9/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5682 gnd XOR2X1_18/Y XOR2X1_17/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5683 XOR2X1_17/Y XOR2X1_17/a_2_6# XOR2X1_17/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M5684 XOR2X1_17/a_13_43# INVX2_48/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5685 XOR2X1_17/a_18_54# XOR2X1_17/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M5686 XOR2X1_17/a_35_6# XOR2X1_18/Y XOR2X1_17/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5687 XOR2X1_17/a_18_6# XOR2X1_17/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5688 vdd XOR2X1_18/Y XOR2X1_17/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M5689 vdd INVX2_48/A XOR2X1_17/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5690 XOR2X1_17/Y XOR2X1_18/Y XOR2X1_17/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M5691 XOR2X1_17/a_35_54# XOR2X1_17/a_2_6# XOR2X1_17/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5692 XOR2X1_17/a_13_43# INVX2_48/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5693 gnd INVX2_48/A XOR2X1_17/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5694 gnd XOR2X1_28/A XOR2X1_28/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5695 XOR2X1_28/Y XOR2X1_28/a_2_6# XOR2X1_28/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M5696 XOR2X1_28/a_13_43# XOR2X1_29/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5697 XOR2X1_28/a_18_54# XOR2X1_28/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M5698 XOR2X1_28/a_35_6# XOR2X1_28/A XOR2X1_28/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5699 XOR2X1_28/a_18_6# XOR2X1_28/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5700 vdd XOR2X1_28/A XOR2X1_28/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M5701 vdd XOR2X1_29/Y XOR2X1_28/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5702 XOR2X1_28/Y XOR2X1_28/A XOR2X1_28/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M5703 XOR2X1_28/a_35_54# XOR2X1_28/a_2_6# XOR2X1_28/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5704 XOR2X1_28/a_13_43# XOR2X1_29/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5705 gnd XOR2X1_29/Y XOR2X1_28/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5706 NAND3X1_7/Y BUFX2_8/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M5707 NAND3X1_7/a_9_6# BUFX2_8/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M5708 NAND3X1_7/Y NAND3X1_7/C vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5709 NAND3X1_7/Y NAND3X1_7/C NAND3X1_7/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M5710 vdd NOR2X1_66/A NAND3X1_7/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5711 NAND3X1_7/a_14_6# NOR2X1_66/A NAND3X1_7/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M5712 DFFNEGX1_109/a_76_6# BUFX2_9/Y DFFNEGX1_109/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M5713 gnd BUFX2_9/Y DFFNEGX1_109/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5714 DFFNEGX1_109/a_66_6# DFFNEGX1_109/a_2_6# DFFNEGX1_109/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5715 out_global_score[15] DFFNEGX1_109/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5716 DFFNEGX1_109/a_23_6# BUFX2_9/Y DFFNEGX1_109/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M5717 DFFNEGX1_109/a_23_6# DFFNEGX1_109/a_2_6# DFFNEGX1_109/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M5718 gnd DFFNEGX1_109/a_34_4# DFFNEGX1_109/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5719 vdd DFFNEGX1_109/a_34_4# DFFNEGX1_109/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M5720 DFFNEGX1_109/a_61_74# DFFNEGX1_109/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5721 DFFNEGX1_109/a_34_4# DFFNEGX1_109/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5722 DFFNEGX1_109/a_34_4# DFFNEGX1_109/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M5723 vdd out_global_score[15] DFFNEGX1_109/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5724 gnd out_global_score[15] DFFNEGX1_109/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5725 DFFNEGX1_109/a_61_6# DFFNEGX1_109/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5726 DFFNEGX1_109/a_76_84# DFFNEGX1_109/a_2_6# DFFNEGX1_109/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M5727 out_global_score[15] DFFNEGX1_109/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5728 vdd BUFX2_9/Y DFFNEGX1_109/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M5729 DFFNEGX1_109/a_31_6# DFFNEGX1_109/a_2_6# DFFNEGX1_109/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5730 DFFNEGX1_109/a_66_6# BUFX2_9/Y DFFNEGX1_109/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5731 DFFNEGX1_109/a_17_74# INVX2_201/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5732 DFFNEGX1_109/a_31_74# BUFX2_9/Y DFFNEGX1_109/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5733 DFFNEGX1_109/a_17_6# INVX2_201/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5734 gnd INVX2_59/Y OAI21X1_103/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M5735 vdd NAND2X1_90/Y OAI21X1_103/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M5736 OAI21X1_103/Y NAND2X1_90/Y OAI21X1_103/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5737 OAI21X1_103/Y BUFX2_23/Y OAI21X1_103/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5738 OAI21X1_103/a_9_54# INVX2_59/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5739 OAI21X1_103/a_2_6# BUFX2_23/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5740 gnd OAI22X1_42/Y OAI21X1_125/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M5741 vdd INVX2_52/Y AOI21X1_11/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M5742 AOI21X1_11/B INVX2_52/Y OAI21X1_125/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5743 AOI21X1_11/B OAI22X1_41/Y OAI21X1_125/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5744 OAI21X1_125/a_9_54# OAI22X1_42/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5745 OAI21X1_125/a_2_6# OAI22X1_41/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5746 gnd NOR2X1_108/Y OAI21X1_114/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M5747 vdd INVX2_251/Y OAI21X1_114/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M5748 OAI21X1_114/Y INVX2_251/Y OAI21X1_114/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5749 OAI21X1_114/Y OAI22X1_39/Y OAI21X1_114/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5750 OAI21X1_114/a_9_54# NOR2X1_108/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5751 OAI21X1_114/a_2_6# OAI22X1_39/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5752 gnd AOI22X1_75/Y OAI21X1_147/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M5753 vdd OAI21X1_148/Y XOR2X1_28/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M5754 XOR2X1_28/A OAI21X1_148/Y OAI21X1_147/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5755 XOR2X1_28/A XOR2X1_12/Y OAI21X1_147/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5756 OAI21X1_147/a_9_54# AOI22X1_75/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5757 OAI21X1_147/a_2_6# XOR2X1_12/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5758 gnd OAI22X1_60/Y OAI21X1_136/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M5759 vdd OAI21X1_1/B AOI21X1_14/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M5760 AOI21X1_14/A OAI21X1_1/B OAI21X1_136/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5761 AOI21X1_14/A OAI22X1_59/Y OAI21X1_136/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5762 OAI21X1_136/a_9_54# OAI22X1_60/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5763 OAI21X1_136/a_2_6# OAI22X1_59/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5764 gnd INVX2_127/A OAI21X1_158/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M5765 vdd NAND3X1_50/Y OAI21X1_158/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M5766 OAI21X1_158/Y NAND3X1_50/Y OAI21X1_158/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5767 OAI21X1_158/Y OR2X1_15/A OAI21X1_158/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5768 OAI21X1_158/a_9_54# INVX2_127/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5769 OAI21X1_158/a_2_6# OR2X1_15/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5770 vdd in_clka BUFX2_1/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5771 gnd in_clka BUFX2_1/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M5772 BUFX2_1/Y BUFX2_1/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5773 BUFX2_1/Y BUFX2_1/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5774 AOI21X1_26/C INVX2_116/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M5775 NAND2X1_131/a_9_6# INVX2_116/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5776 vdd INVX2_118/Y AOI21X1_26/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5777 AOI21X1_26/C INVX2_118/Y NAND2X1_131/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5778 OAI22X1_75/D INVX2_37/A vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M5779 NAND2X1_120/a_9_6# INVX2_37/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5780 vdd out_temp_data_in[0] OAI22X1_75/D vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5781 OAI22X1_75/D out_temp_data_in[0] NAND2X1_120/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5782 INVX2_1/Y out_temp_index[0] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5783 INVX2_1/Y out_temp_index[0] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5784 AOI21X1_1/a_2_54# out_temp_index[2] vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M5785 AOI21X1_1/a_12_6# NOR2X1_67/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5786 gnd NOR2X1_66/Y INVX2_245/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0.11n ps=52u
M5787 vdd NOR2X1_67/Y AOI21X1_1/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5788 INVX2_245/A NOR2X1_66/Y AOI21X1_1/a_2_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5789 INVX2_245/A out_temp_index[2] AOI21X1_1/a_12_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5790 gnd XOR2X1_20/Y XNOR2X1_20/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5791 XNOR2X1_20/Y XOR2X1_20/Y XNOR2X1_20/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M5792 XNOR2X1_20/a_12_41# INVX2_48/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5793 XNOR2X1_20/a_18_54# XNOR2X1_20/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M5794 XNOR2X1_20/a_35_6# XNOR2X1_20/a_2_6# XNOR2X1_20/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5795 XNOR2X1_20/a_18_6# XNOR2X1_20/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5796 vdd XOR2X1_20/Y XNOR2X1_20/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M5797 vdd INVX2_48/Y XNOR2X1_20/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5798 XNOR2X1_20/Y XNOR2X1_20/a_2_6# XNOR2X1_20/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M5799 XNOR2X1_20/a_35_54# XOR2X1_20/Y XNOR2X1_20/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5800 XNOR2X1_20/a_12_41# INVX2_48/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5801 gnd INVX2_48/Y XNOR2X1_20/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5802 vdd out_global_score[18] HAX1_12/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M5803 HAX1_12/a_41_74# HAX1_12/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M5804 HAX1_12/a_9_6# out_global_score[18] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5805 HAX1_12/a_41_74# HAX1_12/B HAX1_12/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M5806 vdd out_global_score[18] HAX1_12/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5807 vdd HAX1_12/a_2_74# HAX1_11/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5808 HAX1_12/a_38_6# HAX1_12/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5809 HAX1_12/YS HAX1_12/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5810 HAX1_12/a_38_6# out_global_score[18] HAX1_12/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5811 HAX1_12/YS HAX1_12/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M5812 HAX1_12/a_2_74# HAX1_12/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5813 HAX1_12/a_2_74# HAX1_12/B HAX1_12/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5814 HAX1_12/a_49_54# HAX1_12/B HAX1_12/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5815 gnd HAX1_12/a_2_74# HAX1_11/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M5816 vdd out_global_score[7] HAX1_23/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M5817 HAX1_23/a_41_74# HAX1_23/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M5818 HAX1_23/a_9_6# out_global_score[7] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5819 HAX1_23/a_41_74# HAX1_23/B HAX1_23/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M5820 vdd out_global_score[7] HAX1_23/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5821 vdd HAX1_23/a_2_74# HAX1_22/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5822 HAX1_23/a_38_6# HAX1_23/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5823 HAX1_23/YS HAX1_23/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5824 HAX1_23/a_38_6# out_global_score[7] HAX1_23/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5825 HAX1_23/YS HAX1_23/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M5826 HAX1_23/a_2_74# HAX1_23/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5827 HAX1_23/a_2_74# HAX1_23/B HAX1_23/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5828 HAX1_23/a_49_54# HAX1_23/B HAX1_23/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5829 gnd HAX1_23/a_2_74# HAX1_22/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M5830 AOI21X1_20/a_2_54# INVX2_133/Y vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M5831 AOI21X1_20/a_12_6# AOI21X1_22/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5832 gnd BUFX2_3/Y AOI21X1_20/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0.11n ps=52u
M5833 vdd AOI21X1_22/Y AOI21X1_20/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5834 AOI21X1_20/Y BUFX2_3/Y AOI21X1_20/a_2_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5835 AOI21X1_20/Y INVX2_133/Y AOI21X1_20/a_12_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5836 vdd HAX1_45/A HAX1_45/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M5837 HAX1_45/a_41_74# HAX1_45/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M5838 HAX1_45/a_9_6# HAX1_45/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5839 HAX1_45/a_41_74# HAX1_45/B HAX1_45/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M5840 vdd HAX1_45/A HAX1_45/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5841 vdd HAX1_45/a_2_74# OR2X1_2/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5842 HAX1_45/a_38_6# HAX1_45/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5843 HAX1_45/YS HAX1_45/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5844 HAX1_45/a_38_6# HAX1_45/A HAX1_45/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5845 HAX1_45/YS HAX1_45/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M5846 HAX1_45/a_2_74# HAX1_45/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5847 HAX1_45/a_2_74# HAX1_45/B HAX1_45/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5848 HAX1_45/a_49_54# HAX1_45/B HAX1_45/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5849 gnd HAX1_45/a_2_74# OR2X1_2/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M5850 vdd HAX1_34/A HAX1_34/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M5851 HAX1_34/a_41_74# HAX1_34/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M5852 HAX1_34/a_9_6# HAX1_34/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5853 HAX1_34/a_41_74# HAX1_34/B HAX1_34/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M5854 vdd HAX1_34/A HAX1_34/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5855 vdd HAX1_34/a_2_74# FAX1_18/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5856 HAX1_34/a_38_6# HAX1_34/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5857 FAX1_10/C HAX1_34/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5858 HAX1_34/a_38_6# HAX1_34/A HAX1_34/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5859 FAX1_10/C HAX1_34/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M5860 HAX1_34/a_2_74# HAX1_34/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5861 HAX1_34/a_2_74# HAX1_34/B HAX1_34/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5862 HAX1_34/a_49_54# HAX1_34/B HAX1_34/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5863 gnd HAX1_34/a_2_74# FAX1_18/C Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M5864 gnd OAI21X1_4/A OAI21X1_4/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M5865 vdd BUFX2_19/Y OAI21X1_4/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M5866 OAI21X1_4/Y BUFX2_19/Y OAI21X1_4/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5867 OAI21X1_4/Y OR2X1_12/Y OAI21X1_4/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5868 OAI21X1_4/a_9_54# OAI21X1_4/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5869 OAI21X1_4/a_2_6# OR2X1_12/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5870 gnd out_mines[17] OAI22X1_50/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M5871 OAI22X1_50/a_2_6# out_mines[16] OAI22X1_50/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M5872 OAI22X1_50/Y OAI22X1_52/D OAI22X1_50/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5873 OAI22X1_50/Y OAI22X1_52/B OAI22X1_50/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M5874 OAI22X1_50/a_28_54# OAI22X1_52/D OAI22X1_50/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M5875 OAI22X1_50/a_9_54# out_mines[17] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5876 OAI22X1_50/a_2_6# OAI22X1_52/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5877 vdd out_mines[16] OAI22X1_50/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5878 gnd out_mines[19] OAI22X1_61/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M5879 OAI22X1_61/a_2_6# out_mines[18] OAI22X1_61/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M5880 OAI22X1_61/Y OAI22X1_63/D OAI22X1_61/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5881 OAI22X1_61/Y OAI22X1_63/B OAI22X1_61/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M5882 OAI22X1_61/a_28_54# OAI22X1_63/D OAI22X1_61/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M5883 OAI22X1_61/a_9_54# out_mines[19] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5884 OAI22X1_61/a_2_6# OAI22X1_63/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5885 vdd out_mines[18] OAI22X1_61/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5886 gnd out_mines[13] OAI22X1_72/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M5887 OAI22X1_72/a_2_6# out_mines[12] OAI22X1_72/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M5888 OAI22X1_72/Y OAI22X1_76/D OAI22X1_72/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5889 OAI22X1_72/Y OAI22X1_76/B OAI22X1_72/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M5890 OAI22X1_72/a_28_54# OAI22X1_76/D OAI22X1_72/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M5891 OAI22X1_72/a_9_54# out_mines[13] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5892 OAI22X1_72/a_2_6# OAI22X1_76/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5893 vdd out_mines[12] OAI22X1_72/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5894 gnd out_mines[15] OAI22X1_83/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M5895 OAI22X1_83/a_2_6# out_mines[14] OAI22X1_83/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M5896 OAI22X1_83/Y OAI22X1_87/D OAI22X1_83/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5897 OAI22X1_83/Y OAI22X1_87/B OAI22X1_83/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M5898 OAI22X1_83/a_28_54# OAI22X1_87/D OAI22X1_83/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M5899 OAI22X1_83/a_9_54# out_mines[15] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5900 OAI22X1_83/a_2_6# OAI22X1_87/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5901 vdd out_mines[14] OAI22X1_83/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5902 DFFNEGX1_2/a_76_6# BUFX2_17/Y DFFNEGX1_2/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M5903 gnd BUFX2_17/Y DFFNEGX1_2/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5904 DFFNEGX1_2/a_66_6# DFFNEGX1_2/a_2_6# DFFNEGX1_2/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5905 out_temp_index[1] DFFNEGX1_2/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5906 DFFNEGX1_2/a_23_6# BUFX2_17/Y DFFNEGX1_2/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M5907 DFFNEGX1_2/a_23_6# DFFNEGX1_2/a_2_6# DFFNEGX1_2/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M5908 gnd DFFNEGX1_2/a_34_4# DFFNEGX1_2/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5909 vdd DFFNEGX1_2/a_34_4# DFFNEGX1_2/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M5910 DFFNEGX1_2/a_61_74# DFFNEGX1_2/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5911 DFFNEGX1_2/a_34_4# DFFNEGX1_2/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5912 DFFNEGX1_2/a_34_4# DFFNEGX1_2/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M5913 vdd out_temp_index[1] DFFNEGX1_2/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M5914 gnd out_temp_index[1] DFFNEGX1_2/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5915 DFFNEGX1_2/a_61_6# DFFNEGX1_2/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5916 DFFNEGX1_2/a_76_84# DFFNEGX1_2/a_2_6# DFFNEGX1_2/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M5917 out_temp_index[1] DFFNEGX1_2/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5918 vdd BUFX2_17/Y DFFNEGX1_2/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M5919 DFFNEGX1_2/a_31_6# DFFNEGX1_2/a_2_6# DFFNEGX1_2/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5920 DFFNEGX1_2/a_66_6# BUFX2_17/Y DFFNEGX1_2/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5921 DFFNEGX1_2/a_17_74# OAI21X1_55/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5922 DFFNEGX1_2/a_31_74# BUFX2_17/Y DFFNEGX1_2/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5923 DFFNEGX1_2/a_17_6# OAI21X1_55/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M5924 gnd XOR2X1_7/A XOR2X1_7/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5925 XOR2X1_7/Y XOR2X1_7/a_2_6# XOR2X1_7/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M5926 XOR2X1_7/a_13_43# FAX1_5/YS gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5927 XOR2X1_7/a_18_54# XOR2X1_7/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M5928 XOR2X1_7/a_35_6# XOR2X1_7/A XOR2X1_7/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5929 XOR2X1_7/a_18_6# XOR2X1_7/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5930 vdd XOR2X1_7/A XOR2X1_7/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M5931 vdd FAX1_5/YS XOR2X1_7/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5932 XOR2X1_7/Y XOR2X1_7/A XOR2X1_7/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M5933 XOR2X1_7/a_35_54# XOR2X1_7/a_2_6# XOR2X1_7/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5934 XOR2X1_7/a_13_43# FAX1_5/YS vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5935 gnd FAX1_5/YS XOR2X1_7/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5936 gnd MUX2X1_8/A MUX2X1_8/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M5937 MUX2X1_8/a_17_50# NOR2X1_5/A vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M5938 MUX2X1_8/Y OR2X1_5/Y MUX2X1_8/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M5939 MUX2X1_8/a_30_54# MUX2X1_8/a_2_10# MUX2X1_8/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M5940 MUX2X1_8/a_17_10# NOR2X1_5/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5941 vdd OR2X1_5/Y MUX2X1_8/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5942 MUX2X1_8/a_30_10# OR2X1_5/Y MUX2X1_8/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M5943 gnd OR2X1_5/Y MUX2X1_8/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M5944 vdd MUX2X1_8/A MUX2X1_8/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5945 MUX2X1_8/Y MUX2X1_8/a_2_10# MUX2X1_8/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5946 INVX2_114/Y out_global_score[0] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5947 INVX2_114/Y out_global_score[0] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5948 INVX2_103/Y out_temp_cleared[10] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5949 INVX2_103/Y out_temp_cleared[10] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5950 OR2X1_5/A MUX2X1_0/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5951 OR2X1_5/A MUX2X1_0/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5952 NOR2X1_17/B in_mult[1] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5953 NOR2X1_17/B in_mult[1] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5954 INVX2_125/Y out_state_main[1] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5955 INVX2_125/Y out_state_main[1] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5956 HAX1_43/A MUX2X1_11/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5957 HAX1_43/A MUX2X1_11/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5958 NOR2X1_1/A MUX2X1_24/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5959 NOR2X1_1/A MUX2X1_24/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5960 FAX1_10/a_46_54# FAX1_10/A vdd vdd pfet w=40 l=2
+  ad=0.118n pd=46u as=0.12n ps=46u
M5961 gnd FAX1_10/A FAX1_10/a_2_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=26u as=100p ps=50u
M5962 gnd FAX1_10/A FAX1_10/a_84_6# Gnd nfet w=20 l=2
+  ad=55p pd=26u as=29.999998p ps=23u
M5963 FAX1_10/a_33_6# FAX1_10/B FAX1_10/a_25_6# Gnd nfet w=20 l=2
+  ad=29.999998p pd=23u as=59.999996p ps=26u
M5964 FAX1_10/a_79_6# FAX1_10/C FAX1_10/a_70_6# Gnd nfet w=20 l=2
+  ad=29.999998p pd=23u as=70p ps=27u
M5965 FAX1_10/a_46_6# FAX1_10/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=26u as=59.999996p ps=26u
M5966 FAX1_2/A FAX1_10/a_70_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0.13n ps=54u
M5967 FAX1_10/a_46_6# FAX1_10/C gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=26u as=59.999996p ps=26u
M5968 FAX1_10/a_79_46# FAX1_10/C FAX1_10/a_70_6# vdd pfet w=48 l=2
+  ad=72p pd=51u as=0.158n ps=55u
M5969 FAX1_9/C FAX1_10/a_25_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M5970 FAX1_10/a_2_54# FAX1_10/B vdd vdd pfet w=40 l=2
+  ad=0.12n pd=46u as=0.12n ps=46u
M5971 FAX1_10/a_25_6# FAX1_10/C FAX1_10/a_2_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=26u as=59.999996p ps=26u
M5972 gnd FAX1_10/A FAX1_10/a_33_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=26u as=29.999998p ps=23u
M5973 FAX1_10/a_70_6# FAX1_10/a_25_6# FAX1_10/a_46_54# vdd pfet w=36 l=2
+  ad=0.158n pd=55u as=0.108n ps=42u
M5974 FAX1_10/a_84_6# FAX1_10/B FAX1_10/a_79_6# Gnd nfet w=20 l=2
+  ad=29.999998p pd=23u as=29.999998p ps=23u
M5975 vdd FAX1_10/B FAX1_10/a_46_54# vdd pfet w=36 l=2
+  ad=0.108n pd=42u as=0.118n ps=46u
M5976 vdd FAX1_10/A FAX1_10/a_84_46# vdd pfet w=48 l=2
+  ad=0.13n pd=54u as=72p ps=51u
M5977 vdd FAX1_10/A FAX1_10/a_2_54# vdd pfet w=40 l=2
+  ad=0.12n pd=46u as=0.2n ps=90u
M5978 FAX1_2/A FAX1_10/a_70_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=55p ps=26u
M5979 FAX1_10/a_25_6# FAX1_10/C FAX1_10/a_2_54# vdd pfet w=40 l=2
+  ad=0.12n pd=46u as=0.12n ps=46u
M5980 gnd FAX1_10/B FAX1_10/a_46_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=26u as=59.999996p ps=26u
M5981 vdd FAX1_10/A FAX1_10/a_33_54# vdd pfet w=40 l=2
+  ad=0.12n pd=46u as=59.999996p ps=43u
M5982 FAX1_10/a_84_46# FAX1_10/B FAX1_10/a_79_46# vdd pfet w=48 l=2
+  ad=72p pd=51u as=72p ps=51u
M5983 FAX1_10/a_70_6# FAX1_10/a_25_6# FAX1_10/a_46_6# Gnd nfet w=20 l=2
+  ad=70p pd=27u as=59.999996p ps=26u
M5984 FAX1_10/a_46_54# FAX1_10/C vdd vdd pfet w=36 l=2
+  ad=0.108n pd=42u as=0.108n ps=42u
M5985 FAX1_9/C FAX1_10/a_25_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M5986 FAX1_10/a_2_6# FAX1_10/B gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=26u as=59.999996p ps=26u
M5987 FAX1_10/a_33_54# FAX1_10/B FAX1_10/a_25_6# vdd pfet w=40 l=2
+  ad=59.999996p pd=43u as=0.12n ps=46u
M5988 gnd XOR2X1_28/A XOR2X1_18/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M5989 XOR2X1_18/Y XOR2X1_18/a_2_6# XOR2X1_18/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M5990 XOR2X1_18/a_13_43# XOR2X1_19/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M5991 XOR2X1_18/a_18_54# XOR2X1_18/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M5992 XOR2X1_18/a_35_6# XOR2X1_28/A XOR2X1_18/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M5993 XOR2X1_18/a_18_6# XOR2X1_18/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M5994 vdd XOR2X1_28/A XOR2X1_18/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M5995 vdd XOR2X1_19/Y XOR2X1_18/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M5996 XOR2X1_18/Y XOR2X1_28/A XOR2X1_18/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M5997 XOR2X1_18/a_35_54# XOR2X1_18/a_2_6# XOR2X1_18/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M5998 XOR2X1_18/a_13_43# XOR2X1_19/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M5999 gnd XOR2X1_19/Y XOR2X1_18/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6000 gnd INVX2_40/Y XOR2X1_29/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6001 XOR2X1_29/Y XOR2X1_29/a_2_6# XOR2X1_29/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M6002 XOR2X1_29/a_13_43# XOR2X1_29/B gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6003 XOR2X1_29/a_18_54# XOR2X1_29/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M6004 XOR2X1_29/a_35_6# INVX2_40/Y XOR2X1_29/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6005 XOR2X1_29/a_18_6# XOR2X1_29/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6006 vdd INVX2_40/Y XOR2X1_29/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M6007 vdd XOR2X1_29/B XOR2X1_29/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6008 XOR2X1_29/Y INVX2_40/Y XOR2X1_29/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M6009 XOR2X1_29/a_35_54# XOR2X1_29/a_2_6# XOR2X1_29/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6010 XOR2X1_29/a_13_43# XOR2X1_29/B vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6011 gnd XOR2X1_29/B XOR2X1_29/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6012 NAND3X1_8/Y NAND3X1_9/A vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M6013 NAND3X1_8/a_9_6# NAND3X1_9/A gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M6014 NAND3X1_8/Y NOR2X1_63/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6015 NAND3X1_8/Y NOR2X1_63/Y NAND3X1_8/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M6016 vdd NOR2X1_66/A NAND3X1_8/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6017 NAND3X1_8/a_14_6# NOR2X1_66/A NAND3X1_8/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M6018 gnd INVX2_57/Y OAI21X1_104/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M6019 vdd NAND2X1_91/Y OAI21X1_104/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M6020 OAI21X1_104/Y NAND2X1_91/Y OAI21X1_104/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6021 OAI21X1_104/Y BUFX2_23/Y OAI21X1_104/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6022 OAI21X1_104/a_9_54# INVX2_57/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6023 OAI21X1_104/a_2_6# BUFX2_23/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6024 gnd OAI22X1_62/Y OAI21X1_137/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M6025 vdd out_temp_data_in[2] OAI21X1_137/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M6026 OAI21X1_137/Y out_temp_data_in[2] OAI21X1_137/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6027 OAI21X1_137/Y OAI22X1_61/Y OAI21X1_137/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6028 OAI21X1_137/a_9_54# OAI22X1_62/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6029 OAI21X1_137/a_2_6# OAI22X1_61/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6030 gnd out_temp_data_in[2] OAI21X1_115/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M6031 vdd OAI21X1_116/Y INVX2_43/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M6032 INVX2_43/A OAI21X1_116/Y OAI21X1_115/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6033 INVX2_43/A AOI22X1_59/Y OAI21X1_115/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6034 OAI21X1_115/a_9_54# out_temp_data_in[2] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6035 OAI21X1_115/a_2_6# AOI22X1_59/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6036 gnd OAI22X1_44/Y OAI21X1_126/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M6037 vdd INVX2_52/A AOI21X1_11/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M6038 AOI21X1_11/A INVX2_52/A OAI21X1_126/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6039 AOI21X1_11/A OAI22X1_43/Y OAI21X1_126/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6040 OAI21X1_126/a_9_54# OAI22X1_44/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6041 OAI21X1_126/a_2_6# OAI22X1_43/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6042 gnd INVX2_130/Y OAI21X1_159/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M6043 vdd NAND3X1_52/Y OAI21X1_159/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M6044 OAI21X1_159/Y NAND3X1_52/Y OAI21X1_159/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6045 OAI21X1_159/Y OAI21X1_160/Y OAI21X1_159/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6046 OAI21X1_159/a_9_54# INVX2_130/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6047 OAI21X1_159/a_2_6# OAI21X1_160/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6048 gnd AOI21X1_18/Y OAI21X1_148/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M6049 vdd XOR2X1_12/Y OAI21X1_148/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M6050 OAI21X1_148/Y XOR2X1_12/Y OAI21X1_148/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6051 OAI21X1_148/Y AOI21X1_17/Y OAI21X1_148/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6052 OAI21X1_148/a_9_54# AOI21X1_18/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6053 OAI21X1_148/a_2_6# AOI21X1_17/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6054 vdd in_clka BUFX2_2/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6055 gnd in_clka BUFX2_2/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M6056 BUFX2_2/Y BUFX2_2/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6057 BUFX2_2/Y BUFX2_2/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6058 OAI22X1_51/D INVX2_53/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M6059 NAND2X1_110/a_9_6# INVX2_53/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6060 vdd out_temp_data_in[0] OAI22X1_51/D vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6061 OAI22X1_51/D out_temp_data_in[0] NAND2X1_110/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6062 FAX1_0/a_46_54# FAX1_0/A vdd vdd pfet w=40 l=2
+  ad=0.452n pd=0.176m as=0 ps=0
M6063 gnd FAX1_0/A FAX1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M6064 gnd FAX1_0/A FAX1_0/a_84_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M6065 FAX1_0/a_33_6# in_incr[4] FAX1_0/a_25_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.12n ps=52u
M6066 FAX1_0/a_79_6# FAX1_0/C FAX1_0/a_70_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.14n ps=54u
M6067 FAX1_0/a_46_6# FAX1_0/A gnd Gnd nfet w=20 l=2
+  ad=0.24n pd=0.104m as=0 ps=0
M6068 FAX1_0/YS FAX1_0/a_70_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6069 FAX1_0/a_46_6# FAX1_0/C gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6070 FAX1_0/a_79_46# FAX1_0/C FAX1_0/a_70_6# vdd pfet w=48 l=2
+  ad=0.144n pd=0.102m as=0.317n ps=0.11m
M6071 FAX1_0/YC FAX1_0/a_25_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6072 FAX1_0/a_2_54# in_incr[4] vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M6073 FAX1_0/a_25_6# FAX1_0/C FAX1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6074 gnd FAX1_0/A FAX1_0/a_33_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6075 FAX1_0/a_70_6# FAX1_0/a_25_6# FAX1_0/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M6076 FAX1_0/a_84_6# in_incr[4] FAX1_0/a_79_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6077 vdd in_incr[4] FAX1_0/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M6078 vdd FAX1_0/A FAX1_0/a_84_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0.144n ps=0.102m
M6079 vdd FAX1_0/A FAX1_0/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6080 FAX1_0/YS FAX1_0/a_70_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M6081 FAX1_0/a_25_6# FAX1_0/C FAX1_0/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M6082 gnd in_incr[4] FAX1_0/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6083 vdd FAX1_0/A FAX1_0/a_33_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6084 FAX1_0/a_84_46# in_incr[4] FAX1_0/a_79_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0 ps=0
M6085 FAX1_0/a_70_6# FAX1_0/a_25_6# FAX1_0/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6086 FAX1_0/a_46_54# FAX1_0/C vdd vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M6087 FAX1_0/YC FAX1_0/a_25_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M6088 FAX1_0/a_2_6# in_incr[4] gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6089 FAX1_0/a_33_54# in_incr[4] FAX1_0/a_25_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6090 NOR2X1_124/B NOR2X1_125/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M6091 NAND2X1_132/a_9_6# NOR2X1_125/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6092 vdd INVX2_119/Y NOR2X1_124/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6093 NOR2X1_124/B INVX2_119/Y NAND2X1_132/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6094 OAI22X1_75/B INVX2_37/A vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M6095 NAND2X1_121/a_9_6# INVX2_37/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6096 vdd INVX2_251/Y OAI22X1_75/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6097 OAI22X1_75/B INVX2_251/Y NAND2X1_121/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6098 INVX2_2/Y out_temp_index[1] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6099 INVX2_2/Y out_temp_index[1] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6100 AOI21X1_2/a_2_54# out_gameover vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M6101 AOI21X1_2/a_12_6# AOI21X1_2/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6102 gnd AOI21X1_3/Y INVX2_218/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0.11n ps=52u
M6103 vdd AOI21X1_2/A AOI21X1_2/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6104 INVX2_218/A AOI21X1_3/Y AOI21X1_2/a_2_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6105 INVX2_218/A out_gameover AOI21X1_2/a_12_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6106 gnd NOR2X1_5/A XNOR2X1_10/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6107 MUX2X1_8/A NOR2X1_5/A XNOR2X1_10/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M6108 XNOR2X1_10/a_12_41# XOR2X1_9/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6109 XNOR2X1_10/a_18_54# XNOR2X1_10/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M6110 XNOR2X1_10/a_35_6# XNOR2X1_10/a_2_6# MUX2X1_8/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6111 XNOR2X1_10/a_18_6# XNOR2X1_10/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6112 vdd NOR2X1_5/A XNOR2X1_10/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M6113 vdd XOR2X1_9/Y XNOR2X1_10/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6114 MUX2X1_8/A XNOR2X1_10/a_2_6# XNOR2X1_10/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M6115 XNOR2X1_10/a_35_54# NOR2X1_5/A MUX2X1_8/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6116 XNOR2X1_10/a_12_41# XOR2X1_9/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6117 gnd XOR2X1_9/Y XNOR2X1_10/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6118 gnd out_temp_data_in[4] XNOR2X1_21/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6119 XNOR2X1_21/Y out_temp_data_in[4] XNOR2X1_21/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M6120 XNOR2X1_21/a_12_41# NOR2X1_33/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6121 XNOR2X1_21/a_18_54# XNOR2X1_21/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M6122 XNOR2X1_21/a_35_6# XNOR2X1_21/a_2_6# XNOR2X1_21/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6123 XNOR2X1_21/a_18_6# XNOR2X1_21/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6124 vdd out_temp_data_in[4] XNOR2X1_21/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M6125 vdd NOR2X1_33/Y XNOR2X1_21/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6126 XNOR2X1_21/Y XNOR2X1_21/a_2_6# XNOR2X1_21/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M6127 XNOR2X1_21/a_35_54# out_temp_data_in[4] XNOR2X1_21/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6128 XNOR2X1_21/a_12_41# NOR2X1_33/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6129 gnd NOR2X1_33/Y XNOR2X1_21/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6130 vdd BUFX2_21/A BUFX2_20/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6131 gnd BUFX2_21/A BUFX2_20/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M6132 BUFX2_20/Y BUFX2_20/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6133 BUFX2_20/Y BUFX2_20/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6134 NOR2X1_0/Y NOR2X1_0/A gnd Gnd nfet w=10 l=2
+  ad=29.999998p pd=16u as=50p ps=30u
M6135 NOR2X1_0/Y NOR2X1_0/B NOR2X1_0/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=59.999996p ps=43u
M6136 NOR2X1_0/a_9_54# NOR2X1_0/A vdd vdd pfet w=40 l=2
+  ad=59.999996p pd=43u as=0.2n ps=90u
M6137 gnd NOR2X1_0/B NOR2X1_0/Y Gnd nfet w=10 l=2
+  ad=50p pd=30u as=29.999998p ps=16u
M6138 AOI21X1_10/a_2_54# AOI22X1_60/Y vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M6139 AOI21X1_10/a_12_6# AOI22X1_61/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6140 gnd INVX2_32/A AOI21X1_9/C Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0.11n ps=52u
M6141 vdd AOI22X1_61/Y AOI21X1_10/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6142 AOI21X1_9/C INVX2_32/A AOI21X1_10/a_2_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6143 AOI21X1_9/C AOI22X1_60/Y AOI21X1_10/a_12_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6144 vdd out_global_score[17] HAX1_13/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M6145 HAX1_13/a_41_74# HAX1_13/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M6146 HAX1_13/a_9_6# out_global_score[17] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6147 HAX1_13/a_41_74# HAX1_13/B HAX1_13/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M6148 vdd out_global_score[17] HAX1_13/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6149 vdd HAX1_13/a_2_74# HAX1_12/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6150 HAX1_13/a_38_6# HAX1_13/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6151 HAX1_13/YS HAX1_13/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6152 HAX1_13/a_38_6# out_global_score[17] HAX1_13/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6153 HAX1_13/YS HAX1_13/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M6154 HAX1_13/a_2_74# HAX1_13/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6155 HAX1_13/a_2_74# HAX1_13/B HAX1_13/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6156 HAX1_13/a_49_54# HAX1_13/B HAX1_13/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6157 gnd HAX1_13/a_2_74# HAX1_12/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M6158 AOI21X1_21/a_2_54# out_display_done vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M6159 AOI21X1_21/a_12_6# in_data_in gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6160 gnd INVX2_122/A INVX2_133/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0.11n ps=52u
M6161 vdd in_data_in AOI21X1_21/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6162 INVX2_133/A INVX2_122/A AOI21X1_21/a_2_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6163 INVX2_133/A out_display_done AOI21X1_21/a_12_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6164 vdd HAX1_46/A HAX1_46/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M6165 HAX1_46/a_41_74# HAX1_46/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M6166 HAX1_46/a_9_6# HAX1_46/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6167 HAX1_46/a_41_74# HAX1_46/B HAX1_46/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M6168 vdd HAX1_46/A HAX1_46/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6169 vdd HAX1_46/a_2_74# HAX1_47/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6170 HAX1_46/a_38_6# HAX1_46/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6171 HAX1_46/YS HAX1_46/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6172 HAX1_46/a_38_6# HAX1_46/A HAX1_46/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6173 HAX1_46/YS HAX1_46/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M6174 HAX1_46/a_2_74# HAX1_46/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6175 HAX1_46/a_2_74# HAX1_46/B HAX1_46/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6176 HAX1_46/a_49_54# HAX1_46/B HAX1_46/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6177 gnd HAX1_46/a_2_74# HAX1_47/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M6178 vdd out_global_score[6] HAX1_24/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M6179 HAX1_24/a_41_74# HAX1_24/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M6180 HAX1_24/a_9_6# out_global_score[6] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6181 HAX1_24/a_41_74# HAX1_24/B HAX1_24/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M6182 vdd out_global_score[6] HAX1_24/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6183 vdd HAX1_24/a_2_74# HAX1_23/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6184 HAX1_24/a_38_6# HAX1_24/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6185 HAX1_24/YS HAX1_24/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6186 HAX1_24/a_38_6# out_global_score[6] HAX1_24/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6187 HAX1_24/YS HAX1_24/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M6188 HAX1_24/a_2_74# HAX1_24/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6189 HAX1_24/a_2_74# HAX1_24/B HAX1_24/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6190 HAX1_24/a_49_54# HAX1_24/B HAX1_24/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6191 gnd HAX1_24/a_2_74# HAX1_23/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M6192 vdd out_temp_mine_cnt[3] HAX1_35/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M6193 HAX1_35/a_41_74# HAX1_35/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M6194 HAX1_35/a_9_6# out_temp_mine_cnt[3] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6195 HAX1_35/a_41_74# HAX1_35/B HAX1_35/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M6196 vdd out_temp_mine_cnt[3] HAX1_35/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6197 vdd HAX1_35/a_2_74# XOR2X1_1/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6198 HAX1_35/a_38_6# HAX1_35/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6199 HAX1_35/YS HAX1_35/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6200 HAX1_35/a_38_6# out_temp_mine_cnt[3] HAX1_35/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6201 HAX1_35/YS HAX1_35/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M6202 HAX1_35/a_2_74# HAX1_35/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6203 HAX1_35/a_2_74# HAX1_35/B HAX1_35/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6204 HAX1_35/a_49_54# HAX1_35/B HAX1_35/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6205 gnd HAX1_35/a_2_74# XOR2X1_1/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M6206 gnd OAI21X1_5/A OAI21X1_5/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M6207 vdd OAI21X1_5/C OAI21X1_5/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M6208 OAI21X1_5/Y OAI21X1_5/C OAI21X1_5/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6209 OAI21X1_5/Y OAI21X1_9/B OAI21X1_5/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6210 OAI21X1_5/a_9_54# OAI21X1_5/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6211 OAI21X1_5/a_2_6# OAI21X1_9/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6212 gnd out_mines[23] OAI22X1_51/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M6213 OAI22X1_51/a_2_6# out_mines[22] OAI22X1_51/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M6214 OAI22X1_51/Y OAI22X1_51/D OAI22X1_51/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6215 OAI22X1_51/Y OAI22X1_51/B OAI22X1_51/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M6216 OAI22X1_51/a_28_54# OAI22X1_51/D OAI22X1_51/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M6217 OAI22X1_51/a_9_54# out_mines[23] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6218 OAI22X1_51/a_2_6# OAI22X1_51/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6219 vdd out_mines[22] OAI22X1_51/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6220 gnd INVX2_26/Y OAI22X1_40/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M6221 OAI22X1_40/a_2_6# out_temp_data_in[0] OAI22X1_40/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M6222 OAI22X1_40/Y OAI22X1_40/D OAI22X1_40/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6223 OAI22X1_40/Y INVX2_41/A OAI22X1_40/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M6224 OAI22X1_40/a_28_54# OAI22X1_40/D OAI22X1_40/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M6225 OAI22X1_40/a_9_54# INVX2_26/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6226 OAI22X1_40/a_2_6# INVX2_41/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6227 vdd out_temp_data_in[0] OAI22X1_40/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6228 gnd out_mines[19] OAI22X1_73/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M6229 OAI22X1_73/a_2_6# out_mines[18] OAI22X1_73/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M6230 OAI22X1_73/Y OAI22X1_75/D OAI22X1_73/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6231 OAI22X1_73/Y OAI22X1_75/B OAI22X1_73/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M6232 OAI22X1_73/a_28_54# OAI22X1_75/D OAI22X1_73/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M6233 OAI22X1_73/a_9_54# out_mines[19] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6234 OAI22X1_73/a_2_6# OAI22X1_75/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6235 vdd out_mines[18] OAI22X1_73/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6236 gnd out_mines[13] OAI22X1_84/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M6237 OAI22X1_84/a_2_6# out_mines[12] OAI22X1_84/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M6238 OAI22X1_84/Y OAI22X1_88/D OAI22X1_84/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6239 OAI22X1_84/Y OAI22X1_88/B OAI22X1_84/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M6240 OAI22X1_84/a_28_54# OAI22X1_88/D OAI22X1_84/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M6241 OAI22X1_84/a_9_54# out_mines[13] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6242 OAI22X1_84/a_2_6# OAI22X1_88/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6243 vdd out_mines[12] OAI22X1_84/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6244 gnd out_mines[17] OAI22X1_62/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M6245 OAI22X1_62/a_2_6# out_mines[16] OAI22X1_62/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M6246 OAI22X1_62/Y OAI22X1_64/D OAI22X1_62/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6247 OAI22X1_62/Y OAI22X1_64/B OAI22X1_62/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M6248 OAI22X1_62/a_28_54# OAI22X1_64/D OAI22X1_62/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M6249 OAI22X1_62/a_9_54# out_mines[17] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6250 OAI22X1_62/a_2_6# OAI22X1_64/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6251 vdd out_mines[16] OAI22X1_62/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6252 DFFNEGX1_3/a_76_6# BUFX2_17/Y DFFNEGX1_3/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M6253 gnd BUFX2_17/Y DFFNEGX1_3/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6254 DFFNEGX1_3/a_66_6# DFFNEGX1_3/a_2_6# DFFNEGX1_3/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M6255 out_temp_index[2] DFFNEGX1_3/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6256 DFFNEGX1_3/a_23_6# BUFX2_17/Y DFFNEGX1_3/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M6257 DFFNEGX1_3/a_23_6# DFFNEGX1_3/a_2_6# DFFNEGX1_3/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M6258 gnd DFFNEGX1_3/a_34_4# DFFNEGX1_3/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M6259 vdd DFFNEGX1_3/a_34_4# DFFNEGX1_3/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M6260 DFFNEGX1_3/a_61_74# DFFNEGX1_3/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6261 DFFNEGX1_3/a_34_4# DFFNEGX1_3/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6262 DFFNEGX1_3/a_34_4# DFFNEGX1_3/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M6263 vdd out_temp_index[2] DFFNEGX1_3/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M6264 gnd out_temp_index[2] DFFNEGX1_3/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6265 DFFNEGX1_3/a_61_6# DFFNEGX1_3/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6266 DFFNEGX1_3/a_76_84# DFFNEGX1_3/a_2_6# DFFNEGX1_3/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M6267 out_temp_index[2] DFFNEGX1_3/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6268 vdd BUFX2_17/Y DFFNEGX1_3/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M6269 DFFNEGX1_3/a_31_6# DFFNEGX1_3/a_2_6# DFFNEGX1_3/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6270 DFFNEGX1_3/a_66_6# BUFX2_17/Y DFFNEGX1_3/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6271 DFFNEGX1_3/a_17_74# INVX2_245/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6272 DFFNEGX1_3/a_31_74# BUFX2_17/Y DFFNEGX1_3/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6273 DFFNEGX1_3/a_17_6# INVX2_245/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6274 gnd XOR2X1_8/A XOR2X1_8/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6275 XOR2X1_8/Y XOR2X1_8/a_2_6# XOR2X1_8/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M6276 XOR2X1_8/a_13_43# FAX1_6/YS gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6277 XOR2X1_8/a_18_54# XOR2X1_8/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M6278 XOR2X1_8/a_35_6# XOR2X1_8/A XOR2X1_8/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6279 XOR2X1_8/a_18_6# XOR2X1_8/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6280 vdd XOR2X1_8/A XOR2X1_8/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M6281 vdd FAX1_6/YS XOR2X1_8/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6282 XOR2X1_8/Y XOR2X1_8/A XOR2X1_8/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M6283 XOR2X1_8/a_35_54# XOR2X1_8/a_2_6# XOR2X1_8/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6284 XOR2X1_8/a_13_43# FAX1_6/YS vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6285 gnd FAX1_6/YS XOR2X1_8/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6286 gnd MUX2X1_9/A MUX2X1_9/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M6287 MUX2X1_9/a_17_50# XOR2X1_9/Y vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M6288 MUX2X1_9/Y OR2X1_5/Y MUX2X1_9/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M6289 MUX2X1_9/a_30_54# MUX2X1_9/a_2_10# MUX2X1_9/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M6290 MUX2X1_9/a_17_10# XOR2X1_9/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6291 vdd OR2X1_5/Y MUX2X1_9/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6292 MUX2X1_9/a_30_10# OR2X1_5/Y MUX2X1_9/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M6293 gnd OR2X1_5/Y MUX2X1_9/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M6294 vdd MUX2X1_9/A MUX2X1_9/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6295 MUX2X1_9/Y MUX2X1_9/a_2_10# MUX2X1_9/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6296 INVX2_104/Y out_temp_cleared[9] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6297 INVX2_104/Y out_temp_cleared[9] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6298 MUX2X1_29/A FAX1_3/YS gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6299 MUX2X1_29/A FAX1_3/YS vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6300 OR2X1_16/A out_alu_done gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6301 OR2X1_16/A out_alu_done vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6302 INVX2_126/Y INVX2_126/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6303 INVX2_126/Y INVX2_126/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6304 MUX2X1_17/B XNOR2X1_7/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6305 MUX2X1_17/B XNOR2X1_7/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6306 HAX1_39/A MUX2X1_1/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6307 HAX1_39/A MUX2X1_1/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6308 FAX1_11/a_46_54# FAX1_11/A vdd vdd pfet w=40 l=2
+  ad=0.452n pd=0.176m as=0 ps=0
M6309 gnd FAX1_11/A FAX1_11/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M6310 gnd FAX1_11/A FAX1_11/a_84_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M6311 FAX1_11/a_33_6# FAX1_11/B FAX1_11/a_25_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.12n ps=52u
M6312 FAX1_11/a_79_6# FAX1_11/C FAX1_11/a_70_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.14n ps=54u
M6313 FAX1_11/a_46_6# FAX1_11/A gnd Gnd nfet w=20 l=2
+  ad=0.24n pd=0.104m as=0 ps=0
M6314 FAX1_5/A FAX1_11/a_70_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6315 FAX1_11/a_46_6# FAX1_11/C gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6316 FAX1_11/a_79_46# FAX1_11/C FAX1_11/a_70_6# vdd pfet w=48 l=2
+  ad=0.144n pd=0.102m as=0.317n ps=0.11m
M6317 FAX1_4/B FAX1_11/a_25_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6318 FAX1_11/a_2_54# FAX1_11/B vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M6319 FAX1_11/a_25_6# FAX1_11/C FAX1_11/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6320 gnd FAX1_11/A FAX1_11/a_33_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6321 FAX1_11/a_70_6# FAX1_11/a_25_6# FAX1_11/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M6322 FAX1_11/a_84_6# FAX1_11/B FAX1_11/a_79_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6323 vdd FAX1_11/B FAX1_11/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M6324 vdd FAX1_11/A FAX1_11/a_84_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0.144n ps=0.102m
M6325 vdd FAX1_11/A FAX1_11/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6326 FAX1_5/A FAX1_11/a_70_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M6327 FAX1_11/a_25_6# FAX1_11/C FAX1_11/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M6328 gnd FAX1_11/B FAX1_11/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6329 vdd FAX1_11/A FAX1_11/a_33_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6330 FAX1_11/a_84_46# FAX1_11/B FAX1_11/a_79_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0 ps=0
M6331 FAX1_11/a_70_6# FAX1_11/a_25_6# FAX1_11/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6332 FAX1_11/a_46_54# FAX1_11/C vdd vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M6333 FAX1_4/B FAX1_11/a_25_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M6334 FAX1_11/a_2_6# FAX1_11/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6335 FAX1_11/a_33_54# FAX1_11/B FAX1_11/a_25_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6336 gnd INVX2_40/Y XOR2X1_19/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6337 XOR2X1_19/Y XOR2X1_19/a_2_6# XOR2X1_19/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M6338 XOR2X1_19/a_13_43# XOR2X1_25/B gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6339 XOR2X1_19/a_18_54# XOR2X1_19/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M6340 XOR2X1_19/a_35_6# INVX2_40/Y XOR2X1_19/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6341 XOR2X1_19/a_18_6# XOR2X1_19/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6342 vdd INVX2_40/Y XOR2X1_19/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M6343 vdd XOR2X1_25/B XOR2X1_19/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6344 XOR2X1_19/Y INVX2_40/Y XOR2X1_19/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M6345 XOR2X1_19/a_35_54# XOR2X1_19/a_2_6# XOR2X1_19/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6346 XOR2X1_19/a_13_43# XOR2X1_25/B vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6347 gnd XOR2X1_25/B XOR2X1_19/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6348 OR2X1_12/B NAND3X1_9/A vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M6349 NAND3X1_9/a_9_6# NAND3X1_9/A gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M6350 OR2X1_12/B NOR2X1_65/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6351 OR2X1_12/B NOR2X1_65/Y NAND3X1_9/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M6352 vdd NOR2X1_66/A OR2X1_12/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6353 NAND3X1_9/a_14_6# NOR2X1_66/A NAND3X1_9/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M6354 gnd OAI22X1_46/Y OAI21X1_127/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M6355 vdd INVX2_52/Y AOI21X1_12/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M6356 AOI21X1_12/B INVX2_52/Y OAI21X1_127/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6357 AOI21X1_12/B OAI22X1_45/Y OAI21X1_127/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6358 OAI21X1_127/a_9_54# OAI22X1_46/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6359 OAI21X1_127/a_2_6# OAI22X1_45/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6360 gnd INVX2_56/Y OAI21X1_105/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M6361 vdd NAND2X1_92/Y OAI21X1_105/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M6362 OAI21X1_105/Y NAND2X1_92/Y OAI21X1_105/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6363 OAI21X1_105/Y BUFX2_23/Y OAI21X1_105/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6364 OAI21X1_105/a_9_54# INVX2_56/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6365 OAI21X1_105/a_2_6# BUFX2_23/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6366 gnd NOR2X1_109/Y OAI21X1_116/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M6367 vdd out_temp_data_in[2] OAI21X1_116/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M6368 OAI21X1_116/Y out_temp_data_in[2] OAI21X1_116/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6369 OAI21X1_116/Y OAI22X1_40/Y OAI21X1_116/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6370 OAI21X1_116/a_9_54# NOR2X1_109/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6371 OAI21X1_116/a_2_6# OAI22X1_40/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6372 gnd OAI22X1_64/Y OAI21X1_138/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M6373 vdd OAI21X1_1/B OAI21X1_138/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M6374 OAI21X1_138/Y OAI21X1_1/B OAI21X1_138/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6375 OAI21X1_138/Y OAI22X1_63/Y OAI21X1_138/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6376 OAI21X1_138/a_9_54# OAI22X1_64/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6377 OAI21X1_138/a_2_6# OAI22X1_63/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6378 gnd OAI22X1_78/Y OAI21X1_149/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M6379 vdd INVX2_35/Y AOI21X1_17/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M6380 AOI21X1_17/B INVX2_35/Y OAI21X1_149/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6381 AOI21X1_17/B OAI22X1_77/Y OAI21X1_149/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6382 OAI21X1_149/a_9_54# OAI22X1_78/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6383 OAI21X1_149/a_2_6# OAI22X1_77/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6384 vdd in_restart BUFX2_3/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6385 gnd in_restart BUFX2_3/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M6386 BUFX2_3/Y BUFX2_3/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6387 BUFX2_3/Y BUFX2_3/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6388 OAI21X1_111/C in_data[4] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M6389 NAND2X1_100/a_9_6# in_data[4] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6390 vdd NOR2X1_107/Y OAI21X1_111/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6391 OAI21X1_111/C NOR2X1_107/Y NAND2X1_100/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6392 FAX1_1/a_46_54# FAX1_1/A vdd vdd pfet w=40 l=2
+  ad=0.452n pd=0.176m as=0 ps=0
M6393 gnd FAX1_1/A FAX1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M6394 gnd FAX1_1/A FAX1_1/a_84_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M6395 FAX1_1/a_33_6# in_incr[3] FAX1_1/a_25_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.12n ps=52u
M6396 FAX1_1/a_79_6# FAX1_1/C FAX1_1/a_70_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.14n ps=54u
M6397 FAX1_1/a_46_6# FAX1_1/A gnd Gnd nfet w=20 l=2
+  ad=0.24n pd=0.104m as=0 ps=0
M6398 FAX1_1/YS FAX1_1/a_70_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6399 FAX1_1/a_46_6# FAX1_1/C gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6400 FAX1_1/a_79_46# FAX1_1/C FAX1_1/a_70_6# vdd pfet w=48 l=2
+  ad=0.144n pd=0.102m as=0.317n ps=0.11m
M6401 FAX1_0/C FAX1_1/a_25_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6402 FAX1_1/a_2_54# in_incr[3] vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M6403 FAX1_1/a_25_6# FAX1_1/C FAX1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6404 gnd FAX1_1/A FAX1_1/a_33_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6405 FAX1_1/a_70_6# FAX1_1/a_25_6# FAX1_1/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M6406 FAX1_1/a_84_6# in_incr[3] FAX1_1/a_79_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6407 vdd in_incr[3] FAX1_1/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M6408 vdd FAX1_1/A FAX1_1/a_84_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0.144n ps=0.102m
M6409 vdd FAX1_1/A FAX1_1/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6410 FAX1_1/YS FAX1_1/a_70_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M6411 FAX1_1/a_25_6# FAX1_1/C FAX1_1/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M6412 gnd in_incr[3] FAX1_1/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6413 vdd FAX1_1/A FAX1_1/a_33_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6414 FAX1_1/a_84_46# in_incr[3] FAX1_1/a_79_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0 ps=0
M6415 FAX1_1/a_70_6# FAX1_1/a_25_6# FAX1_1/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6416 FAX1_1/a_46_54# FAX1_1/C vdd vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M6417 FAX1_0/C FAX1_1/a_25_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M6418 FAX1_1/a_2_6# in_incr[3] gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6419 FAX1_1/a_33_54# in_incr[3] FAX1_1/a_25_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6420 OAI22X1_76/D out_temp_data_in[0] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M6421 NAND2X1_122/a_9_6# out_temp_data_in[0] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6422 vdd INVX2_37/Y OAI22X1_76/D vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6423 OAI22X1_76/D INVX2_37/Y NAND2X1_122/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6424 OAI22X1_51/B INVX2_53/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M6425 NAND2X1_111/a_9_6# INVX2_53/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6426 vdd INVX2_251/Y OAI22X1_51/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6427 OAI22X1_51/B INVX2_251/Y NAND2X1_111/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6428 INVX2_3/Y out_temp_index[2] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6429 INVX2_3/Y out_temp_index[2] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6430 AOI21X1_3/a_2_54# NOR2X1_79/Y vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M6431 AOI21X1_3/a_12_6# AOI21X1_3/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6432 gnd OR2X1_11/A AOI21X1_3/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0.11n ps=52u
M6433 vdd AOI21X1_3/A AOI21X1_3/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6434 AOI21X1_3/Y OR2X1_11/A AOI21X1_3/a_2_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6435 AOI21X1_3/Y NOR2X1_79/Y AOI21X1_3/a_12_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6436 gnd MUX2X1_3/Y XNOR2X1_11/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6437 MUX2X1_7/A MUX2X1_3/Y XNOR2X1_11/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M6438 XNOR2X1_11/a_12_41# NOR2X1_5/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6439 XNOR2X1_11/a_18_54# XNOR2X1_11/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M6440 XNOR2X1_11/a_35_6# XNOR2X1_11/a_2_6# MUX2X1_7/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6441 XNOR2X1_11/a_18_6# XNOR2X1_11/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6442 vdd MUX2X1_3/Y XNOR2X1_11/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M6443 vdd NOR2X1_5/Y XNOR2X1_11/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6444 MUX2X1_7/A XNOR2X1_11/a_2_6# XNOR2X1_11/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M6445 XNOR2X1_11/a_35_54# MUX2X1_3/Y MUX2X1_7/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6446 XNOR2X1_11/a_12_41# NOR2X1_5/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6447 gnd NOR2X1_5/Y XNOR2X1_11/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6448 gnd out_temp_mine_cnt[0] XNOR2X1_22/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6449 XNOR2X1_22/Y out_temp_mine_cnt[0] XNOR2X1_22/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M6450 XNOR2X1_22/a_12_41# in_n_mines[0] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6451 XNOR2X1_22/a_18_54# XNOR2X1_22/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M6452 XNOR2X1_22/a_35_6# XNOR2X1_22/a_2_6# XNOR2X1_22/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6453 XNOR2X1_22/a_18_6# XNOR2X1_22/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6454 vdd out_temp_mine_cnt[0] XNOR2X1_22/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M6455 vdd in_n_mines[0] XNOR2X1_22/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6456 XNOR2X1_22/Y XNOR2X1_22/a_2_6# XNOR2X1_22/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M6457 XNOR2X1_22/a_35_54# out_temp_mine_cnt[0] XNOR2X1_22/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6458 XNOR2X1_22/a_12_41# in_n_mines[0] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6459 gnd in_n_mines[0] XNOR2X1_22/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6460 vdd BUFX2_9/A BUFX2_10/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6461 gnd BUFX2_9/A BUFX2_10/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M6462 BUFX2_10/Y BUFX2_10/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6463 BUFX2_10/Y BUFX2_10/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6464 vdd BUFX2_21/A BUFX2_21/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6465 gnd BUFX2_21/A BUFX2_21/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M6466 BUFX2_21/Y BUFX2_21/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6467 BUFX2_21/Y BUFX2_21/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6468 NOR2X1_1/Y NOR2X1_1/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M6469 NOR2X1_1/Y FAX1_3/YS NOR2X1_1/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M6470 NOR2X1_1/a_9_54# NOR2X1_1/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6471 gnd FAX1_3/YS NOR2X1_1/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6472 vdd out_global_score[16] HAX1_14/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M6473 HAX1_14/a_41_74# HAX1_14/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M6474 HAX1_14/a_9_6# out_global_score[16] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6475 HAX1_14/a_41_74# HAX1_14/B HAX1_14/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M6476 vdd out_global_score[16] HAX1_14/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6477 vdd HAX1_14/a_2_74# HAX1_13/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6478 HAX1_14/a_38_6# HAX1_14/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6479 HAX1_14/YS HAX1_14/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6480 HAX1_14/a_38_6# out_global_score[16] HAX1_14/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6481 HAX1_14/YS HAX1_14/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M6482 HAX1_14/a_2_74# HAX1_14/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6483 HAX1_14/a_2_74# HAX1_14/B HAX1_14/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6484 HAX1_14/a_49_54# HAX1_14/B HAX1_14/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6485 gnd HAX1_14/a_2_74# HAX1_13/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M6486 AOI21X1_22/a_2_54# NOR2X1_117/Y vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M6487 AOI21X1_22/a_12_6# AND2X2_18/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6488 gnd INVX2_124/Y AOI21X1_22/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0.11n ps=52u
M6489 vdd AND2X2_18/Y AOI21X1_22/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6490 AOI21X1_22/Y INVX2_124/Y AOI21X1_22/a_2_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6491 AOI21X1_22/Y NOR2X1_117/Y AOI21X1_22/a_12_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6492 AOI21X1_11/a_2_54# AOI21X1_11/B vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M6493 AOI21X1_11/a_12_6# AOI21X1_11/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6494 gnd INVX2_51/A AOI21X1_11/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0.11n ps=52u
M6495 vdd AOI21X1_11/A AOI21X1_11/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6496 AOI21X1_11/Y INVX2_51/A AOI21X1_11/a_2_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6497 AOI21X1_11/Y AOI21X1_11/B AOI21X1_11/a_12_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6498 vdd HAX1_47/A HAX1_47/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M6499 HAX1_47/a_41_74# HAX1_47/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M6500 HAX1_47/a_9_6# HAX1_47/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6501 HAX1_47/a_41_74# HAX1_47/B HAX1_47/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M6502 vdd HAX1_47/A HAX1_47/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6503 vdd HAX1_47/a_2_74# OR2X1_1/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6504 HAX1_47/a_38_6# HAX1_47/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6505 HAX1_47/YS HAX1_47/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6506 HAX1_47/a_38_6# HAX1_47/A HAX1_47/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6507 HAX1_47/YS HAX1_47/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M6508 HAX1_47/a_2_74# HAX1_47/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6509 HAX1_47/a_2_74# HAX1_47/B HAX1_47/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6510 HAX1_47/a_49_54# HAX1_47/B HAX1_47/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6511 gnd HAX1_47/a_2_74# OR2X1_1/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M6512 vdd out_global_score[5] HAX1_25/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M6513 HAX1_25/a_41_74# HAX1_25/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M6514 HAX1_25/a_9_6# out_global_score[5] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6515 HAX1_25/a_41_74# HAX1_25/B HAX1_25/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M6516 vdd out_global_score[5] HAX1_25/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6517 vdd HAX1_25/a_2_74# HAX1_24/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6518 HAX1_25/a_38_6# HAX1_25/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6519 HAX1_25/YS HAX1_25/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6520 HAX1_25/a_38_6# out_global_score[5] HAX1_25/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6521 HAX1_25/YS HAX1_25/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M6522 HAX1_25/a_2_74# HAX1_25/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6523 HAX1_25/a_2_74# HAX1_25/B HAX1_25/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6524 HAX1_25/a_49_54# HAX1_25/B HAX1_25/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6525 gnd HAX1_25/a_2_74# HAX1_24/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M6526 vdd out_temp_mine_cnt[2] HAX1_36/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M6527 HAX1_36/a_41_74# HAX1_36/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M6528 HAX1_36/a_9_6# out_temp_mine_cnt[2] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6529 HAX1_36/a_41_74# HAX1_36/B HAX1_36/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M6530 vdd out_temp_mine_cnt[2] HAX1_36/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6531 vdd HAX1_36/a_2_74# HAX1_35/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6532 HAX1_36/a_38_6# HAX1_36/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6533 HAX1_36/YS HAX1_36/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6534 HAX1_36/a_38_6# out_temp_mine_cnt[2] HAX1_36/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6535 HAX1_36/YS HAX1_36/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M6536 HAX1_36/a_2_74# HAX1_36/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6537 HAX1_36/a_2_74# HAX1_36/B HAX1_36/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6538 HAX1_36/a_49_54# HAX1_36/B HAX1_36/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6539 gnd HAX1_36/a_2_74# HAX1_35/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M6540 gnd OAI21X1_6/A OAI21X1_6/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M6541 vdd BUFX2_19/Y OAI21X1_6/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M6542 OAI21X1_6/Y BUFX2_19/Y OAI21X1_6/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6543 OAI21X1_6/Y OAI21X1_8/A OAI21X1_6/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6544 OAI21X1_6/a_9_54# OAI21X1_6/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6545 OAI21X1_6/a_2_6# OAI21X1_8/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6546 gnd out_mines[21] OAI22X1_52/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M6547 OAI22X1_52/a_2_6# out_mines[20] OAI22X1_52/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M6548 OAI22X1_52/Y OAI22X1_52/D OAI22X1_52/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6549 OAI22X1_52/Y OAI22X1_52/B OAI22X1_52/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M6550 OAI22X1_52/a_28_54# OAI22X1_52/D OAI22X1_52/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M6551 OAI22X1_52/a_9_54# out_mines[21] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6552 OAI22X1_52/a_2_6# OAI22X1_52/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6553 vdd out_mines[20] OAI22X1_52/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6554 gnd out_mines[3] OAI22X1_41/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M6555 OAI22X1_41/a_2_6# out_mines[2] OAI22X1_41/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M6556 OAI22X1_41/Y OAI22X1_51/D OAI22X1_41/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6557 OAI22X1_41/Y OAI22X1_51/B OAI22X1_41/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M6558 OAI22X1_41/a_28_54# OAI22X1_51/D OAI22X1_41/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M6559 OAI22X1_41/a_9_54# out_mines[3] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6560 OAI22X1_41/a_2_6# OAI22X1_51/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6561 vdd out_mines[2] OAI22X1_41/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6562 gnd INVX2_50/Y OAI22X1_30/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M6563 OAI22X1_30/a_2_6# INVX2_40/A XNOR2X1_26/B Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M6564 XNOR2X1_26/B XOR2X1_22/Y OAI22X1_30/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6565 XNOR2X1_26/B XOR2X1_29/B OAI22X1_30/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M6566 OAI22X1_30/a_28_54# XOR2X1_22/Y XNOR2X1_26/B vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M6567 OAI22X1_30/a_9_54# INVX2_50/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6568 OAI22X1_30/a_2_6# XOR2X1_29/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6569 vdd INVX2_40/A OAI22X1_30/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6570 gnd out_mines[17] OAI22X1_74/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M6571 OAI22X1_74/a_2_6# out_mines[16] OAI22X1_74/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M6572 OAI22X1_74/Y OAI22X1_76/D OAI22X1_74/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6573 OAI22X1_74/Y OAI22X1_76/B OAI22X1_74/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M6574 OAI22X1_74/a_28_54# OAI22X1_76/D OAI22X1_74/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M6575 OAI22X1_74/a_9_54# out_mines[17] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6576 OAI22X1_74/a_2_6# OAI22X1_76/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6577 vdd out_mines[16] OAI22X1_74/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6578 gnd out_mines[19] OAI22X1_85/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M6579 OAI22X1_85/a_2_6# out_mines[18] OAI22X1_85/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M6580 OAI22X1_85/Y OAI22X1_87/D OAI22X1_85/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6581 OAI22X1_85/Y OAI22X1_87/B OAI22X1_85/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M6582 OAI22X1_85/a_28_54# OAI22X1_87/D OAI22X1_85/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M6583 OAI22X1_85/a_9_54# out_mines[19] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6584 OAI22X1_85/a_2_6# OAI22X1_87/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6585 vdd out_mines[18] OAI22X1_85/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6586 gnd out_mines[23] OAI22X1_63/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M6587 OAI22X1_63/a_2_6# out_mines[22] OAI22X1_63/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M6588 OAI22X1_63/Y OAI22X1_63/D OAI22X1_63/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6589 OAI22X1_63/Y OAI22X1_63/B OAI22X1_63/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M6590 OAI22X1_63/a_28_54# OAI22X1_63/D OAI22X1_63/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M6591 OAI22X1_63/a_9_54# out_mines[23] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6592 OAI22X1_63/a_2_6# OAI22X1_63/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6593 vdd out_mines[22] OAI22X1_63/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6594 DFFNEGX1_4/a_76_6# BUFX2_17/Y DFFNEGX1_4/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M6595 gnd BUFX2_17/Y DFFNEGX1_4/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6596 DFFNEGX1_4/a_66_6# DFFNEGX1_4/a_2_6# DFFNEGX1_4/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M6597 out_temp_index[3] DFFNEGX1_4/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6598 DFFNEGX1_4/a_23_6# BUFX2_17/Y DFFNEGX1_4/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M6599 DFFNEGX1_4/a_23_6# DFFNEGX1_4/a_2_6# DFFNEGX1_4/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M6600 gnd DFFNEGX1_4/a_34_4# DFFNEGX1_4/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M6601 vdd DFFNEGX1_4/a_34_4# DFFNEGX1_4/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M6602 DFFNEGX1_4/a_61_74# DFFNEGX1_4/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6603 DFFNEGX1_4/a_34_4# DFFNEGX1_4/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6604 DFFNEGX1_4/a_34_4# DFFNEGX1_4/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M6605 vdd out_temp_index[3] DFFNEGX1_4/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M6606 gnd out_temp_index[3] DFFNEGX1_4/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6607 DFFNEGX1_4/a_61_6# DFFNEGX1_4/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6608 DFFNEGX1_4/a_76_84# DFFNEGX1_4/a_2_6# DFFNEGX1_4/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M6609 out_temp_index[3] DFFNEGX1_4/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6610 vdd BUFX2_17/Y DFFNEGX1_4/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M6611 DFFNEGX1_4/a_31_6# DFFNEGX1_4/a_2_6# DFFNEGX1_4/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6612 DFFNEGX1_4/a_66_6# BUFX2_17/Y DFFNEGX1_4/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6613 DFFNEGX1_4/a_17_74# OAI21X1_54/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6614 DFFNEGX1_4/a_31_74# BUFX2_17/Y DFFNEGX1_4/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6615 DFFNEGX1_4/a_17_6# OAI21X1_54/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6616 gnd FAX1_0/YC XOR2X1_9/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6617 XOR2X1_9/Y XOR2X1_9/a_2_6# XOR2X1_9/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M6618 XOR2X1_9/a_13_43# FAX1_7/YS gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6619 XOR2X1_9/a_18_54# XOR2X1_9/a_13_43# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M6620 XOR2X1_9/a_35_6# FAX1_0/YC XOR2X1_9/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6621 XOR2X1_9/a_18_6# XOR2X1_9/a_13_43# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6622 vdd FAX1_0/YC XOR2X1_9/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M6623 vdd FAX1_7/YS XOR2X1_9/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6624 XOR2X1_9/Y FAX1_0/YC XOR2X1_9/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M6625 XOR2X1_9/a_35_54# XOR2X1_9/a_2_6# XOR2X1_9/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6626 XOR2X1_9/a_13_43# FAX1_7/YS vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6627 gnd FAX1_7/YS XOR2X1_9/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6628 OAI22X1_1/B out_temp_cleared[8] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6629 OAI22X1_1/B out_temp_cleared[8] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6630 NOR2X1_22/B in_mult[2] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6631 NOR2X1_22/B in_mult[2] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6632 OR2X1_15/B INVX2_127/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6633 OR2X1_15/B INVX2_127/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6634 INVX2_116/Y out_state_main[0] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6635 INVX2_116/Y out_state_main[0] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6636 HAX1_38/A MUX2X1_2/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6637 HAX1_38/A MUX2X1_2/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6638 FAX1_12/a_46_54# FAX1_12/A vdd vdd pfet w=40 l=2
+  ad=0.452n pd=0.176m as=0 ps=0
M6639 gnd FAX1_12/A FAX1_12/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M6640 gnd FAX1_12/A FAX1_12/a_84_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M6641 FAX1_12/a_33_6# FAX1_12/B FAX1_12/a_25_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.12n ps=52u
M6642 FAX1_12/a_79_6# FAX1_12/C FAX1_12/a_70_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.14n ps=54u
M6643 FAX1_12/a_46_6# FAX1_12/A gnd Gnd nfet w=20 l=2
+  ad=0.24n pd=0.104m as=0 ps=0
M6644 FAX1_6/B FAX1_12/a_70_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6645 FAX1_12/a_46_6# FAX1_12/C gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6646 FAX1_12/a_79_46# FAX1_12/C FAX1_12/a_70_6# vdd pfet w=48 l=2
+  ad=0.144n pd=0.102m as=0.317n ps=0.11m
M6647 FAX1_5/B FAX1_12/a_25_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6648 FAX1_12/a_2_54# FAX1_12/B vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M6649 FAX1_12/a_25_6# FAX1_12/C FAX1_12/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6650 gnd FAX1_12/A FAX1_12/a_33_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6651 FAX1_12/a_70_6# FAX1_12/a_25_6# FAX1_12/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M6652 FAX1_12/a_84_6# FAX1_12/B FAX1_12/a_79_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6653 vdd FAX1_12/B FAX1_12/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M6654 vdd FAX1_12/A FAX1_12/a_84_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0.144n ps=0.102m
M6655 vdd FAX1_12/A FAX1_12/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6656 FAX1_6/B FAX1_12/a_70_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M6657 FAX1_12/a_25_6# FAX1_12/C FAX1_12/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M6658 gnd FAX1_12/B FAX1_12/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6659 vdd FAX1_12/A FAX1_12/a_33_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6660 FAX1_12/a_84_46# FAX1_12/B FAX1_12/a_79_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0 ps=0
M6661 FAX1_12/a_70_6# FAX1_12/a_25_6# FAX1_12/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6662 FAX1_12/a_46_54# FAX1_12/C vdd vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M6663 FAX1_5/B FAX1_12/a_25_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M6664 FAX1_12/a_2_6# FAX1_12/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6665 FAX1_12/a_33_54# FAX1_12/B FAX1_12/a_25_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6666 gnd OAI22X1_48/Y OAI21X1_128/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M6667 vdd INVX2_52/A AOI21X1_12/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M6668 AOI21X1_12/A INVX2_52/A OAI21X1_128/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6669 AOI21X1_12/A OAI22X1_47/Y OAI21X1_128/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6670 OAI21X1_128/a_9_54# OAI22X1_48/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6671 OAI21X1_128/a_2_6# OAI22X1_47/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6672 gnd INVX2_55/Y OAI21X1_106/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M6673 vdd NAND2X1_93/Y OAI21X1_106/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M6674 OAI21X1_106/Y NAND2X1_93/Y OAI21X1_106/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6675 OAI21X1_106/Y BUFX2_23/Y OAI21X1_106/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6676 OAI21X1_106/a_9_54# INVX2_55/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6677 OAI21X1_106/a_2_6# BUFX2_23/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6678 gnd AND2X2_16/Y OAI21X1_117/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M6679 vdd OAI21X1_118/Y INVX2_50/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M6680 INVX2_50/A OAI21X1_118/Y OAI21X1_117/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6681 INVX2_50/A OAI21X1_1/B OAI21X1_117/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6682 OAI21X1_117/a_9_54# AND2X2_16/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6683 OAI21X1_117/a_2_6# OAI21X1_1/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6684 gnd AOI22X1_74/Y OAI21X1_139/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M6685 vdd OAI21X1_140/Y INVX2_40/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M6686 INVX2_40/A OAI21X1_140/Y OAI21X1_139/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6687 INVX2_40/A XOR2X1_11/Y OAI21X1_139/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6688 OAI21X1_139/a_9_54# AOI22X1_74/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6689 OAI21X1_139/a_2_6# XOR2X1_11/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6690 vdd in_clka BUFX2_4/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6691 gnd in_clka BUFX2_4/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M6692 BUFX2_5/A BUFX2_4/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6693 BUFX2_5/A BUFX2_4/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6694 XNOR2X1_28/A XOR2X1_24/A vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M6695 NAND2X1_101/a_9_6# XOR2X1_24/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6696 vdd XOR2X1_25/Y XNOR2X1_28/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6697 XNOR2X1_28/A XOR2X1_25/Y NAND2X1_101/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6698 FAX1_2/a_46_54# FAX1_2/A vdd vdd pfet w=40 l=2
+  ad=0.452n pd=0.176m as=0 ps=0
M6699 gnd FAX1_2/A FAX1_2/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M6700 gnd FAX1_2/A FAX1_2/a_84_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M6701 FAX1_2/a_33_6# in_incr[2] FAX1_2/a_25_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.12n ps=52u
M6702 FAX1_2/a_79_6# FAX1_2/C FAX1_2/a_70_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.14n ps=54u
M6703 FAX1_2/a_46_6# FAX1_2/A gnd Gnd nfet w=20 l=2
+  ad=0.24n pd=0.104m as=0 ps=0
M6704 FAX1_2/YS FAX1_2/a_70_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6705 FAX1_2/a_46_6# FAX1_2/C gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6706 FAX1_2/a_79_46# FAX1_2/C FAX1_2/a_70_6# vdd pfet w=48 l=2
+  ad=0.144n pd=0.102m as=0.317n ps=0.11m
M6707 FAX1_1/C FAX1_2/a_25_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6708 FAX1_2/a_2_54# in_incr[2] vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M6709 FAX1_2/a_25_6# FAX1_2/C FAX1_2/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6710 gnd FAX1_2/A FAX1_2/a_33_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6711 FAX1_2/a_70_6# FAX1_2/a_25_6# FAX1_2/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M6712 FAX1_2/a_84_6# in_incr[2] FAX1_2/a_79_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6713 vdd in_incr[2] FAX1_2/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M6714 vdd FAX1_2/A FAX1_2/a_84_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0.144n ps=0.102m
M6715 vdd FAX1_2/A FAX1_2/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6716 FAX1_2/YS FAX1_2/a_70_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M6717 FAX1_2/a_25_6# FAX1_2/C FAX1_2/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M6718 gnd in_incr[2] FAX1_2/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6719 vdd FAX1_2/A FAX1_2/a_33_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6720 FAX1_2/a_84_46# in_incr[2] FAX1_2/a_79_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0 ps=0
M6721 FAX1_2/a_70_6# FAX1_2/a_25_6# FAX1_2/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6722 FAX1_2/a_46_54# FAX1_2/C vdd vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M6723 FAX1_1/C FAX1_2/a_25_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M6724 FAX1_2/a_2_6# in_incr[2] gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6725 FAX1_2/a_33_54# in_incr[2] FAX1_2/a_25_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6726 OAI22X1_76/B INVX2_251/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M6727 NAND2X1_123/a_9_6# INVX2_251/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6728 vdd INVX2_37/Y OAI22X1_76/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6729 OAI22X1_76/B INVX2_37/Y NAND2X1_123/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6730 OAI22X1_52/D out_temp_data_in[0] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M6731 NAND2X1_112/a_9_6# out_temp_data_in[0] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6732 vdd INVX2_53/A OAI22X1_52/D vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6733 OAI22X1_52/D INVX2_53/A NAND2X1_112/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6734 INVX2_4/Y out_temp_index[3] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6735 INVX2_4/Y out_temp_index[3] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6736 AOI21X1_4/a_2_54# out_temp_decoded[2] vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M6737 AOI21X1_4/a_12_6# out_mines[2] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6738 gnd OAI22X1_0/Y AOI21X1_4/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0.11n ps=52u
M6739 vdd out_mines[2] AOI21X1_4/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6740 AOI21X1_4/Y OAI22X1_0/Y AOI21X1_4/a_2_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6741 AOI21X1_4/Y out_temp_decoded[2] AOI21X1_4/a_12_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6742 gnd XOR2X1_7/Y XNOR2X1_12/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6743 MUX2X1_3/A XOR2X1_7/Y XNOR2X1_12/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M6744 XNOR2X1_12/a_12_41# XOR2X1_8/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6745 XNOR2X1_12/a_18_54# XNOR2X1_12/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M6746 XNOR2X1_12/a_35_6# XNOR2X1_12/a_2_6# MUX2X1_3/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6747 XNOR2X1_12/a_18_6# XNOR2X1_12/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6748 vdd XOR2X1_7/Y XNOR2X1_12/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M6749 vdd XOR2X1_8/Y XNOR2X1_12/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6750 MUX2X1_3/A XNOR2X1_12/a_2_6# XNOR2X1_12/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M6751 XNOR2X1_12/a_35_54# XOR2X1_7/Y MUX2X1_3/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6752 XNOR2X1_12/a_12_41# XOR2X1_8/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6753 gnd XOR2X1_8/Y XNOR2X1_12/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6754 gnd out_temp_mine_cnt[1] XNOR2X1_23/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6755 XNOR2X1_23/Y out_temp_mine_cnt[1] XNOR2X1_23/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M6756 XNOR2X1_23/a_12_41# in_n_mines[1] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6757 XNOR2X1_23/a_18_54# XNOR2X1_23/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M6758 XNOR2X1_23/a_35_6# XNOR2X1_23/a_2_6# XNOR2X1_23/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6759 XNOR2X1_23/a_18_6# XNOR2X1_23/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6760 vdd out_temp_mine_cnt[1] XNOR2X1_23/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M6761 vdd in_n_mines[1] XNOR2X1_23/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6762 XNOR2X1_23/Y XNOR2X1_23/a_2_6# XNOR2X1_23/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M6763 XNOR2X1_23/a_35_54# out_temp_mine_cnt[1] XNOR2X1_23/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6764 XNOR2X1_23/a_12_41# in_n_mines[1] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6765 gnd in_n_mines[1] XNOR2X1_23/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6766 vdd BUFX2_9/A BUFX2_11/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6767 gnd BUFX2_9/A BUFX2_11/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M6768 BUFX2_11/Y BUFX2_11/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6769 BUFX2_11/Y BUFX2_11/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6770 vdd BUFX2_23/A BUFX2_22/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6771 gnd BUFX2_23/A BUFX2_22/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M6772 BUFX2_22/Y BUFX2_22/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6773 BUFX2_22/Y BUFX2_22/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6774 NOR2X1_2/Y NOR2X1_2/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M6775 NOR2X1_2/Y FAX1_2/YS NOR2X1_2/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M6776 NOR2X1_2/a_9_54# NOR2X1_2/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6777 gnd FAX1_2/YS NOR2X1_2/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6778 AOI21X1_12/a_2_54# AOI21X1_12/B vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M6779 AOI21X1_12/a_12_6# AOI21X1_12/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6780 gnd INVX2_51/Y AOI21X1_12/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0.11n ps=52u
M6781 vdd AOI21X1_12/A AOI21X1_12/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6782 AOI21X1_12/Y INVX2_51/Y AOI21X1_12/a_2_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6783 AOI21X1_12/Y AOI21X1_12/B AOI21X1_12/a_12_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6784 AOI21X1_23/a_2_54# OR2X1_16/Y vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M6785 AOI21X1_23/a_12_6# INVX2_123/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6786 gnd AOI21X1_23/C NOR2X1_119/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0.11n ps=52u
M6787 vdd INVX2_123/Y AOI21X1_23/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6788 NOR2X1_119/B AOI21X1_23/C AOI21X1_23/a_2_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6789 NOR2X1_119/B OR2X1_16/Y AOI21X1_23/a_12_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6790 vdd out_global_score[15] HAX1_15/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M6791 HAX1_15/a_41_74# HAX1_15/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M6792 HAX1_15/a_9_6# out_global_score[15] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6793 HAX1_15/a_41_74# HAX1_15/B HAX1_15/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M6794 vdd out_global_score[15] HAX1_15/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6795 vdd HAX1_15/a_2_74# HAX1_14/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6796 HAX1_15/a_38_6# HAX1_15/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6797 HAX1_15/YS HAX1_15/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6798 HAX1_15/a_38_6# out_global_score[15] HAX1_15/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6799 HAX1_15/YS HAX1_15/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M6800 HAX1_15/a_2_74# HAX1_15/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6801 HAX1_15/a_2_74# HAX1_15/B HAX1_15/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6802 HAX1_15/a_49_54# HAX1_15/B HAX1_15/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6803 gnd HAX1_15/a_2_74# HAX1_14/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M6804 vdd HAX1_48/A HAX1_48/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M6805 HAX1_48/a_41_74# HAX1_48/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M6806 HAX1_48/a_9_6# HAX1_48/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6807 HAX1_48/a_41_74# HAX1_48/B HAX1_48/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M6808 vdd HAX1_48/A HAX1_48/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6809 vdd HAX1_48/a_2_74# HAX1_49/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6810 HAX1_48/a_38_6# HAX1_48/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6811 HAX1_48/YS HAX1_48/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6812 HAX1_48/a_38_6# HAX1_48/A HAX1_48/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6813 HAX1_48/YS HAX1_48/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M6814 HAX1_48/a_2_74# HAX1_48/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6815 HAX1_48/a_2_74# HAX1_48/B HAX1_48/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6816 HAX1_48/a_49_54# HAX1_48/B HAX1_48/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6817 gnd HAX1_48/a_2_74# HAX1_49/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M6818 vdd out_global_score[4] HAX1_26/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M6819 HAX1_26/a_41_74# HAX1_26/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M6820 HAX1_26/a_9_6# out_global_score[4] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6821 HAX1_26/a_41_74# HAX1_26/B HAX1_26/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M6822 vdd out_global_score[4] HAX1_26/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6823 vdd HAX1_26/a_2_74# HAX1_25/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6824 HAX1_26/a_38_6# HAX1_26/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6825 HAX1_26/YS HAX1_26/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6826 HAX1_26/a_38_6# out_global_score[4] HAX1_26/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6827 HAX1_26/YS HAX1_26/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M6828 HAX1_26/a_2_74# HAX1_26/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6829 HAX1_26/a_2_74# HAX1_26/B HAX1_26/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6830 HAX1_26/a_49_54# HAX1_26/B HAX1_26/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6831 gnd HAX1_26/a_2_74# HAX1_25/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M6832 vdd out_temp_mine_cnt[1] HAX1_37/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M6833 HAX1_37/a_41_74# HAX1_37/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M6834 HAX1_37/a_9_6# out_temp_mine_cnt[1] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6835 HAX1_37/a_41_74# out_temp_mine_cnt[0] HAX1_37/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M6836 vdd out_temp_mine_cnt[1] HAX1_37/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6837 vdd HAX1_37/a_2_74# HAX1_36/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6838 HAX1_37/a_38_6# HAX1_37/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6839 HAX1_37/YS HAX1_37/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6840 HAX1_37/a_38_6# out_temp_mine_cnt[1] HAX1_37/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6841 HAX1_37/YS HAX1_37/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M6842 HAX1_37/a_2_74# out_temp_mine_cnt[0] vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6843 HAX1_37/a_2_74# out_temp_mine_cnt[0] HAX1_37/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6844 HAX1_37/a_49_54# out_temp_mine_cnt[0] HAX1_37/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6845 gnd HAX1_37/a_2_74# HAX1_36/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M6846 gnd OAI21X1_7/A OAI21X1_7/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M6847 vdd OAI21X1_7/C OAI21X1_7/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M6848 OAI21X1_7/Y OAI21X1_7/C OAI21X1_7/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6849 OAI21X1_7/Y OAI21X1_9/B OAI21X1_7/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6850 OAI21X1_7/a_9_54# OAI21X1_7/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6851 OAI21X1_7/a_2_6# OAI21X1_9/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6852 gnd out_mines[1] OAI22X1_42/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M6853 OAI22X1_42/a_2_6# out_mines[0] OAI22X1_42/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M6854 OAI22X1_42/Y OAI22X1_52/D OAI22X1_42/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6855 OAI22X1_42/Y OAI22X1_52/B OAI22X1_42/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M6856 OAI22X1_42/a_28_54# OAI22X1_52/D OAI22X1_42/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M6857 OAI22X1_42/a_9_54# out_mines[1] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6858 OAI22X1_42/a_2_6# OAI22X1_52/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6859 vdd out_mines[0] OAI22X1_42/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6860 gnd BUFX2_24/Y OAI22X1_20/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M6861 OAI22X1_20/a_2_6# OR2X1_11/A OAI22X1_20/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M6862 OAI22X1_20/Y INVX2_74/Y OAI22X1_20/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6863 OAI22X1_20/Y OAI22X1_1/B OAI22X1_20/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M6864 OAI22X1_20/a_28_54# INVX2_74/Y OAI22X1_20/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M6865 OAI22X1_20/a_9_54# BUFX2_24/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6866 OAI22X1_20/a_2_6# OAI22X1_1/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6867 vdd OR2X1_11/A OAI22X1_20/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6868 gnd INVX2_44/Y OAI22X1_31/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M6869 OAI22X1_31/a_2_6# INVX2_48/Y XNOR2X1_26/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M6870 XNOR2X1_26/A XOR2X1_20/Y OAI22X1_31/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6871 XNOR2X1_26/A INVX2_49/A OAI22X1_31/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M6872 OAI22X1_31/a_28_54# XOR2X1_20/Y XNOR2X1_26/A vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M6873 OAI22X1_31/a_9_54# INVX2_44/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6874 OAI22X1_31/a_2_6# INVX2_49/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6875 vdd INVX2_48/Y OAI22X1_31/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6876 gnd out_mines[23] OAI22X1_75/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M6877 OAI22X1_75/a_2_6# out_mines[22] OAI22X1_75/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M6878 OAI22X1_75/Y OAI22X1_75/D OAI22X1_75/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6879 OAI22X1_75/Y OAI22X1_75/B OAI22X1_75/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M6880 OAI22X1_75/a_28_54# OAI22X1_75/D OAI22X1_75/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M6881 OAI22X1_75/a_9_54# out_mines[23] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6882 OAI22X1_75/a_2_6# OAI22X1_75/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6883 vdd out_mines[22] OAI22X1_75/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6884 gnd out_mines[3] OAI22X1_53/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M6885 OAI22X1_53/a_2_6# out_mines[2] OAI22X1_53/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M6886 OAI22X1_53/Y OAI22X1_63/D OAI22X1_53/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6887 OAI22X1_53/Y OAI22X1_63/B OAI22X1_53/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M6888 OAI22X1_53/a_28_54# OAI22X1_63/D OAI22X1_53/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M6889 OAI22X1_53/a_9_54# out_mines[3] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6890 OAI22X1_53/a_2_6# OAI22X1_63/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6891 vdd out_mines[2] OAI22X1_53/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6892 gnd out_mines[21] OAI22X1_64/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M6893 OAI22X1_64/a_2_6# out_mines[20] OAI22X1_64/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M6894 OAI22X1_64/Y OAI22X1_64/D OAI22X1_64/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6895 OAI22X1_64/Y OAI22X1_64/B OAI22X1_64/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M6896 OAI22X1_64/a_28_54# OAI22X1_64/D OAI22X1_64/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M6897 OAI22X1_64/a_9_54# out_mines[21] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6898 OAI22X1_64/a_2_6# OAI22X1_64/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6899 vdd out_mines[20] OAI22X1_64/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6900 gnd out_mines[17] OAI22X1_86/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M6901 OAI22X1_86/a_2_6# out_mines[16] OAI22X1_86/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M6902 OAI22X1_86/Y OAI22X1_88/D OAI22X1_86/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6903 OAI22X1_86/Y OAI22X1_88/B OAI22X1_86/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M6904 OAI22X1_86/a_28_54# OAI22X1_88/D OAI22X1_86/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M6905 OAI22X1_86/a_9_54# out_mines[17] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6906 OAI22X1_86/a_2_6# OAI22X1_88/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6907 vdd out_mines[16] OAI22X1_86/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6908 DFFNEGX1_5/a_76_6# BUFX2_17/Y DFFNEGX1_5/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M6909 gnd BUFX2_17/Y DFFNEGX1_5/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6910 DFFNEGX1_5/a_66_6# DFFNEGX1_5/a_2_6# DFFNEGX1_5/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M6911 out_mines[7] DFFNEGX1_5/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6912 DFFNEGX1_5/a_23_6# BUFX2_17/Y DFFNEGX1_5/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M6913 DFFNEGX1_5/a_23_6# DFFNEGX1_5/a_2_6# DFFNEGX1_5/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M6914 gnd DFFNEGX1_5/a_34_4# DFFNEGX1_5/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M6915 vdd DFFNEGX1_5/a_34_4# DFFNEGX1_5/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M6916 DFFNEGX1_5/a_61_74# DFFNEGX1_5/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M6917 DFFNEGX1_5/a_34_4# DFFNEGX1_5/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6918 DFFNEGX1_5/a_34_4# DFFNEGX1_5/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M6919 vdd out_mines[7] DFFNEGX1_5/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M6920 gnd out_mines[7] DFFNEGX1_5/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6921 DFFNEGX1_5/a_61_6# DFFNEGX1_5/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6922 DFFNEGX1_5/a_76_84# DFFNEGX1_5/a_2_6# DFFNEGX1_5/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M6923 out_mines[7] DFFNEGX1_5/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6924 vdd BUFX2_17/Y DFFNEGX1_5/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M6925 DFFNEGX1_5/a_31_6# DFFNEGX1_5/a_2_6# DFFNEGX1_5/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6926 DFFNEGX1_5/a_66_6# BUFX2_17/Y DFFNEGX1_5/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6927 DFFNEGX1_5/a_17_74# OAI21X1_37/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6928 DFFNEGX1_5/a_31_74# BUFX2_17/Y DFFNEGX1_5/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6929 DFFNEGX1_5/a_17_6# OAI21X1_37/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M6930 OAI22X1_1/D out_temp_cleared[7] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6931 OAI22X1_1/D out_temp_cleared[7] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6932 INVX2_128/Y INVX2_128/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6933 INVX2_128/Y INVX2_128/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6934 INVX2_117/Y INVX2_117/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6935 INVX2_117/Y INVX2_117/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6936 MUX2X1_24/A FAX1_2/YS gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6937 MUX2X1_24/A FAX1_2/YS vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6938 FAX1_13/a_46_54# FAX1_13/A vdd vdd pfet w=40 l=2
+  ad=0.452n pd=0.176m as=0 ps=0
M6939 gnd FAX1_13/A FAX1_13/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M6940 gnd FAX1_13/A FAX1_13/a_84_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M6941 FAX1_13/a_33_6# FAX1_13/B FAX1_13/a_25_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.12n ps=52u
M6942 FAX1_13/a_79_6# FAX1_13/C FAX1_13/a_70_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.14n ps=54u
M6943 FAX1_13/a_46_6# FAX1_13/A gnd Gnd nfet w=20 l=2
+  ad=0.24n pd=0.104m as=0 ps=0
M6944 FAX1_12/B FAX1_13/a_70_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6945 FAX1_13/a_46_6# FAX1_13/C gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6946 FAX1_13/a_79_46# FAX1_13/C FAX1_13/a_70_6# vdd pfet w=48 l=2
+  ad=0.144n pd=0.102m as=0.317n ps=0.11m
M6947 FAX1_11/C FAX1_13/a_25_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6948 FAX1_13/a_2_54# FAX1_13/B vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M6949 FAX1_13/a_25_6# FAX1_13/C FAX1_13/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6950 gnd FAX1_13/A FAX1_13/a_33_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6951 FAX1_13/a_70_6# FAX1_13/a_25_6# FAX1_13/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M6952 FAX1_13/a_84_6# FAX1_13/B FAX1_13/a_79_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6953 vdd FAX1_13/B FAX1_13/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M6954 vdd FAX1_13/A FAX1_13/a_84_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0.144n ps=0.102m
M6955 vdd FAX1_13/A FAX1_13/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6956 FAX1_12/B FAX1_13/a_70_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M6957 FAX1_13/a_25_6# FAX1_13/C FAX1_13/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M6958 gnd FAX1_13/B FAX1_13/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6959 vdd FAX1_13/A FAX1_13/a_33_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6960 FAX1_13/a_84_46# FAX1_13/B FAX1_13/a_79_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0 ps=0
M6961 FAX1_13/a_70_6# FAX1_13/a_25_6# FAX1_13/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6962 FAX1_13/a_46_54# FAX1_13/C vdd vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M6963 FAX1_11/C FAX1_13/a_25_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M6964 FAX1_13/a_2_6# FAX1_13/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6965 FAX1_13/a_33_54# FAX1_13/B FAX1_13/a_25_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6966 gnd OAI22X1_50/Y OAI21X1_129/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M6967 vdd INVX2_52/Y OAI21X1_129/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M6968 OAI21X1_129/Y INVX2_52/Y OAI21X1_129/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6969 OAI21X1_129/Y OAI22X1_49/Y OAI21X1_129/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6970 OAI21X1_129/a_9_54# OAI22X1_50/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6971 OAI21X1_129/a_2_6# OAI22X1_49/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6972 gnd INVX2_251/Y OAI21X1_107/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M6973 vdd NAND2X1_96/Y OAI21X1_107/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M6974 OAI21X1_107/Y NAND2X1_96/Y OAI21X1_107/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6975 OAI21X1_107/Y INVX2_217/Y OAI21X1_107/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6976 OAI21X1_107/a_9_54# INVX2_251/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6977 OAI21X1_107/a_2_6# INVX2_217/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6978 gnd NOR2X1_110/Y OAI21X1_118/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M6979 vdd OAI21X1_1/B OAI21X1_118/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M6980 OAI21X1_118/Y OAI21X1_1/B OAI21X1_118/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6981 OAI21X1_118/Y INVX2_46/Y OAI21X1_118/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M6982 OAI21X1_118/a_9_54# NOR2X1_110/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M6983 OAI21X1_118/a_2_6# INVX2_46/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6984 vdd BUFX2_5/A BUFX2_5/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M6985 gnd BUFX2_5/A BUFX2_5/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M6986 BUFX2_5/Y BUFX2_5/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M6987 BUFX2_5/Y BUFX2_5/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6988 FAX1_3/a_46_54# FAX1_3/A vdd vdd pfet w=40 l=2
+  ad=0.452n pd=0.176m as=0 ps=0
M6989 gnd FAX1_3/A FAX1_3/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M6990 gnd FAX1_3/A FAX1_3/a_84_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M6991 FAX1_3/a_33_6# in_incr[1] FAX1_3/a_25_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.12n ps=52u
M6992 FAX1_3/a_79_6# FAX1_3/C FAX1_3/a_70_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.14n ps=54u
M6993 FAX1_3/a_46_6# FAX1_3/A gnd Gnd nfet w=20 l=2
+  ad=0.24n pd=0.104m as=0 ps=0
M6994 FAX1_3/YS FAX1_3/a_70_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6995 FAX1_3/a_46_6# FAX1_3/C gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M6996 FAX1_3/a_79_46# FAX1_3/C FAX1_3/a_70_6# vdd pfet w=48 l=2
+  ad=0.144n pd=0.102m as=0.317n ps=0.11m
M6997 FAX1_2/C FAX1_3/a_25_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M6998 FAX1_3/a_2_54# in_incr[1] vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M6999 FAX1_3/a_25_6# FAX1_3/C FAX1_3/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7000 gnd FAX1_3/A FAX1_3/a_33_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7001 FAX1_3/a_70_6# FAX1_3/a_25_6# FAX1_3/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M7002 FAX1_3/a_84_6# in_incr[1] FAX1_3/a_79_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7003 vdd in_incr[1] FAX1_3/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M7004 vdd FAX1_3/A FAX1_3/a_84_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0.144n ps=0.102m
M7005 vdd FAX1_3/A FAX1_3/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7006 FAX1_3/YS FAX1_3/a_70_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M7007 FAX1_3/a_25_6# FAX1_3/C FAX1_3/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M7008 gnd in_incr[1] FAX1_3/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7009 vdd FAX1_3/A FAX1_3/a_33_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7010 FAX1_3/a_84_46# in_incr[1] FAX1_3/a_79_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0 ps=0
M7011 FAX1_3/a_70_6# FAX1_3/a_25_6# FAX1_3/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7012 FAX1_3/a_46_54# FAX1_3/C vdd vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M7013 FAX1_2/C FAX1_3/a_25_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M7014 FAX1_3/a_2_6# in_incr[1] gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7015 FAX1_3/a_33_54# in_incr[1] FAX1_3/a_25_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7016 AOI22X1_75/A OAI21X1_154/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M7017 NAND2X1_124/a_9_6# OAI21X1_154/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7018 vdd OAI21X1_153/Y AOI22X1_75/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7019 AOI22X1_75/A OAI21X1_153/Y NAND2X1_124/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7020 INVX2_41/A out_temp_data_in[0] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M7021 NAND2X1_102/a_9_6# out_temp_data_in[0] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7022 vdd INVX2_32/Y INVX2_41/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7023 INVX2_41/A INVX2_32/Y NAND2X1_102/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7024 OAI22X1_52/B INVX2_251/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M7025 NAND2X1_113/a_9_6# INVX2_251/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7026 vdd INVX2_53/A OAI22X1_52/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7027 OAI22X1_52/B INVX2_53/A NAND2X1_113/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7028 HAX1_48/B NOR2X1_0/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M7029 NAND2X1_0/a_9_6# NOR2X1_0/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7030 vdd XNOR2X1_1/A HAX1_48/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7031 HAX1_48/B XNOR2X1_1/A NAND2X1_0/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7032 INVX2_5/Y out_mines[7] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7033 INVX2_5/Y out_mines[7] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7034 AOI21X1_5/a_2_54# INVX2_18/Y vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M7035 AOI21X1_5/a_12_6# NOR2X1_92/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7036 gnd AOI21X1_5/C AOI21X1_5/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0.11n ps=52u
M7037 vdd NOR2X1_92/Y AOI21X1_5/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7038 AOI21X1_5/Y AOI21X1_5/C AOI21X1_5/a_2_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7039 AOI21X1_5/Y INVX2_18/Y AOI21X1_5/a_12_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7040 gnd NAND2X1_6/B XNOR2X1_13/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M7041 MUX2X1_2/A NAND2X1_6/B XNOR2X1_13/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M7042 XNOR2X1_13/a_12_41# NOR2X1_6/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7043 XNOR2X1_13/a_18_54# XNOR2X1_13/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7044 XNOR2X1_13/a_35_6# XNOR2X1_13/a_2_6# MUX2X1_2/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7045 XNOR2X1_13/a_18_6# XNOR2X1_13/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7046 vdd NAND2X1_6/B XNOR2X1_13/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M7047 vdd NOR2X1_6/Y XNOR2X1_13/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7048 MUX2X1_2/A XNOR2X1_13/a_2_6# XNOR2X1_13/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M7049 XNOR2X1_13/a_35_54# NAND2X1_6/B MUX2X1_2/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7050 XNOR2X1_13/a_12_41# NOR2X1_6/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7051 gnd NOR2X1_6/Y XNOR2X1_13/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7052 gnd out_temp_mine_cnt[3] XNOR2X1_24/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M7053 XNOR2X1_24/Y out_temp_mine_cnt[3] XNOR2X1_24/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M7054 XNOR2X1_24/a_12_41# in_n_mines[3] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7055 XNOR2X1_24/a_18_54# XNOR2X1_24/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7056 XNOR2X1_24/a_35_6# XNOR2X1_24/a_2_6# XNOR2X1_24/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7057 XNOR2X1_24/a_18_6# XNOR2X1_24/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7058 vdd out_temp_mine_cnt[3] XNOR2X1_24/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M7059 vdd in_n_mines[3] XNOR2X1_24/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7060 XNOR2X1_24/Y XNOR2X1_24/a_2_6# XNOR2X1_24/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M7061 XNOR2X1_24/a_35_54# out_temp_mine_cnt[3] XNOR2X1_24/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7062 XNOR2X1_24/a_12_41# in_n_mines[3] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7063 gnd in_n_mines[3] XNOR2X1_24/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7064 vdd BUFX2_23/A BUFX2_23/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M7065 gnd BUFX2_23/A BUFX2_23/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M7066 BUFX2_23/Y BUFX2_23/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7067 BUFX2_23/Y BUFX2_23/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7068 vdd BUFX2_1/Y BUFX2_12/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M7069 gnd BUFX2_1/Y BUFX2_12/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M7070 BUFX2_12/Y BUFX2_12/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7071 BUFX2_12/Y BUFX2_12/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7072 NOR2X1_3/Y NOR2X1_3/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M7073 NOR2X1_3/Y FAX1_1/YS NOR2X1_3/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M7074 NOR2X1_3/a_9_54# NOR2X1_3/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7075 gnd FAX1_1/YS NOR2X1_3/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7076 AOI21X1_24/a_2_54# AND2X2_19/Y vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M7077 AOI21X1_24/a_12_6# AOI21X1_25/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7078 gnd BUFX2_3/Y AOI21X1_24/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0.11n ps=52u
M7079 vdd AOI21X1_25/Y AOI21X1_24/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7080 AOI21X1_24/Y BUFX2_3/Y AOI21X1_24/a_2_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7081 AOI21X1_24/Y AND2X2_19/Y AOI21X1_24/a_12_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7082 AOI21X1_13/a_2_54# AOI21X1_13/B vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M7083 AOI21X1_13/a_12_6# AOI21X1_13/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7084 gnd INVX2_34/A AOI21X1_13/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0.11n ps=52u
M7085 vdd AOI21X1_13/A AOI21X1_13/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7086 AOI21X1_13/Y INVX2_34/A AOI21X1_13/a_2_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7087 AOI21X1_13/Y AOI21X1_13/B AOI21X1_13/a_12_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7088 vdd HAX1_38/A HAX1_38/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M7089 HAX1_38/a_41_74# HAX1_38/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M7090 HAX1_38/a_9_6# HAX1_38/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7091 HAX1_38/a_41_74# HAX1_38/B HAX1_38/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M7092 vdd HAX1_38/A HAX1_38/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7093 vdd HAX1_38/a_2_74# HAX1_39/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M7094 HAX1_38/a_38_6# HAX1_38/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7095 MUX2X1_6/A HAX1_38/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7096 HAX1_38/a_38_6# HAX1_38/A HAX1_38/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7097 MUX2X1_6/A HAX1_38/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M7098 HAX1_38/a_2_74# HAX1_38/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7099 HAX1_38/a_2_74# HAX1_38/B HAX1_38/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7100 HAX1_38/a_49_54# HAX1_38/B HAX1_38/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7101 gnd HAX1_38/a_2_74# HAX1_39/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M7102 vdd out_global_score[14] HAX1_16/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M7103 HAX1_16/a_41_74# HAX1_16/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M7104 HAX1_16/a_9_6# out_global_score[14] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7105 HAX1_16/a_41_74# HAX1_16/B HAX1_16/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M7106 vdd out_global_score[14] HAX1_16/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7107 vdd HAX1_16/a_2_74# HAX1_15/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M7108 HAX1_16/a_38_6# HAX1_16/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7109 HAX1_16/YS HAX1_16/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7110 HAX1_16/a_38_6# out_global_score[14] HAX1_16/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7111 HAX1_16/YS HAX1_16/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M7112 HAX1_16/a_2_74# HAX1_16/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7113 HAX1_16/a_2_74# HAX1_16/B HAX1_16/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7114 HAX1_16/a_49_54# HAX1_16/B HAX1_16/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7115 gnd HAX1_16/a_2_74# HAX1_15/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M7116 vdd out_global_score[3] HAX1_27/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M7117 HAX1_27/a_41_74# HAX1_27/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M7118 HAX1_27/a_9_6# out_global_score[3] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7119 HAX1_27/a_41_74# HAX1_27/B HAX1_27/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M7120 vdd out_global_score[3] HAX1_27/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7121 vdd HAX1_27/a_2_74# HAX1_26/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M7122 HAX1_27/a_38_6# HAX1_27/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7123 HAX1_27/YS HAX1_27/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7124 HAX1_27/a_38_6# out_global_score[3] HAX1_27/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7125 HAX1_27/YS HAX1_27/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M7126 HAX1_27/a_2_74# HAX1_27/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7127 HAX1_27/a_2_74# HAX1_27/B HAX1_27/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7128 HAX1_27/a_49_54# HAX1_27/B HAX1_27/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7129 gnd HAX1_27/a_2_74# HAX1_26/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M7130 vdd HAX1_49/A HAX1_49/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M7131 HAX1_49/a_41_74# HAX1_49/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M7132 HAX1_49/a_9_6# HAX1_49/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7133 HAX1_49/a_41_74# HAX1_49/B HAX1_49/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M7134 vdd HAX1_49/A HAX1_49/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7135 vdd HAX1_49/a_2_74# OR2X1_0/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M7136 HAX1_49/a_38_6# HAX1_49/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7137 HAX1_49/YS HAX1_49/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7138 HAX1_49/a_38_6# HAX1_49/A HAX1_49/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7139 HAX1_49/YS HAX1_49/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M7140 HAX1_49/a_2_74# HAX1_49/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7141 HAX1_49/a_2_74# HAX1_49/B HAX1_49/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7142 HAX1_49/a_49_54# HAX1_49/B HAX1_49/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7143 gnd HAX1_49/a_2_74# OR2X1_0/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M7144 OR2X1_0/a_2_54# OR2X1_0/A gnd Gnd nfet w=10 l=2
+  ad=29.999998p pd=16u as=50p ps=30u
M7145 OR2X1_0/Y OR2X1_0/a_2_54# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0.11n ps=46u
M7146 OR2X1_0/Y OR2X1_0/a_2_54# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=29.999998p ps=16u
M7147 vdd OR2X1_0/B OR2X1_0/a_9_54# vdd pfet w=40 l=2
+  ad=0.11n pd=46u as=59.999996p ps=43u
M7148 OR2X1_0/a_9_54# OR2X1_0/A OR2X1_0/a_2_54# vdd pfet w=40 l=2
+  ad=59.999996p pd=43u as=0.2n ps=90u
M7149 gnd OR2X1_0/B OR2X1_0/a_2_54# Gnd nfet w=10 l=2
+  ad=29.999998p pd=16u as=29.999998p ps=16u
M7150 gnd OAI21X1_8/A OAI21X1_8/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M7151 vdd BUFX2_19/Y OAI21X1_8/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M7152 OAI21X1_8/Y BUFX2_19/Y OAI21X1_8/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7153 OAI21X1_8/Y OAI21X1_8/B OAI21X1_8/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7154 OAI21X1_8/a_9_54# OAI21X1_8/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7155 OAI21X1_8/a_2_6# OAI21X1_8/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7156 gnd BUFX2_24/Y OAI22X1_21/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M7157 OAI22X1_21/a_2_6# OAI22X1_5/C OAI22X1_21/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M7158 OAI22X1_21/Y INVX2_75/Y OAI22X1_21/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7159 OAI22X1_21/Y OAI22X1_1/D OAI22X1_21/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M7160 OAI22X1_21/a_28_54# INVX2_75/Y OAI22X1_21/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7161 OAI22X1_21/a_9_54# BUFX2_24/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7162 OAI22X1_21/a_2_6# OAI22X1_1/D gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7163 vdd OAI22X1_5/C OAI22X1_21/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7164 gnd BUFX2_25/Y OAI22X1_10/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M7165 OAI22X1_10/a_2_6# OR2X1_11/A OAI22X1_10/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M7166 OAI22X1_10/Y INVX2_63/Y OAI22X1_10/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7167 OAI22X1_10/Y INVX2_95/Y OAI22X1_10/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M7168 OAI22X1_10/a_28_54# INVX2_63/Y OAI22X1_10/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7169 OAI22X1_10/a_9_54# BUFX2_25/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7170 OAI22X1_10/a_2_6# INVX2_95/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7171 vdd OR2X1_11/A OAI22X1_10/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7172 gnd XOR2X1_29/Y OAI22X1_32/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M7173 OAI22X1_32/a_2_6# INVX2_40/A XNOR2X1_27/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M7174 XNOR2X1_27/A XOR2X1_29/B OAI22X1_32/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7175 XNOR2X1_27/A XOR2X1_28/A OAI22X1_32/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M7176 OAI22X1_32/a_28_54# XOR2X1_29/B XNOR2X1_27/A vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7177 OAI22X1_32/a_9_54# XOR2X1_29/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7178 OAI22X1_32/a_2_6# XOR2X1_28/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7179 vdd INVX2_40/A OAI22X1_32/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7180 gnd out_mines[7] OAI22X1_43/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M7181 OAI22X1_43/a_2_6# out_mines[6] OAI22X1_43/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M7182 OAI22X1_43/Y OAI22X1_51/D OAI22X1_43/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7183 OAI22X1_43/Y OAI22X1_51/B OAI22X1_43/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M7184 OAI22X1_43/a_28_54# OAI22X1_51/D OAI22X1_43/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7185 OAI22X1_43/a_9_54# out_mines[7] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7186 OAI22X1_43/a_2_6# OAI22X1_51/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7187 vdd out_mines[6] OAI22X1_43/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7188 gnd out_mines[21] OAI22X1_76/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M7189 OAI22X1_76/a_2_6# out_mines[20] OAI22X1_76/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M7190 OAI22X1_76/Y OAI22X1_76/D OAI22X1_76/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7191 OAI22X1_76/Y OAI22X1_76/B OAI22X1_76/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M7192 OAI22X1_76/a_28_54# OAI22X1_76/D OAI22X1_76/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7193 OAI22X1_76/a_9_54# out_mines[21] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7194 OAI22X1_76/a_2_6# OAI22X1_76/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7195 vdd out_mines[20] OAI22X1_76/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7196 gnd out_mines[3] OAI22X1_65/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M7197 OAI22X1_65/a_2_6# out_mines[2] OAI22X1_65/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M7198 OAI22X1_65/Y OAI22X1_75/D OAI22X1_65/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7199 OAI22X1_65/Y OAI22X1_75/B OAI22X1_65/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M7200 OAI22X1_65/a_28_54# OAI22X1_75/D OAI22X1_65/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7201 OAI22X1_65/a_9_54# out_mines[3] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7202 OAI22X1_65/a_2_6# OAI22X1_75/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7203 vdd out_mines[2] OAI22X1_65/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7204 gnd out_mines[1] OAI22X1_54/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M7205 OAI22X1_54/a_2_6# out_mines[0] OAI22X1_54/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M7206 OAI22X1_54/Y OAI22X1_64/D OAI22X1_54/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7207 OAI22X1_54/Y OAI22X1_64/B OAI22X1_54/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M7208 OAI22X1_54/a_28_54# OAI22X1_64/D OAI22X1_54/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7209 OAI22X1_54/a_9_54# out_mines[1] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7210 OAI22X1_54/a_2_6# OAI22X1_64/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7211 vdd out_mines[0] OAI22X1_54/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7212 gnd out_mines[23] OAI22X1_87/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M7213 OAI22X1_87/a_2_6# out_mines[22] OAI22X1_87/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M7214 OAI22X1_87/Y OAI22X1_87/D OAI22X1_87/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7215 OAI22X1_87/Y OAI22X1_87/B OAI22X1_87/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M7216 OAI22X1_87/a_28_54# OAI22X1_87/D OAI22X1_87/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7217 OAI22X1_87/a_9_54# out_mines[23] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7218 OAI22X1_87/a_2_6# OAI22X1_87/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7219 vdd out_mines[22] OAI22X1_87/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7220 DFFNEGX1_6/a_76_6# BUFX2_17/Y DFFNEGX1_6/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M7221 gnd BUFX2_17/Y DFFNEGX1_6/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M7222 DFFNEGX1_6/a_66_6# DFFNEGX1_6/a_2_6# DFFNEGX1_6/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M7223 out_mines[5] DFFNEGX1_6/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7224 DFFNEGX1_6/a_23_6# BUFX2_17/Y DFFNEGX1_6/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M7225 DFFNEGX1_6/a_23_6# DFFNEGX1_6/a_2_6# DFFNEGX1_6/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M7226 gnd DFFNEGX1_6/a_34_4# DFFNEGX1_6/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M7227 vdd DFFNEGX1_6/a_34_4# DFFNEGX1_6/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M7228 DFFNEGX1_6/a_61_74# DFFNEGX1_6/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7229 DFFNEGX1_6/a_34_4# DFFNEGX1_6/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7230 DFFNEGX1_6/a_34_4# DFFNEGX1_6/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M7231 vdd out_mines[5] DFFNEGX1_6/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M7232 gnd out_mines[5] DFFNEGX1_6/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7233 DFFNEGX1_6/a_61_6# DFFNEGX1_6/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7234 DFFNEGX1_6/a_76_84# DFFNEGX1_6/a_2_6# DFFNEGX1_6/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M7235 out_mines[5] DFFNEGX1_6/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7236 vdd BUFX2_17/Y DFFNEGX1_6/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M7237 DFFNEGX1_6/a_31_6# DFFNEGX1_6/a_2_6# DFFNEGX1_6/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7238 DFFNEGX1_6/a_66_6# BUFX2_17/Y DFFNEGX1_6/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7239 DFFNEGX1_6/a_17_74# OAI21X1_41/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7240 DFFNEGX1_6/a_31_74# BUFX2_17/Y DFFNEGX1_6/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7241 DFFNEGX1_6/a_17_6# OAI21X1_41/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7242 INVX2_107/Y out_temp_cleared[6] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7243 INVX2_107/Y out_temp_cleared[6] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7244 INVX2_129/Y out_load gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7245 INVX2_129/Y out_load vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7246 INVX2_118/Y out_state_main[3] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7247 INVX2_118/Y out_state_main[3] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7248 FAX1_14/a_46_54# FAX1_14/A vdd vdd pfet w=40 l=2
+  ad=0.452n pd=0.176m as=0 ps=0
M7249 gnd FAX1_14/A FAX1_14/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M7250 gnd FAX1_14/A FAX1_14/a_84_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M7251 FAX1_14/a_33_6# FAX1_14/B FAX1_14/a_25_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.12n ps=52u
M7252 FAX1_14/a_79_6# FAX1_14/C FAX1_14/a_70_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.14n ps=54u
M7253 FAX1_14/a_46_6# FAX1_14/A gnd Gnd nfet w=20 l=2
+  ad=0.24n pd=0.104m as=0 ps=0
M7254 FAX1_7/B FAX1_14/a_70_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7255 FAX1_14/a_46_6# FAX1_14/C gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7256 FAX1_14/a_79_46# FAX1_14/C FAX1_14/a_70_6# vdd pfet w=48 l=2
+  ad=0.144n pd=0.102m as=0.317n ps=0.11m
M7257 FAX1_6/A FAX1_14/a_25_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7258 FAX1_14/a_2_54# FAX1_14/B vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M7259 FAX1_14/a_25_6# FAX1_14/C FAX1_14/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7260 gnd FAX1_14/A FAX1_14/a_33_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7261 FAX1_14/a_70_6# FAX1_14/a_25_6# FAX1_14/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M7262 FAX1_14/a_84_6# FAX1_14/B FAX1_14/a_79_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7263 vdd FAX1_14/B FAX1_14/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M7264 vdd FAX1_14/A FAX1_14/a_84_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0.144n ps=0.102m
M7265 vdd FAX1_14/A FAX1_14/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7266 FAX1_7/B FAX1_14/a_70_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M7267 FAX1_14/a_25_6# FAX1_14/C FAX1_14/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M7268 gnd FAX1_14/B FAX1_14/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7269 vdd FAX1_14/A FAX1_14/a_33_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7270 FAX1_14/a_84_46# FAX1_14/B FAX1_14/a_79_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0 ps=0
M7271 FAX1_14/a_70_6# FAX1_14/a_25_6# FAX1_14/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7272 FAX1_14/a_46_54# FAX1_14/C vdd vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M7273 FAX1_6/A FAX1_14/a_25_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M7274 FAX1_14/a_2_6# FAX1_14/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7275 FAX1_14/a_33_54# FAX1_14/B FAX1_14/a_25_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7276 NOR2X1_90/Y NOR2X1_90/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M7277 NOR2X1_90/Y OAI22X1_3/Y NOR2X1_90/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M7278 NOR2X1_90/a_9_54# NOR2X1_90/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7279 gnd OAI22X1_3/Y NOR2X1_90/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7280 gnd OR2X1_6/A OAI21X1_108/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M7281 vdd NAND2X1_97/Y OAI21X1_108/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M7282 OAI21X1_108/Y NAND2X1_97/Y OAI21X1_108/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7283 OAI21X1_108/Y INVX2_217/Y OAI21X1_108/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7284 OAI21X1_108/a_9_54# OR2X1_6/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7285 OAI21X1_108/a_2_6# INVX2_217/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7286 gnd INVX2_20/Y OAI21X1_119/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M7287 vdd AOI22X1_67/Y AOI22X1_66/D vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M7288 AOI22X1_66/D AOI22X1_67/Y OAI21X1_119/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7289 AOI22X1_66/D NOR2X1_110/B OAI21X1_119/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7290 OAI21X1_119/a_9_54# INVX2_20/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7291 OAI21X1_119/a_2_6# NOR2X1_110/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7292 vdd BUFX2_8/A BUFX2_6/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M7293 gnd BUFX2_8/A BUFX2_6/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M7294 BUFX2_6/Y BUFX2_6/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7295 BUFX2_6/Y BUFX2_6/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7296 FAX1_4/a_46_54# FAX1_4/A vdd vdd pfet w=40 l=2
+  ad=0.452n pd=0.176m as=0 ps=0
M7297 gnd FAX1_4/A FAX1_4/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M7298 gnd FAX1_4/A FAX1_4/a_84_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M7299 FAX1_4/a_33_6# FAX1_4/B FAX1_4/a_25_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.12n ps=52u
M7300 FAX1_4/a_79_6# FAX1_4/C FAX1_4/a_70_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.14n ps=54u
M7301 FAX1_4/a_46_6# FAX1_4/A gnd Gnd nfet w=20 l=2
+  ad=0.24n pd=0.104m as=0 ps=0
M7302 FAX1_4/YS FAX1_4/a_70_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7303 FAX1_4/a_46_6# FAX1_4/C gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7304 FAX1_4/a_79_46# FAX1_4/C FAX1_4/a_70_6# vdd pfet w=48 l=2
+  ad=0.144n pd=0.102m as=0.317n ps=0.11m
M7305 FAX1_4/YC FAX1_4/a_25_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7306 FAX1_4/a_2_54# FAX1_4/B vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M7307 FAX1_4/a_25_6# FAX1_4/C FAX1_4/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7308 gnd FAX1_4/A FAX1_4/a_33_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7309 FAX1_4/a_70_6# FAX1_4/a_25_6# FAX1_4/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M7310 FAX1_4/a_84_6# FAX1_4/B FAX1_4/a_79_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7311 vdd FAX1_4/B FAX1_4/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M7312 vdd FAX1_4/A FAX1_4/a_84_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0.144n ps=0.102m
M7313 vdd FAX1_4/A FAX1_4/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7314 FAX1_4/YS FAX1_4/a_70_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M7315 FAX1_4/a_25_6# FAX1_4/C FAX1_4/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M7316 gnd FAX1_4/B FAX1_4/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7317 vdd FAX1_4/A FAX1_4/a_33_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7318 FAX1_4/a_84_46# FAX1_4/B FAX1_4/a_79_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0 ps=0
M7319 FAX1_4/a_70_6# FAX1_4/a_25_6# FAX1_4/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7320 FAX1_4/a_46_54# FAX1_4/C vdd vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M7321 FAX1_4/YC FAX1_4/a_25_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M7322 FAX1_4/a_2_6# FAX1_4/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7323 FAX1_4/a_33_54# FAX1_4/B FAX1_4/a_25_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7324 OAI22X1_87/D OR2X1_6/A vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M7325 NAND2X1_125/a_9_6# OR2X1_6/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7326 vdd INVX2_251/Y OAI22X1_87/D vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7327 OAI22X1_87/D INVX2_251/Y NAND2X1_125/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7328 OAI22X1_38/C out_temp_data_in[0] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M7329 NAND2X1_103/a_9_6# out_temp_data_in[0] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7330 vdd INVX2_31/Y OAI22X1_38/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7331 OAI22X1_38/C INVX2_31/Y NAND2X1_103/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7332 AOI22X1_73/A OAI21X1_138/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M7333 NAND2X1_114/a_9_6# OAI21X1_138/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7334 vdd OAI21X1_137/Y AOI22X1_73/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7335 AOI22X1_73/A OAI21X1_137/Y NAND2X1_114/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7336 HAX1_46/B NOR2X1_1/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M7337 NAND2X1_1/a_9_6# NOR2X1_1/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7338 vdd XNOR2X1_3/A HAX1_46/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7339 HAX1_46/B XNOR2X1_3/A NAND2X1_1/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7340 INVX2_6/Y out_mines[5] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7341 INVX2_6/Y out_mines[5] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7342 AOI21X1_6/a_2_54# INVX2_6/Y vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M7343 AOI21X1_6/a_12_6# NOR2X1_98/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7344 gnd AOI21X1_6/C AOI21X1_6/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0.11n ps=52u
M7345 vdd NOR2X1_98/Y AOI21X1_6/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7346 AOI21X1_6/Y AOI21X1_6/C AOI21X1_6/a_2_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7347 AOI21X1_6/Y INVX2_6/Y AOI21X1_6/a_12_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7348 gnd MUX2X1_0/B XNOR2X1_14/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M7349 MUX2X1_0/A MUX2X1_0/B XNOR2X1_14/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M7350 XNOR2X1_14/a_12_41# NOR2X1_7/B gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7351 XNOR2X1_14/a_18_54# XNOR2X1_14/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7352 XNOR2X1_14/a_35_6# XNOR2X1_14/a_2_6# MUX2X1_0/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7353 XNOR2X1_14/a_18_6# XNOR2X1_14/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7354 vdd MUX2X1_0/B XNOR2X1_14/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M7355 vdd NOR2X1_7/B XNOR2X1_14/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7356 MUX2X1_0/A XNOR2X1_14/a_2_6# XNOR2X1_14/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M7357 XNOR2X1_14/a_35_54# MUX2X1_0/B MUX2X1_0/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7358 XNOR2X1_14/a_12_41# NOR2X1_7/B vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7359 gnd NOR2X1_7/B XNOR2X1_14/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7360 gnd XNOR2X1_25/A XNOR2X1_25/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M7361 AOI22X1_1/A XNOR2X1_25/A XNOR2X1_25/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M7362 XNOR2X1_25/a_12_41# XNOR2X1_25/B gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7363 XNOR2X1_25/a_18_54# XNOR2X1_25/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7364 XNOR2X1_25/a_35_6# XNOR2X1_25/a_2_6# AOI22X1_1/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7365 XNOR2X1_25/a_18_6# XNOR2X1_25/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7366 vdd XNOR2X1_25/A XNOR2X1_25/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M7367 vdd XNOR2X1_25/B XNOR2X1_25/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7368 AOI22X1_1/A XNOR2X1_25/a_2_6# XNOR2X1_25/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M7369 XNOR2X1_25/a_35_54# XNOR2X1_25/A AOI22X1_1/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7370 XNOR2X1_25/a_12_41# XNOR2X1_25/B vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7371 gnd XNOR2X1_25/B XNOR2X1_25/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7372 vdd BUFX2_1/Y BUFX2_13/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M7373 gnd BUFX2_1/Y BUFX2_13/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M7374 BUFX2_13/Y BUFX2_13/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7375 BUFX2_13/Y BUFX2_13/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7376 vdd BUFX2_25/A BUFX2_24/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M7377 gnd BUFX2_25/A BUFX2_24/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M7378 BUFX2_24/Y BUFX2_24/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7379 BUFX2_24/Y BUFX2_24/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7380 NOR2X1_4/Y NOR2X1_4/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M7381 NOR2X1_4/Y FAX1_0/YS NOR2X1_4/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M7382 NOR2X1_4/a_9_54# NOR2X1_4/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7383 gnd FAX1_0/YS NOR2X1_4/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7384 AOI21X1_25/a_2_54# INVX2_123/Y vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M7385 AOI21X1_25/a_12_6# OR2X1_16/B gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7386 gnd AOI21X1_26/Y AOI21X1_25/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0.11n ps=52u
M7387 vdd OR2X1_16/B AOI21X1_25/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7388 AOI21X1_25/Y AOI21X1_26/Y AOI21X1_25/a_2_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7389 AOI21X1_25/Y INVX2_123/Y AOI21X1_25/a_12_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7390 AOI21X1_14/a_2_54# AOI21X1_14/B vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M7391 AOI21X1_14/a_12_6# AOI21X1_14/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7392 gnd INVX2_34/Y AOI21X1_14/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0.11n ps=52u
M7393 vdd AOI21X1_14/A AOI21X1_14/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7394 AOI21X1_14/Y INVX2_34/Y AOI21X1_14/a_2_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7395 AOI21X1_14/Y AOI21X1_14/B AOI21X1_14/a_12_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7396 vdd HAX1_39/A HAX1_39/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M7397 HAX1_39/a_41_74# HAX1_39/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M7398 HAX1_39/a_9_6# HAX1_39/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7399 HAX1_39/a_41_74# HAX1_39/B HAX1_39/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M7400 vdd HAX1_39/A HAX1_39/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7401 vdd HAX1_39/a_2_74# OR2X1_5/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M7402 HAX1_39/a_38_6# HAX1_39/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7403 MUX2X1_5/A HAX1_39/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7404 HAX1_39/a_38_6# HAX1_39/A HAX1_39/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7405 MUX2X1_5/A HAX1_39/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M7406 HAX1_39/a_2_74# HAX1_39/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7407 HAX1_39/a_2_74# HAX1_39/B HAX1_39/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7408 HAX1_39/a_49_54# HAX1_39/B HAX1_39/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7409 gnd HAX1_39/a_2_74# OR2X1_5/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M7410 vdd out_global_score[13] HAX1_17/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M7411 HAX1_17/a_41_74# HAX1_17/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M7412 HAX1_17/a_9_6# out_global_score[13] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7413 HAX1_17/a_41_74# HAX1_17/B HAX1_17/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M7414 vdd out_global_score[13] HAX1_17/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7415 vdd HAX1_17/a_2_74# HAX1_16/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M7416 HAX1_17/a_38_6# HAX1_17/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7417 HAX1_17/YS HAX1_17/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7418 HAX1_17/a_38_6# out_global_score[13] HAX1_17/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7419 HAX1_17/YS HAX1_17/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M7420 HAX1_17/a_2_74# HAX1_17/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7421 HAX1_17/a_2_74# HAX1_17/B HAX1_17/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7422 HAX1_17/a_49_54# HAX1_17/B HAX1_17/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7423 gnd HAX1_17/a_2_74# HAX1_16/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M7424 vdd out_global_score[2] HAX1_28/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M7425 HAX1_28/a_41_74# HAX1_28/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M7426 HAX1_28/a_9_6# out_global_score[2] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7427 HAX1_28/a_41_74# HAX1_28/B HAX1_28/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M7428 vdd out_global_score[2] HAX1_28/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7429 vdd HAX1_28/a_2_74# HAX1_27/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M7430 HAX1_28/a_38_6# HAX1_28/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7431 HAX1_28/YS HAX1_28/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7432 HAX1_28/a_38_6# out_global_score[2] HAX1_28/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7433 HAX1_28/YS HAX1_28/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M7434 HAX1_28/a_2_74# HAX1_28/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7435 HAX1_28/a_2_74# HAX1_28/B HAX1_28/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7436 HAX1_28/a_49_54# HAX1_28/B HAX1_28/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7437 gnd HAX1_28/a_2_74# HAX1_27/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M7438 OR2X1_1/a_2_54# OR2X1_1/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M7439 OR2X1_1/Y OR2X1_1/a_2_54# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7440 OR2X1_1/Y OR2X1_1/a_2_54# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M7441 vdd OR2X1_1/B OR2X1_1/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7442 OR2X1_1/a_9_54# OR2X1_1/A OR2X1_1/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M7443 gnd OR2X1_1/B OR2X1_1/a_2_54# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7444 gnd OAI21X1_9/A OAI21X1_9/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M7445 vdd OAI21X1_9/C OAI21X1_9/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M7446 OAI21X1_9/Y OAI21X1_9/C OAI21X1_9/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7447 OAI21X1_9/Y OAI21X1_9/B OAI21X1_9/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7448 OAI21X1_9/a_9_54# OAI21X1_9/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7449 OAI21X1_9/a_2_6# OAI21X1_9/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7450 gnd BUFX2_24/Y OAI22X1_22/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M7451 OAI22X1_22/a_2_6# OR2X1_11/A OAI22X1_22/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M7452 OAI22X1_22/Y INVX2_77/Y OAI22X1_22/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7453 OAI22X1_22/Y INVX2_107/Y OAI22X1_22/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M7454 OAI22X1_22/a_28_54# INVX2_77/Y OAI22X1_22/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7455 OAI22X1_22/a_9_54# BUFX2_24/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7456 OAI22X1_22/a_2_6# INVX2_107/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7457 vdd OR2X1_11/A OAI22X1_22/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7458 gnd BUFX2_25/Y OAI22X1_11/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M7459 OAI22X1_11/a_2_6# OAI22X1_5/C OAI22X1_11/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M7460 OAI22X1_11/Y INVX2_64/Y OAI22X1_11/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7461 OAI22X1_11/Y INVX2_96/Y OAI22X1_11/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M7462 OAI22X1_11/a_28_54# INVX2_64/Y OAI22X1_11/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7463 OAI22X1_11/a_9_54# BUFX2_25/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7464 OAI22X1_11/a_2_6# INVX2_96/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7465 vdd OAI22X1_5/C OAI22X1_11/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7466 gnd INVX2_50/Y OAI22X1_33/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M7467 OAI22X1_33/a_2_6# XOR2X1_26/Y XNOR2X1_28/B Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M7468 XNOR2X1_28/B XOR2X1_25/B OAI22X1_33/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7469 XNOR2X1_28/B INVX2_45/Y OAI22X1_33/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M7470 OAI22X1_33/a_28_54# XOR2X1_25/B XNOR2X1_28/B vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7471 OAI22X1_33/a_9_54# INVX2_50/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7472 OAI22X1_33/a_2_6# INVX2_45/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7473 vdd XOR2X1_26/Y OAI22X1_33/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7474 gnd out_mines[1] OAI22X1_66/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M7475 OAI22X1_66/a_2_6# out_mines[0] OAI22X1_66/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M7476 OAI22X1_66/Y OAI22X1_76/D OAI22X1_66/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7477 OAI22X1_66/Y OAI22X1_76/B OAI22X1_66/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M7478 OAI22X1_66/a_28_54# OAI22X1_76/D OAI22X1_66/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7479 OAI22X1_66/a_9_54# out_mines[1] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7480 OAI22X1_66/a_2_6# OAI22X1_76/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7481 vdd out_mines[0] OAI22X1_66/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7482 gnd out_mines[7] OAI22X1_55/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M7483 OAI22X1_55/a_2_6# out_mines[6] OAI22X1_55/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M7484 OAI22X1_55/Y OAI22X1_63/D OAI22X1_55/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7485 OAI22X1_55/Y OAI22X1_63/B OAI22X1_55/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M7486 OAI22X1_55/a_28_54# OAI22X1_63/D OAI22X1_55/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7487 OAI22X1_55/a_9_54# out_mines[7] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7488 OAI22X1_55/a_2_6# OAI22X1_63/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7489 vdd out_mines[6] OAI22X1_55/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7490 gnd out_mines[5] OAI22X1_44/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M7491 OAI22X1_44/a_2_6# out_mines[4] OAI22X1_44/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M7492 OAI22X1_44/Y OAI22X1_52/D OAI22X1_44/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7493 OAI22X1_44/Y OAI22X1_52/B OAI22X1_44/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M7494 OAI22X1_44/a_28_54# OAI22X1_52/D OAI22X1_44/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7495 OAI22X1_44/a_9_54# out_mines[5] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7496 OAI22X1_44/a_2_6# OAI22X1_52/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7497 vdd out_mines[4] OAI22X1_44/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7498 gnd out_mines[21] OAI22X1_88/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M7499 OAI22X1_88/a_2_6# out_mines[20] OAI22X1_88/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M7500 OAI22X1_88/Y OAI22X1_88/D OAI22X1_88/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7501 OAI22X1_88/Y OAI22X1_88/B OAI22X1_88/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M7502 OAI22X1_88/a_28_54# OAI22X1_88/D OAI22X1_88/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7503 OAI22X1_88/a_9_54# out_mines[21] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7504 OAI22X1_88/a_2_6# OAI22X1_88/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7505 vdd out_mines[20] OAI22X1_88/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7506 gnd out_mines[3] OAI22X1_77/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M7507 OAI22X1_77/a_2_6# out_mines[2] OAI22X1_77/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M7508 OAI22X1_77/Y OAI22X1_87/D OAI22X1_77/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7509 OAI22X1_77/Y OAI22X1_87/B OAI22X1_77/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M7510 OAI22X1_77/a_28_54# OAI22X1_87/D OAI22X1_77/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7511 OAI22X1_77/a_9_54# out_mines[3] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7512 OAI22X1_77/a_2_6# OAI22X1_87/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7513 vdd out_mines[2] OAI22X1_77/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7514 DFFNEGX1_7/a_76_6# BUFX2_17/Y DFFNEGX1_7/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M7515 gnd BUFX2_17/Y DFFNEGX1_7/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M7516 DFFNEGX1_7/a_66_6# DFFNEGX1_7/a_2_6# DFFNEGX1_7/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M7517 out_mines[6] DFFNEGX1_7/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7518 DFFNEGX1_7/a_23_6# BUFX2_17/Y DFFNEGX1_7/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M7519 DFFNEGX1_7/a_23_6# DFFNEGX1_7/a_2_6# DFFNEGX1_7/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M7520 gnd DFFNEGX1_7/a_34_4# DFFNEGX1_7/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M7521 vdd DFFNEGX1_7/a_34_4# DFFNEGX1_7/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M7522 DFFNEGX1_7/a_61_74# DFFNEGX1_7/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7523 DFFNEGX1_7/a_34_4# DFFNEGX1_7/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7524 DFFNEGX1_7/a_34_4# DFFNEGX1_7/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M7525 vdd out_mines[6] DFFNEGX1_7/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M7526 gnd out_mines[6] DFFNEGX1_7/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7527 DFFNEGX1_7/a_61_6# DFFNEGX1_7/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7528 DFFNEGX1_7/a_76_84# DFFNEGX1_7/a_2_6# DFFNEGX1_7/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M7529 out_mines[6] DFFNEGX1_7/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7530 vdd BUFX2_17/Y DFFNEGX1_7/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M7531 DFFNEGX1_7/a_31_6# DFFNEGX1_7/a_2_6# DFFNEGX1_7/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7532 DFFNEGX1_7/a_66_6# BUFX2_17/Y DFFNEGX1_7/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7533 DFFNEGX1_7/a_17_74# OAI21X1_39/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7534 DFFNEGX1_7/a_31_74# BUFX2_17/Y DFFNEGX1_7/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7535 DFFNEGX1_7/a_17_6# OAI21X1_39/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7536 INVX2_119/Y INVX2_119/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7537 INVX2_119/Y INVX2_119/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7538 INVX2_108/Y out_temp_cleared[5] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7539 INVX2_108/Y out_temp_cleared[5] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7540 FAX1_15/a_46_54# FAX1_15/A vdd vdd pfet w=40 l=2
+  ad=0.452n pd=0.176m as=0 ps=0
M7541 gnd FAX1_15/A FAX1_15/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M7542 gnd FAX1_15/A FAX1_15/a_84_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M7543 FAX1_15/a_33_6# FAX1_15/B FAX1_15/a_25_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.12n ps=52u
M7544 FAX1_15/a_79_6# FAX1_15/C FAX1_15/a_70_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.14n ps=54u
M7545 FAX1_15/a_46_6# FAX1_15/A gnd Gnd nfet w=20 l=2
+  ad=0.24n pd=0.104m as=0 ps=0
M7546 FAX1_14/C FAX1_15/a_70_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7547 FAX1_15/a_46_6# FAX1_15/C gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7548 FAX1_15/a_79_46# FAX1_15/C FAX1_15/a_70_6# vdd pfet w=48 l=2
+  ad=0.144n pd=0.102m as=0.317n ps=0.11m
M7549 FAX1_12/C FAX1_15/a_25_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7550 FAX1_15/a_2_54# FAX1_15/B vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M7551 FAX1_15/a_25_6# FAX1_15/C FAX1_15/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7552 gnd FAX1_15/A FAX1_15/a_33_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7553 FAX1_15/a_70_6# FAX1_15/a_25_6# FAX1_15/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M7554 FAX1_15/a_84_6# FAX1_15/B FAX1_15/a_79_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7555 vdd FAX1_15/B FAX1_15/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M7556 vdd FAX1_15/A FAX1_15/a_84_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0.144n ps=0.102m
M7557 vdd FAX1_15/A FAX1_15/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7558 FAX1_14/C FAX1_15/a_70_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M7559 FAX1_15/a_25_6# FAX1_15/C FAX1_15/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M7560 gnd FAX1_15/B FAX1_15/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7561 vdd FAX1_15/A FAX1_15/a_33_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7562 FAX1_15/a_84_46# FAX1_15/B FAX1_15/a_79_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0 ps=0
M7563 FAX1_15/a_70_6# FAX1_15/a_25_6# FAX1_15/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7564 FAX1_15/a_46_54# FAX1_15/C vdd vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M7565 FAX1_12/C FAX1_15/a_25_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M7566 FAX1_15/a_2_6# FAX1_15/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7567 FAX1_15/a_33_54# FAX1_15/B FAX1_15/a_25_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7568 NOR2X1_91/Y NOR2X1_91/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M7569 NOR2X1_91/Y NOR2X1_91/B NOR2X1_91/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M7570 NOR2X1_91/a_9_54# NOR2X1_91/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7571 gnd NOR2X1_91/B NOR2X1_91/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7572 NOR2X1_80/Y INVX2_73/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M7573 NOR2X1_80/Y INVX2_58/A NOR2X1_80/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M7574 NOR2X1_80/a_9_54# INVX2_73/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7575 gnd INVX2_58/A NOR2X1_80/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7576 gnd OAI21X1_1/B OAI21X1_109/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M7577 vdd NAND2X1_98/Y OAI21X1_109/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M7578 OAI21X1_109/Y NAND2X1_98/Y OAI21X1_109/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7579 OAI21X1_109/Y INVX2_217/Y OAI21X1_109/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7580 OAI21X1_109/a_9_54# OAI21X1_1/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7581 OAI21X1_109/a_2_6# INVX2_217/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7582 vdd BUFX2_7/A BUFX2_7/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M7583 gnd BUFX2_7/A BUFX2_7/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M7584 BUFX2_7/Y BUFX2_7/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7585 BUFX2_7/Y BUFX2_7/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7586 OAI22X1_87/B OR2X1_6/A vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M7587 NAND2X1_126/a_9_6# OR2X1_6/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7588 vdd out_temp_data_in[0] OAI22X1_87/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7589 OAI22X1_87/B out_temp_data_in[0] NAND2X1_126/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7590 OAI22X1_63/D out_temp_data_in[1] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M7591 NAND2X1_115/a_9_6# out_temp_data_in[1] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7592 vdd INVX2_251/Y OAI22X1_63/D vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7593 OAI22X1_63/D INVX2_251/Y NAND2X1_115/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7594 AOI21X1_9/A AOI22X1_63/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M7595 NAND2X1_104/a_9_6# AOI22X1_63/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7596 vdd AOI22X1_62/Y AOI21X1_9/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7597 AOI21X1_9/A AOI22X1_62/Y NAND2X1_104/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7598 FAX1_5/a_46_54# FAX1_5/A vdd vdd pfet w=40 l=2
+  ad=0.452n pd=0.176m as=0 ps=0
M7599 gnd FAX1_5/A FAX1_5/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M7600 gnd FAX1_5/A FAX1_5/a_84_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M7601 FAX1_5/a_33_6# FAX1_5/B FAX1_5/a_25_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.12n ps=52u
M7602 FAX1_5/a_79_6# FAX1_5/C FAX1_5/a_70_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.14n ps=54u
M7603 FAX1_5/a_46_6# FAX1_5/A gnd Gnd nfet w=20 l=2
+  ad=0.24n pd=0.104m as=0 ps=0
M7604 FAX1_5/YS FAX1_5/a_70_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7605 FAX1_5/a_46_6# FAX1_5/C gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7606 FAX1_5/a_79_46# FAX1_5/C FAX1_5/a_70_6# vdd pfet w=48 l=2
+  ad=0.144n pd=0.102m as=0.317n ps=0.11m
M7607 FAX1_4/C FAX1_5/a_25_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7608 FAX1_5/a_2_54# FAX1_5/B vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M7609 FAX1_5/a_25_6# FAX1_5/C FAX1_5/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7610 gnd FAX1_5/A FAX1_5/a_33_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7611 FAX1_5/a_70_6# FAX1_5/a_25_6# FAX1_5/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M7612 FAX1_5/a_84_6# FAX1_5/B FAX1_5/a_79_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7613 vdd FAX1_5/B FAX1_5/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M7614 vdd FAX1_5/A FAX1_5/a_84_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0.144n ps=0.102m
M7615 vdd FAX1_5/A FAX1_5/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7616 FAX1_5/YS FAX1_5/a_70_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M7617 FAX1_5/a_25_6# FAX1_5/C FAX1_5/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M7618 gnd FAX1_5/B FAX1_5/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7619 vdd FAX1_5/A FAX1_5/a_33_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7620 FAX1_5/a_84_46# FAX1_5/B FAX1_5/a_79_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0 ps=0
M7621 FAX1_5/a_70_6# FAX1_5/a_25_6# FAX1_5/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7622 FAX1_5/a_46_54# FAX1_5/C vdd vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M7623 FAX1_4/C FAX1_5/a_25_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M7624 FAX1_5/a_2_6# FAX1_5/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7625 FAX1_5/a_33_54# FAX1_5/B FAX1_5/a_25_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7626 HAX1_44/B NOR2X1_2/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M7627 NAND2X1_2/a_9_6# NOR2X1_2/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7628 vdd XNOR2X1_5/A HAX1_44/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7629 HAX1_44/B XNOR2X1_5/A NAND2X1_2/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7630 INVX2_7/Y out_mines[6] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7631 INVX2_7/Y out_mines[6] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7632 AOI21X1_7/a_2_54# INVX2_24/Y vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M7633 AOI21X1_7/a_12_6# AOI21X1_7/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7634 gnd AOI21X1_7/C AOI21X1_7/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0.11n ps=52u
M7635 vdd AOI21X1_7/A AOI21X1_7/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7636 AOI21X1_7/Y AOI21X1_7/C AOI21X1_7/a_2_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7637 AOI21X1_7/Y INVX2_24/Y AOI21X1_7/a_12_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7638 gnd out_temp_data_in[3] XNOR2X1_15/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M7639 INVX2_51/A out_temp_data_in[3] XNOR2X1_15/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M7640 XNOR2X1_15/a_12_41# OAI21X1_0/C gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7641 XNOR2X1_15/a_18_54# XNOR2X1_15/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7642 XNOR2X1_15/a_35_6# XNOR2X1_15/a_2_6# INVX2_51/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7643 XNOR2X1_15/a_18_6# XNOR2X1_15/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7644 vdd out_temp_data_in[3] XNOR2X1_15/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M7645 vdd OAI21X1_0/C XNOR2X1_15/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7646 INVX2_51/A XNOR2X1_15/a_2_6# XNOR2X1_15/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M7647 XNOR2X1_15/a_35_54# out_temp_data_in[3] INVX2_51/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7648 XNOR2X1_15/a_12_41# OAI21X1_0/C vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7649 gnd OAI21X1_0/C XNOR2X1_15/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7650 gnd XNOR2X1_26/A XNOR2X1_26/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M7651 NOR2X1_72/A XNOR2X1_26/A XNOR2X1_26/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M7652 XNOR2X1_26/a_12_41# XNOR2X1_26/B gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7653 XNOR2X1_26/a_18_54# XNOR2X1_26/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7654 XNOR2X1_26/a_35_6# XNOR2X1_26/a_2_6# NOR2X1_72/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7655 XNOR2X1_26/a_18_6# XNOR2X1_26/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7656 vdd XNOR2X1_26/A XNOR2X1_26/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M7657 vdd XNOR2X1_26/B XNOR2X1_26/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7658 NOR2X1_72/A XNOR2X1_26/a_2_6# XNOR2X1_26/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M7659 XNOR2X1_26/a_35_54# XNOR2X1_26/A NOR2X1_72/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7660 XNOR2X1_26/a_12_41# XNOR2X1_26/B vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7661 gnd XNOR2X1_26/B XNOR2X1_26/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7662 vdd BUFX2_25/A BUFX2_25/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M7663 gnd BUFX2_25/A BUFX2_25/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M7664 BUFX2_25/Y BUFX2_25/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7665 BUFX2_25/Y BUFX2_25/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7666 vdd BUFX2_1/Y BUFX2_14/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M7667 gnd BUFX2_1/Y BUFX2_14/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M7668 BUFX2_14/Y BUFX2_14/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7669 BUFX2_14/Y BUFX2_14/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7670 NOR2X1_5/Y NOR2X1_5/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M7671 NOR2X1_5/Y XOR2X1_9/Y NOR2X1_5/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M7672 NOR2X1_5/a_9_54# NOR2X1_5/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7673 gnd XOR2X1_9/Y NOR2X1_5/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7674 AOI21X1_26/a_2_54# NAND3X1_57/Y vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M7675 AOI21X1_26/a_12_6# AOI21X1_26/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7676 gnd AOI21X1_26/C AOI21X1_26/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0.11n ps=52u
M7677 vdd AOI21X1_26/A AOI21X1_26/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7678 AOI21X1_26/Y AOI21X1_26/C AOI21X1_26/a_2_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7679 AOI21X1_26/Y NAND3X1_57/Y AOI21X1_26/a_12_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7680 AOI21X1_15/a_2_54# AOI21X1_15/B vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M7681 AOI21X1_15/a_12_6# AOI21X1_15/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7682 gnd INVX2_39/A AOI21X1_15/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0.11n ps=52u
M7683 vdd AOI21X1_15/A AOI21X1_15/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7684 AOI21X1_15/Y INVX2_39/A AOI21X1_15/a_2_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7685 AOI21X1_15/Y AOI21X1_15/B AOI21X1_15/a_12_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7686 vdd out_global_score[12] HAX1_18/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M7687 HAX1_18/a_41_74# HAX1_18/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M7688 HAX1_18/a_9_6# out_global_score[12] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7689 HAX1_18/a_41_74# HAX1_18/B HAX1_18/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M7690 vdd out_global_score[12] HAX1_18/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7691 vdd HAX1_18/a_2_74# HAX1_17/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M7692 HAX1_18/a_38_6# HAX1_18/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7693 HAX1_18/YS HAX1_18/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7694 HAX1_18/a_38_6# out_global_score[12] HAX1_18/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7695 HAX1_18/YS HAX1_18/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M7696 HAX1_18/a_2_74# HAX1_18/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7697 HAX1_18/a_2_74# HAX1_18/B HAX1_18/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7698 HAX1_18/a_49_54# HAX1_18/B HAX1_18/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7699 gnd HAX1_18/a_2_74# HAX1_17/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M7700 vdd out_global_score[1] HAX1_29/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M7701 HAX1_29/a_41_74# HAX1_29/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M7702 HAX1_29/a_9_6# out_global_score[1] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7703 HAX1_29/a_41_74# out_global_score[0] HAX1_29/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M7704 vdd out_global_score[1] HAX1_29/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7705 vdd HAX1_29/a_2_74# HAX1_28/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M7706 HAX1_29/a_38_6# HAX1_29/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7707 HAX1_29/YS HAX1_29/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7708 HAX1_29/a_38_6# out_global_score[1] HAX1_29/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7709 HAX1_29/YS HAX1_29/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M7710 HAX1_29/a_2_74# out_global_score[0] vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7711 HAX1_29/a_2_74# out_global_score[0] HAX1_29/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7712 HAX1_29/a_49_54# out_global_score[0] HAX1_29/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7713 gnd HAX1_29/a_2_74# HAX1_28/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M7714 OR2X1_2/a_2_54# OR2X1_2/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M7715 OR2X1_2/Y OR2X1_2/a_2_54# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7716 OR2X1_2/Y OR2X1_2/a_2_54# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M7717 vdd OR2X1_2/B OR2X1_2/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7718 OR2X1_2/a_9_54# OR2X1_2/A OR2X1_2/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M7719 gnd OR2X1_2/B OR2X1_2/a_2_54# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7720 gnd BUFX2_25/Y OAI22X1_12/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M7721 OAI22X1_12/a_2_6# OR2X1_11/A OAI22X1_12/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M7722 OAI22X1_12/Y INVX2_65/Y OAI22X1_12/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7723 OAI22X1_12/Y INVX2_97/Y OAI22X1_12/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M7724 OAI22X1_12/a_28_54# INVX2_65/Y OAI22X1_12/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7725 OAI22X1_12/a_9_54# BUFX2_25/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7726 OAI22X1_12/a_2_6# INVX2_97/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7727 vdd OR2X1_11/A OAI22X1_12/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7728 gnd BUFX2_24/Y OAI22X1_23/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M7729 OAI22X1_23/a_2_6# OAI22X1_5/C OAI22X1_23/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M7730 OAI22X1_23/Y INVX2_78/Y OAI22X1_23/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7731 OAI22X1_23/Y INVX2_108/Y OAI22X1_23/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M7732 OAI22X1_23/a_28_54# INVX2_78/Y OAI22X1_23/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7733 OAI22X1_23/a_9_54# BUFX2_24/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7734 OAI22X1_23/a_2_6# INVX2_108/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7735 vdd OAI22X1_5/C OAI22X1_23/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7736 gnd out_temp_data_in[1] OAI22X1_34/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M7737 OAI22X1_34/a_2_6# OAI22X1_34/C INVX2_44/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M7738 INVX2_44/A OR2X1_6/A OAI22X1_34/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7739 INVX2_44/A INVX2_43/Y OAI22X1_34/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M7740 OAI22X1_34/a_28_54# OR2X1_6/A INVX2_44/A vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7741 OAI22X1_34/a_9_54# out_temp_data_in[1] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7742 OAI22X1_34/a_2_6# INVX2_43/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7743 vdd OAI22X1_34/C OAI22X1_34/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7744 gnd out_mines[11] OAI22X1_45/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M7745 OAI22X1_45/a_2_6# out_mines[10] OAI22X1_45/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M7746 OAI22X1_45/Y OAI22X1_51/D OAI22X1_45/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7747 OAI22X1_45/Y OAI22X1_51/B OAI22X1_45/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M7748 OAI22X1_45/a_28_54# OAI22X1_51/D OAI22X1_45/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7749 OAI22X1_45/a_9_54# out_mines[11] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7750 OAI22X1_45/a_2_6# OAI22X1_51/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7751 vdd out_mines[10] OAI22X1_45/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7752 gnd out_mines[5] OAI22X1_56/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M7753 OAI22X1_56/a_2_6# out_mines[4] OAI22X1_56/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M7754 OAI22X1_56/Y OAI22X1_64/D OAI22X1_56/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7755 OAI22X1_56/Y OAI22X1_64/B OAI22X1_56/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M7756 OAI22X1_56/a_28_54# OAI22X1_64/D OAI22X1_56/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7757 OAI22X1_56/a_9_54# out_mines[5] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7758 OAI22X1_56/a_2_6# OAI22X1_64/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7759 vdd out_mines[4] OAI22X1_56/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7760 gnd out_mines[7] OAI22X1_67/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M7761 OAI22X1_67/a_2_6# out_mines[6] OAI22X1_67/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M7762 OAI22X1_67/Y OAI22X1_75/D OAI22X1_67/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7763 OAI22X1_67/Y OAI22X1_75/B OAI22X1_67/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M7764 OAI22X1_67/a_28_54# OAI22X1_75/D OAI22X1_67/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7765 OAI22X1_67/a_9_54# out_mines[7] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7766 OAI22X1_67/a_2_6# OAI22X1_75/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7767 vdd out_mines[6] OAI22X1_67/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7768 gnd out_mines[1] OAI22X1_78/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M7769 OAI22X1_78/a_2_6# out_mines[0] OAI22X1_78/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M7770 OAI22X1_78/Y OAI22X1_88/D OAI22X1_78/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7771 OAI22X1_78/Y OAI22X1_88/B OAI22X1_78/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M7772 OAI22X1_78/a_28_54# OAI22X1_88/D OAI22X1_78/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7773 OAI22X1_78/a_9_54# out_mines[1] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7774 OAI22X1_78/a_2_6# OAI22X1_88/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7775 vdd out_mines[0] OAI22X1_78/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7776 DFFNEGX1_8/a_76_6# BUFX2_17/Y DFFNEGX1_8/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M7777 gnd BUFX2_17/Y DFFNEGX1_8/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M7778 DFFNEGX1_8/a_66_6# DFFNEGX1_8/a_2_6# DFFNEGX1_8/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M7779 out_mines[4] DFFNEGX1_8/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7780 DFFNEGX1_8/a_23_6# BUFX2_17/Y DFFNEGX1_8/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M7781 DFFNEGX1_8/a_23_6# DFFNEGX1_8/a_2_6# DFFNEGX1_8/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M7782 gnd DFFNEGX1_8/a_34_4# DFFNEGX1_8/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M7783 vdd DFFNEGX1_8/a_34_4# DFFNEGX1_8/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M7784 DFFNEGX1_8/a_61_74# DFFNEGX1_8/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7785 DFFNEGX1_8/a_34_4# DFFNEGX1_8/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7786 DFFNEGX1_8/a_34_4# DFFNEGX1_8/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M7787 vdd out_mines[4] DFFNEGX1_8/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M7788 gnd out_mines[4] DFFNEGX1_8/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7789 DFFNEGX1_8/a_61_6# DFFNEGX1_8/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7790 DFFNEGX1_8/a_76_84# DFFNEGX1_8/a_2_6# DFFNEGX1_8/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M7791 out_mines[4] DFFNEGX1_8/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7792 vdd BUFX2_17/Y DFFNEGX1_8/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M7793 DFFNEGX1_8/a_31_6# DFFNEGX1_8/a_2_6# DFFNEGX1_8/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7794 DFFNEGX1_8/a_66_6# BUFX2_17/Y DFFNEGX1_8/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7795 DFFNEGX1_8/a_17_74# OAI21X1_43/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7796 DFFNEGX1_8/a_31_74# BUFX2_17/Y DFFNEGX1_8/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7797 DFFNEGX1_8/a_17_6# OAI21X1_43/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7798 OAI22X1_2/B out_temp_cleared[4] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7799 OAI22X1_2/B out_temp_cleared[4] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7800 FAX1_16/a_46_54# FAX1_16/A vdd vdd pfet w=40 l=2
+  ad=0.452n pd=0.176m as=0 ps=0
M7801 gnd FAX1_16/A FAX1_16/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M7802 gnd FAX1_16/A FAX1_16/a_84_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M7803 FAX1_16/a_33_6# FAX1_16/B FAX1_16/a_25_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.12n ps=52u
M7804 FAX1_16/a_79_6# FAX1_16/C FAX1_16/a_70_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.14n ps=54u
M7805 FAX1_16/a_46_6# FAX1_16/A gnd Gnd nfet w=20 l=2
+  ad=0.24n pd=0.104m as=0 ps=0
M7806 FAX1_8/B FAX1_16/a_70_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7807 FAX1_16/a_46_6# FAX1_16/C gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7808 FAX1_16/a_79_46# FAX1_16/C FAX1_16/a_70_6# vdd pfet w=48 l=2
+  ad=0.144n pd=0.102m as=0.317n ps=0.11m
M7809 FAX1_7/A FAX1_16/a_25_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7810 FAX1_16/a_2_54# FAX1_16/B vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M7811 FAX1_16/a_25_6# FAX1_16/C FAX1_16/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7812 gnd FAX1_16/A FAX1_16/a_33_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7813 FAX1_16/a_70_6# FAX1_16/a_25_6# FAX1_16/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M7814 FAX1_16/a_84_6# FAX1_16/B FAX1_16/a_79_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7815 vdd FAX1_16/B FAX1_16/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M7816 vdd FAX1_16/A FAX1_16/a_84_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0.144n ps=0.102m
M7817 vdd FAX1_16/A FAX1_16/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7818 FAX1_8/B FAX1_16/a_70_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M7819 FAX1_16/a_25_6# FAX1_16/C FAX1_16/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M7820 gnd FAX1_16/B FAX1_16/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7821 vdd FAX1_16/A FAX1_16/a_33_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7822 FAX1_16/a_84_46# FAX1_16/B FAX1_16/a_79_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0 ps=0
M7823 FAX1_16/a_70_6# FAX1_16/a_25_6# FAX1_16/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7824 FAX1_16/a_46_54# FAX1_16/C vdd vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M7825 FAX1_7/A FAX1_16/a_25_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M7826 FAX1_16/a_2_6# FAX1_16/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7827 FAX1_16/a_33_54# FAX1_16/B FAX1_16/a_25_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7828 NOR2X1_81/Y NOR2X1_86/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M7829 NOR2X1_81/Y NOR2X1_84/A NOR2X1_81/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M7830 NOR2X1_81/a_9_54# NOR2X1_86/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7831 gnd NOR2X1_84/A NOR2X1_81/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7832 NOR2X1_70/Y out_start gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M7833 NOR2X1_70/Y out_display NOR2X1_70/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M7834 NOR2X1_70/a_9_54# out_start vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7835 gnd out_display NOR2X1_70/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7836 NOR2X1_92/Y out_temp_decoded[23] gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M7837 NOR2X1_92/Y out_temp_cleared[23] NOR2X1_92/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M7838 NOR2X1_92/a_9_54# out_temp_decoded[23] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7839 gnd out_temp_cleared[23] NOR2X1_92/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7840 vdd BUFX2_8/A BUFX2_8/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M7841 gnd BUFX2_8/A BUFX2_8/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M7842 BUFX2_8/Y BUFX2_8/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7843 BUFX2_8/Y BUFX2_8/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7844 OAI22X1_63/B out_temp_data_in[1] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M7845 NAND2X1_116/a_9_6# out_temp_data_in[1] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7846 vdd out_temp_data_in[0] OAI22X1_63/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7847 OAI22X1_63/B out_temp_data_in[0] NAND2X1_116/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7848 INVX2_47/A AOI22X1_65/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M7849 NAND2X1_105/a_9_6# AOI22X1_65/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7850 vdd AOI22X1_64/Y INVX2_47/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7851 INVX2_47/A AOI22X1_64/Y NAND2X1_105/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7852 FAX1_6/a_46_54# FAX1_6/A vdd vdd pfet w=40 l=2
+  ad=0.452n pd=0.176m as=0 ps=0
M7853 gnd FAX1_6/A FAX1_6/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M7854 gnd FAX1_6/A FAX1_6/a_84_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M7855 FAX1_6/a_33_6# FAX1_6/B FAX1_6/a_25_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.12n ps=52u
M7856 FAX1_6/a_79_6# FAX1_6/C FAX1_6/a_70_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.14n ps=54u
M7857 FAX1_6/a_46_6# FAX1_6/A gnd Gnd nfet w=20 l=2
+  ad=0.24n pd=0.104m as=0 ps=0
M7858 FAX1_6/YS FAX1_6/a_70_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7859 FAX1_6/a_46_6# FAX1_6/C gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7860 FAX1_6/a_79_46# FAX1_6/C FAX1_6/a_70_6# vdd pfet w=48 l=2
+  ad=0.144n pd=0.102m as=0.317n ps=0.11m
M7861 FAX1_5/C FAX1_6/a_25_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7862 FAX1_6/a_2_54# FAX1_6/B vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M7863 FAX1_6/a_25_6# FAX1_6/C FAX1_6/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7864 gnd FAX1_6/A FAX1_6/a_33_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7865 FAX1_6/a_70_6# FAX1_6/a_25_6# FAX1_6/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M7866 FAX1_6/a_84_6# FAX1_6/B FAX1_6/a_79_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7867 vdd FAX1_6/B FAX1_6/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M7868 vdd FAX1_6/A FAX1_6/a_84_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0.144n ps=0.102m
M7869 vdd FAX1_6/A FAX1_6/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7870 FAX1_6/YS FAX1_6/a_70_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M7871 FAX1_6/a_25_6# FAX1_6/C FAX1_6/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M7872 gnd FAX1_6/B FAX1_6/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7873 vdd FAX1_6/A FAX1_6/a_33_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7874 FAX1_6/a_84_46# FAX1_6/B FAX1_6/a_79_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0 ps=0
M7875 FAX1_6/a_70_6# FAX1_6/a_25_6# FAX1_6/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7876 FAX1_6/a_46_54# FAX1_6/C vdd vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M7877 FAX1_5/C FAX1_6/a_25_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M7878 FAX1_6/a_2_6# FAX1_6/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7879 FAX1_6/a_33_54# FAX1_6/B FAX1_6/a_25_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7880 OAI22X1_88/D INVX2_251/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M7881 NAND2X1_127/a_9_6# INVX2_251/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7882 vdd out_temp_data_in[1] OAI22X1_88/D vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7883 OAI22X1_88/D out_temp_data_in[1] NAND2X1_127/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7884 HAX1_42/B NOR2X1_3/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M7885 NAND2X1_3/a_9_6# NOR2X1_3/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7886 vdd XNOR2X1_7/A HAX1_42/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7887 HAX1_42/B XNOR2X1_7/A NAND2X1_3/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7888 INVX2_8/Y out_mines[4] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7889 INVX2_8/Y out_mines[4] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7890 AOI21X1_8/a_2_54# AOI21X1_8/B vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M7891 AOI21X1_8/a_12_6# INVX2_251/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7892 gnd AOI21X1_8/C INVX2_42/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0.11n ps=52u
M7893 vdd INVX2_251/Y AOI21X1_8/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7894 INVX2_42/A AOI21X1_8/C AOI21X1_8/a_2_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7895 INVX2_42/A AOI21X1_8/B AOI21X1_8/a_12_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7896 gnd out_temp_data_in[2] XNOR2X1_16/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M7897 INVX2_34/A out_temp_data_in[2] XNOR2X1_16/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M7898 XNOR2X1_16/a_12_41# out_temp_data_in[3] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7899 XNOR2X1_16/a_18_54# XNOR2X1_16/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7900 XNOR2X1_16/a_35_6# XNOR2X1_16/a_2_6# INVX2_34/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7901 XNOR2X1_16/a_18_6# XNOR2X1_16/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7902 vdd out_temp_data_in[2] XNOR2X1_16/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M7903 vdd out_temp_data_in[3] XNOR2X1_16/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7904 INVX2_34/A XNOR2X1_16/a_2_6# XNOR2X1_16/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M7905 XNOR2X1_16/a_35_54# out_temp_data_in[2] INVX2_34/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7906 XNOR2X1_16/a_12_41# out_temp_data_in[3] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7907 gnd out_temp_data_in[3] XNOR2X1_16/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7908 gnd XNOR2X1_27/A XNOR2X1_27/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M7909 XOR2X1_23/B XNOR2X1_27/A XNOR2X1_27/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M7910 XNOR2X1_27/a_12_41# XNOR2X1_27/B gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7911 XNOR2X1_27/a_18_54# XNOR2X1_27/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7912 XNOR2X1_27/a_35_6# XNOR2X1_27/a_2_6# XOR2X1_23/B Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7913 XNOR2X1_27/a_18_6# XNOR2X1_27/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7914 vdd XNOR2X1_27/A XNOR2X1_27/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M7915 vdd XNOR2X1_27/B XNOR2X1_27/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7916 XOR2X1_23/B XNOR2X1_27/a_2_6# XNOR2X1_27/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M7917 XNOR2X1_27/a_35_54# XNOR2X1_27/A XOR2X1_23/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7918 XNOR2X1_27/a_12_41# XNOR2X1_27/B vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7919 gnd XNOR2X1_27/B XNOR2X1_27/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7920 vdd BUFX2_2/Y BUFX2_15/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M7921 gnd BUFX2_2/Y BUFX2_15/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M7922 BUFX2_15/Y BUFX2_15/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7923 BUFX2_15/Y BUFX2_15/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7924 NOR2X1_6/Y XOR2X1_8/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M7925 NOR2X1_6/Y XOR2X1_7/Y NOR2X1_6/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M7926 NOR2X1_6/a_9_54# XOR2X1_8/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7927 gnd XOR2X1_7/Y NOR2X1_6/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7928 AOI21X1_16/a_2_54# AOI21X1_16/B vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M7929 AOI21X1_16/a_12_6# AOI21X1_16/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7930 gnd INVX2_39/Y AOI21X1_16/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0.11n ps=52u
M7931 vdd AOI21X1_16/A AOI21X1_16/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7932 AOI21X1_16/Y INVX2_39/Y AOI21X1_16/a_2_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M7933 AOI21X1_16/Y AOI21X1_16/B AOI21X1_16/a_12_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7934 vdd out_global_score[11] HAX1_19/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M7935 HAX1_19/a_41_74# HAX1_19/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M7936 HAX1_19/a_9_6# out_global_score[11] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M7937 HAX1_19/a_41_74# HAX1_19/B HAX1_19/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M7938 vdd out_global_score[11] HAX1_19/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7939 vdd HAX1_19/a_2_74# HAX1_18/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M7940 HAX1_19/a_38_6# HAX1_19/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7941 HAX1_19/YS HAX1_19/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7942 HAX1_19/a_38_6# out_global_score[11] HAX1_19/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7943 HAX1_19/YS HAX1_19/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M7944 HAX1_19/a_2_74# HAX1_19/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7945 HAX1_19/a_2_74# HAX1_19/B HAX1_19/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7946 HAX1_19/a_49_54# HAX1_19/B HAX1_19/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7947 gnd HAX1_19/a_2_74# HAX1_18/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M7948 OR2X1_3/a_2_54# OR2X1_3/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M7949 OR2X1_3/Y OR2X1_3/a_2_54# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M7950 OR2X1_3/Y OR2X1_3/a_2_54# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M7951 vdd OR2X1_3/B OR2X1_3/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M7952 OR2X1_3/a_9_54# OR2X1_3/A OR2X1_3/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M7953 gnd OR2X1_3/B OR2X1_3/a_2_54# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M7954 gnd BUFX2_25/Y OAI22X1_13/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M7955 OAI22X1_13/a_2_6# OAI22X1_5/C OAI22X1_13/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M7956 OAI22X1_13/Y INVX2_66/Y OAI22X1_13/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7957 OAI22X1_13/Y INVX2_98/Y OAI22X1_13/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M7958 OAI22X1_13/a_28_54# INVX2_66/Y OAI22X1_13/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7959 OAI22X1_13/a_9_54# BUFX2_25/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7960 OAI22X1_13/a_2_6# INVX2_98/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7961 vdd OAI22X1_5/C OAI22X1_13/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7962 gnd BUFX2_24/Y OAI22X1_24/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M7963 OAI22X1_24/a_2_6# OR2X1_11/A OAI22X1_24/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M7964 OAI22X1_24/Y INVX2_79/Y OAI22X1_24/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7965 OAI22X1_24/Y OAI22X1_2/B OAI22X1_24/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M7966 OAI22X1_24/a_28_54# INVX2_79/Y OAI22X1_24/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7967 OAI22X1_24/a_9_54# BUFX2_24/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7968 OAI22X1_24/a_2_6# OAI22X1_2/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7969 vdd OR2X1_11/A OAI22X1_24/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7970 gnd out_mines[9] OAI22X1_46/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M7971 OAI22X1_46/a_2_6# out_mines[8] OAI22X1_46/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M7972 OAI22X1_46/Y OAI22X1_52/D OAI22X1_46/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7973 OAI22X1_46/Y OAI22X1_52/B OAI22X1_46/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M7974 OAI22X1_46/a_28_54# OAI22X1_52/D OAI22X1_46/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7975 OAI22X1_46/a_9_54# out_mines[9] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7976 OAI22X1_46/a_2_6# OAI22X1_52/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7977 vdd out_mines[8] OAI22X1_46/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7978 gnd INVX2_21/Y OAI22X1_35/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M7979 OAI22X1_35/a_2_6# INVX2_14/Y OAI22X1_35/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M7980 OAI22X1_35/Y INVX2_32/A OAI22X1_35/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7981 OAI22X1_35/Y INVX2_31/A OAI22X1_35/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M7982 OAI22X1_35/a_28_54# INVX2_32/A OAI22X1_35/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7983 OAI22X1_35/a_9_54# INVX2_21/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7984 OAI22X1_35/a_2_6# INVX2_31/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7985 vdd INVX2_14/Y OAI22X1_35/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7986 gnd out_mines[11] OAI22X1_57/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M7987 OAI22X1_57/a_2_6# out_mines[10] OAI22X1_57/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M7988 OAI22X1_57/Y OAI22X1_63/D OAI22X1_57/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7989 OAI22X1_57/Y OAI22X1_63/B OAI22X1_57/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M7990 OAI22X1_57/a_28_54# OAI22X1_63/D OAI22X1_57/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7991 OAI22X1_57/a_9_54# out_mines[11] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7992 OAI22X1_57/a_2_6# OAI22X1_63/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7993 vdd out_mines[10] OAI22X1_57/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M7994 gnd out_mines[7] OAI22X1_79/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M7995 OAI22X1_79/a_2_6# out_mines[6] OAI22X1_79/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M7996 OAI22X1_79/Y OAI22X1_87/D OAI22X1_79/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M7997 OAI22X1_79/Y OAI22X1_87/B OAI22X1_79/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M7998 OAI22X1_79/a_28_54# OAI22X1_87/D OAI22X1_79/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M7999 OAI22X1_79/a_9_54# out_mines[7] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8000 OAI22X1_79/a_2_6# OAI22X1_87/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8001 vdd out_mines[6] OAI22X1_79/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8002 gnd out_mines[5] OAI22X1_68/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M8003 OAI22X1_68/a_2_6# out_mines[4] OAI22X1_68/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M8004 OAI22X1_68/Y OAI22X1_76/D OAI22X1_68/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8005 OAI22X1_68/Y OAI22X1_76/B OAI22X1_68/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M8006 OAI22X1_68/a_28_54# OAI22X1_76/D OAI22X1_68/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M8007 OAI22X1_68/a_9_54# out_mines[5] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8008 OAI22X1_68/a_2_6# OAI22X1_76/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8009 vdd out_mines[4] OAI22X1_68/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8010 DFFNEGX1_9/a_76_6# BUFX2_17/Y DFFNEGX1_9/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M8011 gnd BUFX2_17/Y DFFNEGX1_9/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M8012 DFFNEGX1_9/a_66_6# DFFNEGX1_9/a_2_6# DFFNEGX1_9/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M8013 out_mines[0] DFFNEGX1_9/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8014 DFFNEGX1_9/a_23_6# BUFX2_17/Y DFFNEGX1_9/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M8015 DFFNEGX1_9/a_23_6# DFFNEGX1_9/a_2_6# DFFNEGX1_9/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M8016 gnd DFFNEGX1_9/a_34_4# DFFNEGX1_9/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M8017 vdd DFFNEGX1_9/a_34_4# DFFNEGX1_9/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M8018 DFFNEGX1_9/a_61_74# DFFNEGX1_9/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M8019 DFFNEGX1_9/a_34_4# DFFNEGX1_9/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8020 DFFNEGX1_9/a_34_4# DFFNEGX1_9/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M8021 vdd out_mines[0] DFFNEGX1_9/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M8022 gnd out_mines[0] DFFNEGX1_9/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8023 DFFNEGX1_9/a_61_6# DFFNEGX1_9/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8024 DFFNEGX1_9/a_76_84# DFFNEGX1_9/a_2_6# DFFNEGX1_9/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M8025 out_mines[0] DFFNEGX1_9/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M8026 vdd BUFX2_17/Y DFFNEGX1_9/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M8027 DFFNEGX1_9/a_31_6# DFFNEGX1_9/a_2_6# DFFNEGX1_9/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8028 DFFNEGX1_9/a_66_6# BUFX2_17/Y DFFNEGX1_9/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8029 DFFNEGX1_9/a_17_74# OAI21X1_51/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8030 DFFNEGX1_9/a_31_74# BUFX2_17/Y DFFNEGX1_9/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8031 DFFNEGX1_9/a_17_6# OAI21X1_51/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8032 gnd INVX2_74/Y OAI21X1_90/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M8033 vdd OAI21X1_90/C OAI21X1_90/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M8034 OAI21X1_90/Y OAI21X1_90/C OAI21X1_90/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8035 OAI21X1_90/Y BUFX2_22/Y OAI21X1_90/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8036 OAI21X1_90/a_9_54# INVX2_74/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8037 OAI21X1_90/a_2_6# BUFX2_22/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8038 FAX1_17/a_46_54# FAX1_17/A vdd vdd pfet w=40 l=2
+  ad=0.452n pd=0.176m as=0 ps=0
M8039 gnd FAX1_17/A FAX1_17/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M8040 gnd FAX1_17/A FAX1_17/a_84_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M8041 FAX1_17/a_33_6# FAX1_17/B FAX1_17/a_25_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.12n ps=52u
M8042 FAX1_17/a_79_6# FAX1_17/C FAX1_17/a_70_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.14n ps=54u
M8043 FAX1_17/a_46_6# FAX1_17/A gnd Gnd nfet w=20 l=2
+  ad=0.24n pd=0.104m as=0 ps=0
M8044 FAX1_16/C FAX1_17/a_70_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8045 FAX1_17/a_46_6# FAX1_17/C gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8046 FAX1_17/a_79_46# FAX1_17/C FAX1_17/a_70_6# vdd pfet w=48 l=2
+  ad=0.144n pd=0.102m as=0.317n ps=0.11m
M8047 FAX1_14/B FAX1_17/a_25_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8048 FAX1_17/a_2_54# FAX1_17/B vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M8049 FAX1_17/a_25_6# FAX1_17/C FAX1_17/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8050 gnd FAX1_17/A FAX1_17/a_33_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8051 FAX1_17/a_70_6# FAX1_17/a_25_6# FAX1_17/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M8052 FAX1_17/a_84_6# FAX1_17/B FAX1_17/a_79_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8053 vdd FAX1_17/B FAX1_17/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M8054 vdd FAX1_17/A FAX1_17/a_84_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0.144n ps=0.102m
M8055 vdd FAX1_17/A FAX1_17/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8056 FAX1_16/C FAX1_17/a_70_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M8057 FAX1_17/a_25_6# FAX1_17/C FAX1_17/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M8058 gnd FAX1_17/B FAX1_17/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8059 vdd FAX1_17/A FAX1_17/a_33_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8060 FAX1_17/a_84_46# FAX1_17/B FAX1_17/a_79_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0 ps=0
M8061 FAX1_17/a_70_6# FAX1_17/a_25_6# FAX1_17/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8062 FAX1_17/a_46_54# FAX1_17/C vdd vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M8063 FAX1_14/B FAX1_17/a_25_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M8064 FAX1_17/a_2_6# FAX1_17/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8065 FAX1_17/a_33_54# FAX1_17/B FAX1_17/a_25_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8066 NOR2X1_82/Y NOR2X1_82/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8067 NOR2X1_82/Y NOR2X1_82/B NOR2X1_82/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8068 NOR2X1_82/a_9_54# NOR2X1_82/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8069 gnd NOR2X1_82/B NOR2X1_82/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8070 INVX2_54/A out_temp_data_in[0] gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8071 INVX2_54/A out_temp_data_in[1] NOR2X1_60/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8072 NOR2X1_60/a_9_54# out_temp_data_in[0] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8073 gnd out_temp_data_in[1] INVX2_54/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8074 NOR2X1_71/Y NOR2X1_73/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8075 NOR2X1_71/Y NOR2X1_71/B NOR2X1_71/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8076 NOR2X1_71/a_9_54# NOR2X1_73/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8077 gnd NOR2X1_71/B NOR2X1_71/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8078 NOR2X1_93/Y out_temp_decoded[14] gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8079 NOR2X1_93/Y out_temp_cleared[14] NOR2X1_93/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8080 NOR2X1_93/a_9_54# out_temp_decoded[14] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8081 gnd out_temp_cleared[14] NOR2X1_93/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8082 vdd BUFX2_9/A BUFX2_9/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M8083 gnd BUFX2_9/A BUFX2_9/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M8084 BUFX2_9/Y BUFX2_9/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M8085 BUFX2_9/Y BUFX2_9/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8086 INVX2_31/A out_temp_data_in[3] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M8087 NAND2X1_106/a_9_6# out_temp_data_in[3] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M8088 vdd INVX2_30/Y INVX2_31/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8089 INVX2_31/A INVX2_30/Y NAND2X1_106/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8090 OAI22X1_64/D INVX2_251/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M8091 NAND2X1_117/a_9_6# INVX2_251/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M8092 vdd OR2X1_6/A OAI22X1_64/D vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8093 OAI22X1_64/D OR2X1_6/A NAND2X1_117/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8094 FAX1_7/a_46_54# FAX1_7/A vdd vdd pfet w=40 l=2
+  ad=0.452n pd=0.176m as=0 ps=0
M8095 gnd FAX1_7/A FAX1_7/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M8096 gnd FAX1_7/A FAX1_7/a_84_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M8097 FAX1_7/a_33_6# FAX1_7/B FAX1_7/a_25_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.12n ps=52u
M8098 FAX1_7/a_79_6# FAX1_7/C FAX1_7/a_70_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.14n ps=54u
M8099 FAX1_7/a_46_6# FAX1_7/A gnd Gnd nfet w=20 l=2
+  ad=0.24n pd=0.104m as=0 ps=0
M8100 FAX1_7/YS FAX1_7/a_70_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8101 FAX1_7/a_46_6# FAX1_7/C gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8102 FAX1_7/a_79_46# FAX1_7/C FAX1_7/a_70_6# vdd pfet w=48 l=2
+  ad=0.144n pd=0.102m as=0.317n ps=0.11m
M8103 FAX1_6/C FAX1_7/a_25_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8104 FAX1_7/a_2_54# FAX1_7/B vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M8105 FAX1_7/a_25_6# FAX1_7/C FAX1_7/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8106 gnd FAX1_7/A FAX1_7/a_33_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8107 FAX1_7/a_70_6# FAX1_7/a_25_6# FAX1_7/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M8108 FAX1_7/a_84_6# FAX1_7/B FAX1_7/a_79_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8109 vdd FAX1_7/B FAX1_7/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M8110 vdd FAX1_7/A FAX1_7/a_84_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0.144n ps=0.102m
M8111 vdd FAX1_7/A FAX1_7/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8112 FAX1_7/YS FAX1_7/a_70_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M8113 FAX1_7/a_25_6# FAX1_7/C FAX1_7/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M8114 gnd FAX1_7/B FAX1_7/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8115 vdd FAX1_7/A FAX1_7/a_33_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8116 FAX1_7/a_84_46# FAX1_7/B FAX1_7/a_79_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0 ps=0
M8117 FAX1_7/a_70_6# FAX1_7/a_25_6# FAX1_7/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8118 FAX1_7/a_46_54# FAX1_7/C vdd vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M8119 FAX1_6/C FAX1_7/a_25_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M8120 FAX1_7/a_2_6# FAX1_7/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8121 FAX1_7/a_33_54# FAX1_7/B FAX1_7/a_25_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8122 OAI22X1_88/B out_temp_data_in[0] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M8123 NAND2X1_128/a_9_6# out_temp_data_in[0] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M8124 vdd out_temp_data_in[1] OAI22X1_88/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8125 OAI22X1_88/B out_temp_data_in[1] NAND2X1_128/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8126 HAX1_40/B NOR2X1_4/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M8127 NAND2X1_4/a_9_6# NOR2X1_4/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M8128 vdd MUX2X1_8/Y HAX1_40/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8129 HAX1_40/B MUX2X1_8/Y NAND2X1_4/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8130 INVX2_9/Y out_mines[0] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8131 INVX2_9/Y out_mines[0] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M8132 AOI21X1_9/a_2_54# INVX2_31/Y vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M8133 AOI21X1_9/a_12_6# AOI21X1_9/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M8134 gnd AOI21X1_9/C INVX2_46/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0.11n ps=52u
M8135 vdd AOI21X1_9/A AOI21X1_9/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8136 INVX2_46/A AOI21X1_9/C AOI21X1_9/a_2_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M8137 INVX2_46/A INVX2_31/Y AOI21X1_9/a_12_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8138 gnd OR2X1_8/B XNOR2X1_17/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M8139 INVX2_39/A OR2X1_8/B XNOR2X1_17/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M8140 XNOR2X1_17/a_12_41# out_temp_data_in[3] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8141 XNOR2X1_17/a_18_54# XNOR2X1_17/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M8142 XNOR2X1_17/a_35_6# XNOR2X1_17/a_2_6# INVX2_39/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M8143 XNOR2X1_17/a_18_6# XNOR2X1_17/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8144 vdd OR2X1_8/B XNOR2X1_17/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M8145 vdd out_temp_data_in[3] XNOR2X1_17/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8146 INVX2_39/A XNOR2X1_17/a_2_6# XNOR2X1_17/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M8147 XNOR2X1_17/a_35_54# OR2X1_8/B INVX2_39/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8148 XNOR2X1_17/a_12_41# out_temp_data_in[3] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M8149 gnd out_temp_data_in[3] XNOR2X1_17/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8150 gnd XNOR2X1_28/A XNOR2X1_28/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M8151 XOR2X1_23/A XNOR2X1_28/A XNOR2X1_28/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M8152 XNOR2X1_28/a_12_41# XNOR2X1_28/B gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8153 XNOR2X1_28/a_18_54# XNOR2X1_28/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M8154 XNOR2X1_28/a_35_6# XNOR2X1_28/a_2_6# XOR2X1_23/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M8155 XNOR2X1_28/a_18_6# XNOR2X1_28/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8156 vdd XNOR2X1_28/A XNOR2X1_28/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M8157 vdd XNOR2X1_28/B XNOR2X1_28/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8158 XOR2X1_23/A XNOR2X1_28/a_2_6# XNOR2X1_28/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M8159 XNOR2X1_28/a_35_54# XNOR2X1_28/A XOR2X1_23/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8160 XNOR2X1_28/a_12_41# XNOR2X1_28/B vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M8161 gnd XNOR2X1_28/B XNOR2X1_28/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8162 vdd BUFX2_2/Y BUFX2_16/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M8163 gnd BUFX2_2/Y BUFX2_16/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M8164 BUFX2_16/Y BUFX2_16/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M8165 BUFX2_16/Y BUFX2_16/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8166 NOR2X1_7/Y NOR2X1_7/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8167 NOR2X1_7/Y NOR2X1_7/B NOR2X1_7/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8168 NOR2X1_7/a_9_54# NOR2X1_7/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8169 gnd NOR2X1_7/B NOR2X1_7/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8170 AOI21X1_17/a_2_54# AOI21X1_17/B vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M8171 AOI21X1_17/a_12_6# AOI21X1_17/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M8172 gnd INVX2_36/A AOI21X1_17/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0.11n ps=52u
M8173 vdd AOI21X1_17/A AOI21X1_17/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8174 AOI21X1_17/Y INVX2_36/A AOI21X1_17/a_2_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M8175 AOI21X1_17/Y AOI21X1_17/B AOI21X1_17/a_12_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8176 OR2X1_4/a_2_54# OR2X1_4/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8177 OR2X1_4/Y OR2X1_4/a_2_54# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8178 OR2X1_4/Y OR2X1_4/a_2_54# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M8179 vdd OR2X1_4/B OR2X1_4/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8180 OR2X1_4/a_9_54# OR2X1_4/A OR2X1_4/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M8181 gnd OR2X1_4/B OR2X1_4/a_2_54# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8182 gnd BUFX2_25/Y OAI22X1_14/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M8183 OAI22X1_14/a_2_6# OR2X1_11/A OAI22X1_14/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M8184 OAI22X1_14/Y INVX2_67/Y OAI22X1_14/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8185 OAI22X1_14/Y INVX2_99/Y OAI22X1_14/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M8186 OAI22X1_14/a_28_54# INVX2_67/Y OAI22X1_14/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M8187 OAI22X1_14/a_9_54# BUFX2_25/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8188 OAI22X1_14/a_2_6# INVX2_99/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8189 vdd OR2X1_11/A OAI22X1_14/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8190 gnd BUFX2_24/Y OAI22X1_25/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M8191 OAI22X1_25/a_2_6# OAI22X1_5/C OAI22X1_25/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M8192 OAI22X1_25/Y INVX2_81/Y OAI22X1_25/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8193 OAI22X1_25/Y OAI22X1_2/D OAI22X1_25/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M8194 OAI22X1_25/a_28_54# INVX2_81/Y OAI22X1_25/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M8195 OAI22X1_25/a_9_54# BUFX2_24/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8196 OAI22X1_25/a_2_6# OAI22X1_2/D gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8197 vdd OAI22X1_5/C OAI22X1_25/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8198 gnd out_mines[15] OAI22X1_47/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M8199 OAI22X1_47/a_2_6# out_mines[14] OAI22X1_47/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M8200 OAI22X1_47/Y OAI22X1_51/D OAI22X1_47/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8201 OAI22X1_47/Y OAI22X1_51/B OAI22X1_47/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M8202 OAI22X1_47/a_28_54# OAI22X1_51/D OAI22X1_47/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M8203 OAI22X1_47/a_9_54# out_mines[15] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8204 OAI22X1_47/a_2_6# OAI22X1_51/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8205 vdd out_mines[14] OAI22X1_47/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8206 gnd out_mines[9] OAI22X1_58/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M8207 OAI22X1_58/a_2_6# out_mines[8] OAI22X1_58/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M8208 OAI22X1_58/Y OAI22X1_64/D OAI22X1_58/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8209 OAI22X1_58/Y OAI22X1_64/B OAI22X1_58/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M8210 OAI22X1_58/a_28_54# OAI22X1_64/D OAI22X1_58/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M8211 OAI22X1_58/a_9_54# out_mines[9] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8212 OAI22X1_58/a_2_6# OAI22X1_64/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8213 vdd out_mines[8] OAI22X1_58/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8214 gnd out_temp_data_in[2] OAI22X1_36/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M8215 OAI22X1_36/a_2_6# OAI22X1_36/C INVX2_48/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M8216 INVX2_48/A OAI21X1_1/B OAI22X1_36/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8217 INVX2_48/A AND2X2_16/Y OAI22X1_36/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M8218 OAI22X1_36/a_28_54# OAI21X1_1/B INVX2_48/A vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M8219 OAI22X1_36/a_9_54# out_temp_data_in[2] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8220 OAI22X1_36/a_2_6# AND2X2_16/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8221 vdd OAI22X1_36/C OAI22X1_36/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8222 gnd out_mines[11] OAI22X1_69/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M8223 OAI22X1_69/a_2_6# out_mines[10] OAI22X1_69/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M8224 OAI22X1_69/Y OAI22X1_75/D OAI22X1_69/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8225 OAI22X1_69/Y OAI22X1_75/B OAI22X1_69/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M8226 OAI22X1_69/a_28_54# OAI22X1_75/D OAI22X1_69/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M8227 OAI22X1_69/a_9_54# out_mines[11] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8228 OAI22X1_69/a_2_6# OAI22X1_75/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8229 vdd out_mines[10] OAI22X1_69/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8230 gnd out_mines[4] OAI21X1_80/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M8231 vdd OAI21X1_80/C AOI21X1_6/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M8232 AOI21X1_6/C OAI21X1_80/C OAI21X1_80/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8233 AOI21X1_6/C OAI21X1_80/B OAI21X1_80/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8234 OAI21X1_80/a_9_54# out_mines[4] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8235 OAI21X1_80/a_2_6# OAI21X1_80/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8236 gnd INVX2_72/Y OAI21X1_91/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M8237 vdd OAI21X1_91/C OAI21X1_91/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M8238 OAI21X1_91/Y OAI21X1_91/C OAI21X1_91/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8239 OAI21X1_91/Y BUFX2_22/Y OAI21X1_91/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8240 OAI21X1_91/a_9_54# INVX2_72/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8241 OAI21X1_91/a_2_6# BUFX2_22/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8242 FAX1_18/a_46_54# FAX1_18/A vdd vdd pfet w=40 l=2
+  ad=0.452n pd=0.176m as=0 ps=0
M8243 gnd FAX1_18/A FAX1_18/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M8244 gnd FAX1_18/A FAX1_18/a_84_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M8245 FAX1_18/a_33_6# FAX1_18/B FAX1_18/a_25_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.12n ps=52u
M8246 FAX1_18/a_79_6# FAX1_18/C FAX1_18/a_70_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.14n ps=54u
M8247 FAX1_18/a_46_6# FAX1_18/A gnd Gnd nfet w=20 l=2
+  ad=0.24n pd=0.104m as=0 ps=0
M8248 FAX1_9/B FAX1_18/a_70_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8249 FAX1_18/a_46_6# FAX1_18/C gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8250 FAX1_18/a_79_46# FAX1_18/C FAX1_18/a_70_6# vdd pfet w=48 l=2
+  ad=0.144n pd=0.102m as=0.317n ps=0.11m
M8251 FAX1_8/A FAX1_18/a_25_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8252 FAX1_18/a_2_54# FAX1_18/B vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M8253 FAX1_18/a_25_6# FAX1_18/C FAX1_18/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8254 gnd FAX1_18/A FAX1_18/a_33_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8255 FAX1_18/a_70_6# FAX1_18/a_25_6# FAX1_18/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M8256 FAX1_18/a_84_6# FAX1_18/B FAX1_18/a_79_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8257 vdd FAX1_18/B FAX1_18/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M8258 vdd FAX1_18/A FAX1_18/a_84_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0.144n ps=0.102m
M8259 vdd FAX1_18/A FAX1_18/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8260 FAX1_9/B FAX1_18/a_70_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M8261 FAX1_18/a_25_6# FAX1_18/C FAX1_18/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M8262 gnd FAX1_18/B FAX1_18/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8263 vdd FAX1_18/A FAX1_18/a_33_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8264 FAX1_18/a_84_46# FAX1_18/B FAX1_18/a_79_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0 ps=0
M8265 FAX1_18/a_70_6# FAX1_18/a_25_6# FAX1_18/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8266 FAX1_18/a_46_54# FAX1_18/C vdd vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M8267 FAX1_8/A FAX1_18/a_25_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M8268 FAX1_18/a_2_6# FAX1_18/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8269 FAX1_18/a_33_54# FAX1_18/B FAX1_18/a_25_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8270 NAND3X1_50/Y out_decode vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M8271 NAND3X1_50/a_9_6# out_decode gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M8272 NAND3X1_50/Y NOR2X1_115/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8273 NAND3X1_50/Y NOR2X1_115/Y NAND3X1_50/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M8274 vdd AND2X2_17/Y NAND3X1_50/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8275 NAND3X1_50/a_14_6# AND2X2_17/Y NAND3X1_50/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M8276 NOR2X1_61/Y OAI21X1_4/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8277 NOR2X1_61/Y NOR2X1_64/A NOR2X1_61/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8278 NOR2X1_61/a_9_54# OAI21X1_4/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8279 gnd NOR2X1_64/A NOR2X1_61/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8280 NOR2X1_50/Y OR2X1_6/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8281 NOR2X1_50/Y NOR2X1_52/B NOR2X1_50/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8282 NOR2X1_50/a_9_54# OR2X1_6/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8283 gnd NOR2X1_52/B NOR2X1_50/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8284 NOR2X1_72/Y NOR2X1_72/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8285 NOR2X1_72/Y OR2X1_14/Y NOR2X1_72/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8286 NOR2X1_72/a_9_54# NOR2X1_72/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8287 gnd OR2X1_14/Y NOR2X1_72/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8288 NOR2X1_94/Y NOR2X1_94/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8289 NOR2X1_94/Y NOR2X1_94/B NOR2X1_94/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8290 NOR2X1_94/a_9_54# NOR2X1_94/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8291 gnd NOR2X1_94/B NOR2X1_94/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8292 NOR2X1_83/Y NOR2X1_83/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8293 NOR2X1_83/Y NOR2X1_83/B NOR2X1_83/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8294 NOR2X1_83/a_9_54# NOR2X1_83/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8295 gnd NOR2X1_83/B NOR2X1_83/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8296 OR2X1_11/A BUFX2_7/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8297 OR2X1_11/A BUFX2_7/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M8298 INVX2_32/A OAI21X1_1/A vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M8299 NAND2X1_107/a_9_6# OAI21X1_1/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M8300 vdd INVX2_30/Y INVX2_32/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8301 INVX2_32/A INVX2_30/Y NAND2X1_107/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8302 FAX1_8/a_46_54# FAX1_8/A vdd vdd pfet w=40 l=2
+  ad=0.452n pd=0.176m as=0 ps=0
M8303 gnd FAX1_8/A FAX1_8/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M8304 gnd FAX1_8/A FAX1_8/a_84_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M8305 FAX1_8/a_33_6# FAX1_8/B FAX1_8/a_25_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.12n ps=52u
M8306 FAX1_8/a_79_6# FAX1_8/C FAX1_8/a_70_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.14n ps=54u
M8307 FAX1_8/a_46_6# FAX1_8/A gnd Gnd nfet w=20 l=2
+  ad=0.24n pd=0.104m as=0 ps=0
M8308 FAX1_0/A FAX1_8/a_70_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8309 FAX1_8/a_46_6# FAX1_8/C gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8310 FAX1_8/a_79_46# FAX1_8/C FAX1_8/a_70_6# vdd pfet w=48 l=2
+  ad=0.144n pd=0.102m as=0.317n ps=0.11m
M8311 FAX1_7/C FAX1_8/a_25_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8312 FAX1_8/a_2_54# FAX1_8/B vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M8313 FAX1_8/a_25_6# FAX1_8/C FAX1_8/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8314 gnd FAX1_8/A FAX1_8/a_33_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8315 FAX1_8/a_70_6# FAX1_8/a_25_6# FAX1_8/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M8316 FAX1_8/a_84_6# FAX1_8/B FAX1_8/a_79_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8317 vdd FAX1_8/B FAX1_8/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M8318 vdd FAX1_8/A FAX1_8/a_84_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0.144n ps=0.102m
M8319 vdd FAX1_8/A FAX1_8/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8320 FAX1_0/A FAX1_8/a_70_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M8321 FAX1_8/a_25_6# FAX1_8/C FAX1_8/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M8322 gnd FAX1_8/B FAX1_8/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8323 vdd FAX1_8/A FAX1_8/a_33_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8324 FAX1_8/a_84_46# FAX1_8/B FAX1_8/a_79_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0 ps=0
M8325 FAX1_8/a_70_6# FAX1_8/a_25_6# FAX1_8/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8326 FAX1_8/a_46_54# FAX1_8/C vdd vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M8327 FAX1_7/C FAX1_8/a_25_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M8328 FAX1_8/a_2_6# FAX1_8/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8329 FAX1_8/a_33_54# FAX1_8/B FAX1_8/a_25_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8330 OAI21X1_157/B out_alu vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M8331 NAND2X1_129/a_9_6# out_alu gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M8332 vdd AND2X2_17/Y OAI21X1_157/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8333 OAI21X1_157/B AND2X2_17/Y NAND2X1_129/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8334 OAI22X1_64/B out_temp_data_in[0] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M8335 NAND2X1_118/a_9_6# out_temp_data_in[0] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M8336 vdd OR2X1_6/A OAI22X1_64/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8337 OAI22X1_64/B OR2X1_6/A NAND2X1_118/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8338 HAX1_38/B NOR2X1_5/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M8339 NAND2X1_5/a_9_6# NOR2X1_5/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M8340 vdd MUX2X1_3/Y HAX1_38/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8341 HAX1_38/B MUX2X1_3/Y NAND2X1_5/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8342 gnd XOR2X1_27/Y XNOR2X1_29/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M8343 XOR2X1_24/A XOR2X1_27/Y XNOR2X1_29/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M8344 XNOR2X1_29/a_12_41# INVX2_48/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8345 XNOR2X1_29/a_18_54# XNOR2X1_29/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M8346 XNOR2X1_29/a_35_6# XNOR2X1_29/a_2_6# XOR2X1_24/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M8347 XNOR2X1_29/a_18_6# XNOR2X1_29/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8348 vdd XOR2X1_27/Y XNOR2X1_29/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M8349 vdd INVX2_48/Y XNOR2X1_29/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8350 XOR2X1_24/A XNOR2X1_29/a_2_6# XNOR2X1_29/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M8351 XNOR2X1_29/a_35_54# XOR2X1_27/Y XOR2X1_24/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8352 XNOR2X1_29/a_12_41# INVX2_48/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M8353 gnd INVX2_48/Y XNOR2X1_29/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8354 gnd out_temp_data_in[0] XNOR2X1_18/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M8355 INVX2_37/A out_temp_data_in[0] XNOR2X1_18/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M8356 XNOR2X1_18/a_12_41# out_temp_data_in[1] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8357 XNOR2X1_18/a_18_54# XNOR2X1_18/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M8358 XNOR2X1_18/a_35_6# XNOR2X1_18/a_2_6# INVX2_37/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M8359 XNOR2X1_18/a_18_6# XNOR2X1_18/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8360 vdd out_temp_data_in[0] XNOR2X1_18/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M8361 vdd out_temp_data_in[1] XNOR2X1_18/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8362 INVX2_37/A XNOR2X1_18/a_2_6# XNOR2X1_18/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M8363 XNOR2X1_18/a_35_54# out_temp_data_in[0] INVX2_37/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8364 XNOR2X1_18/a_12_41# out_temp_data_in[1] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M8365 gnd out_temp_data_in[1] XNOR2X1_18/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8366 vdd BUFX2_2/Y BUFX2_17/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M8367 gnd BUFX2_2/Y BUFX2_17/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M8368 BUFX2_17/Y BUFX2_17/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M8369 BUFX2_17/Y BUFX2_17/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8370 NOR2X1_8/Y NOR2X1_9/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8371 NOR2X1_8/Y INVX2_1/Y NOR2X1_8/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8372 NOR2X1_8/a_9_54# NOR2X1_9/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8373 gnd INVX2_1/Y NOR2X1_8/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8374 AOI21X1_18/a_2_54# AOI21X1_18/B vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M8375 AOI21X1_18/a_12_6# AOI21X1_18/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M8376 gnd INVX2_36/Y AOI21X1_18/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0.11n ps=52u
M8377 vdd AOI21X1_18/A AOI21X1_18/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8378 AOI21X1_18/Y INVX2_36/Y AOI21X1_18/a_2_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M8379 AOI21X1_18/Y AOI21X1_18/B AOI21X1_18/a_12_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8380 OR2X1_5/a_2_54# OR2X1_5/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8381 OR2X1_5/Y OR2X1_5/a_2_54# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8382 OR2X1_5/Y OR2X1_5/a_2_54# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M8383 vdd OR2X1_5/B OR2X1_5/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8384 OR2X1_5/a_9_54# OR2X1_5/A OR2X1_5/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M8385 gnd OR2X1_5/B OR2X1_5/a_2_54# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8386 gnd BUFX2_25/Y OAI22X1_15/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M8387 OAI22X1_15/a_2_6# OAI22X1_5/C OAI22X1_15/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M8388 OAI22X1_15/Y INVX2_68/Y OAI22X1_15/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8389 OAI22X1_15/Y INVX2_100/Y OAI22X1_15/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M8390 OAI22X1_15/a_28_54# INVX2_68/Y OAI22X1_15/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M8391 OAI22X1_15/a_9_54# BUFX2_25/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8392 OAI22X1_15/a_2_6# INVX2_100/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8393 vdd OAI22X1_5/C OAI22X1_15/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8394 gnd out_mines[13] OAI22X1_48/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M8395 OAI22X1_48/a_2_6# out_mines[12] OAI22X1_48/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M8396 OAI22X1_48/Y OAI22X1_52/D OAI22X1_48/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8397 OAI22X1_48/Y OAI22X1_52/B OAI22X1_48/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M8398 OAI22X1_48/a_28_54# OAI22X1_52/D OAI22X1_48/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M8399 OAI22X1_48/a_9_54# out_mines[13] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8400 OAI22X1_48/a_2_6# OAI22X1_52/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8401 vdd out_mines[12] OAI22X1_48/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8402 gnd BUFX2_24/Y OAI22X1_26/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M8403 OAI22X1_26/a_2_6# OAI22X1_5/C OAI22X1_26/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M8404 OAI22X1_26/Y INVX2_82/Y OAI22X1_26/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8405 OAI22X1_26/Y INVX2_111/Y OAI22X1_26/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M8406 OAI22X1_26/a_28_54# INVX2_82/Y OAI22X1_26/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M8407 OAI22X1_26/a_9_54# BUFX2_24/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8408 OAI22X1_26/a_2_6# INVX2_111/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8409 vdd OAI22X1_5/C OAI22X1_26/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8410 gnd INVX2_43/Y OAI22X1_37/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M8411 OAI22X1_37/a_2_6# out_temp_data_in[1] INVX2_45/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M8412 INVX2_45/A OAI22X1_37/D OAI22X1_37/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8413 INVX2_45/A OR2X1_6/A OAI22X1_37/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M8414 OAI22X1_37/a_28_54# OAI22X1_37/D INVX2_45/A vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M8415 OAI22X1_37/a_9_54# INVX2_43/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8416 OAI22X1_37/a_2_6# OR2X1_6/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8417 vdd out_temp_data_in[1] OAI22X1_37/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8418 gnd out_mines[15] OAI22X1_59/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M8419 OAI22X1_59/a_2_6# out_mines[14] OAI22X1_59/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M8420 OAI22X1_59/Y OAI22X1_63/D OAI22X1_59/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8421 OAI22X1_59/Y OAI22X1_63/B OAI22X1_59/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M8422 OAI22X1_59/a_28_54# OAI22X1_63/D OAI22X1_59/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M8423 OAI22X1_59/a_9_54# out_mines[15] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8424 OAI22X1_59/a_2_6# OAI22X1_63/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8425 vdd out_mines[14] OAI22X1_59/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8426 gnd INVX2_23/Y OAI21X1_81/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M8427 vdd OAI21X1_81/C AOI21X1_7/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M8428 AOI21X1_7/C OAI21X1_81/C OAI21X1_81/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8429 AOI21X1_7/C INVX2_89/Y OAI21X1_81/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8430 OAI21X1_81/a_9_54# INVX2_23/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8431 OAI21X1_81/a_2_6# INVX2_89/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8432 gnd INVX2_6/Y OAI21X1_70/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M8433 vdd OAI21X1_70/C INVX2_80/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M8434 INVX2_80/A OAI21X1_70/C OAI21X1_70/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8435 INVX2_80/A INVX2_78/Y OAI21X1_70/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8436 OAI21X1_70/a_9_54# INVX2_6/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8437 OAI21X1_70/a_2_6# INVX2_78/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8438 gnd INVX2_71/Y OAI21X1_92/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M8439 vdd OAI21X1_92/C OAI21X1_92/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M8440 OAI21X1_92/Y OAI21X1_92/C OAI21X1_92/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8441 OAI21X1_92/Y BUFX2_22/Y OAI21X1_92/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8442 OAI21X1_92/a_9_54# INVX2_71/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8443 OAI21X1_92/a_2_6# BUFX2_22/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8444 OAI21X1_77/C INVX2_92/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M8445 NAND3X1_40/a_9_6# INVX2_92/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M8446 OAI21X1_77/C INVX2_19/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8447 OAI21X1_77/C INVX2_19/Y NAND3X1_40/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M8448 vdd INVX2_59/Y OAI21X1_77/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8449 NAND3X1_40/a_14_6# INVX2_59/Y NAND3X1_40/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M8450 OR2X1_15/A INVX2_120/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M8451 NAND3X1_51/a_9_6# INVX2_120/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M8452 OR2X1_15/A INVX2_119/A vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8453 OR2X1_15/A INVX2_119/A NAND3X1_51/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M8454 vdd INVX2_117/Y OR2X1_15/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8455 NAND3X1_51/a_14_6# INVX2_117/Y NAND3X1_51/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M8456 NOR2X1_62/Y OR2X1_12/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8457 NOR2X1_62/Y NOR2X1_64/B NOR2X1_62/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8458 NOR2X1_62/a_9_54# OR2X1_12/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8459 gnd NOR2X1_64/B NOR2X1_62/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8460 NOR2X1_51/Y NOR2X1_55/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8461 NOR2X1_51/Y NOR2X1_52/B NOR2X1_51/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8462 NOR2X1_51/a_9_54# NOR2X1_55/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8463 gnd NOR2X1_52/B NOR2X1_51/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8464 NOR2X1_40/Y INVX2_54/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8465 NOR2X1_40/Y NOR2X1_40/B NOR2X1_40/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8466 NOR2X1_40/a_9_54# INVX2_54/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8467 gnd NOR2X1_40/B NOR2X1_40/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8468 NOR2X1_73/Y NOR2X1_73/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8469 NOR2X1_73/Y NOR2X1_75/B NOR2X1_73/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8470 NOR2X1_73/a_9_54# NOR2X1_73/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8471 gnd NOR2X1_75/B NOR2X1_73/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8472 NOR2X1_95/Y out_temp_decoded[13] gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8473 NOR2X1_95/Y out_temp_cleared[13] NOR2X1_95/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8474 NOR2X1_95/a_9_54# out_temp_decoded[13] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8475 gnd out_temp_cleared[13] NOR2X1_95/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8476 NOR2X1_84/Y NOR2X1_84/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8477 NOR2X1_84/Y INVX2_62/A NOR2X1_84/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8478 NOR2X1_84/a_9_54# NOR2X1_84/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8479 gnd INVX2_62/A NOR2X1_84/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8480 INVX2_240/Y INVX2_240/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8481 INVX2_240/Y INVX2_240/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M8482 INVX2_251/Y out_temp_data_in[0] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8483 INVX2_251/Y out_temp_data_in[0] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M8484 NOR2X1_110/B out_temp_data_in[4] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M8485 NAND2X1_108/a_9_6# out_temp_data_in[4] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M8486 vdd OAI21X1_1/A NOR2X1_110/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8487 NOR2X1_110/B OAI21X1_1/A NAND2X1_108/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8488 FAX1_9/a_46_54# FAX1_9/A vdd vdd pfet w=40 l=2
+  ad=0.452n pd=0.176m as=0 ps=0
M8489 gnd FAX1_9/A FAX1_9/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M8490 gnd FAX1_9/A FAX1_9/a_84_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M8491 FAX1_9/a_33_6# FAX1_9/B FAX1_9/a_25_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.12n ps=52u
M8492 FAX1_9/a_79_6# FAX1_9/C FAX1_9/a_70_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0.14n ps=54u
M8493 FAX1_9/a_46_6# FAX1_9/A gnd Gnd nfet w=20 l=2
+  ad=0.24n pd=0.104m as=0 ps=0
M8494 FAX1_1/A FAX1_9/a_70_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8495 FAX1_9/a_46_6# FAX1_9/C gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8496 FAX1_9/a_79_46# FAX1_9/C FAX1_9/a_70_6# vdd pfet w=48 l=2
+  ad=0.144n pd=0.102m as=0.317n ps=0.11m
M8497 FAX1_8/C FAX1_9/a_25_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8498 FAX1_9/a_2_54# FAX1_9/B vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M8499 FAX1_9/a_25_6# FAX1_9/C FAX1_9/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8500 gnd FAX1_9/A FAX1_9/a_33_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8501 FAX1_9/a_70_6# FAX1_9/a_25_6# FAX1_9/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M8502 FAX1_9/a_84_6# FAX1_9/B FAX1_9/a_79_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8503 vdd FAX1_9/B FAX1_9/a_46_54# vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M8504 vdd FAX1_9/A FAX1_9/a_84_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0.144n ps=0.102m
M8505 vdd FAX1_9/A FAX1_9/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8506 FAX1_1/A FAX1_9/a_70_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M8507 FAX1_9/a_25_6# FAX1_9/C FAX1_9/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M8508 gnd FAX1_9/B FAX1_9/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8509 vdd FAX1_9/A FAX1_9/a_33_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8510 FAX1_9/a_84_46# FAX1_9/B FAX1_9/a_79_46# vdd pfet w=48 l=2
+  ad=0 pd=0 as=0 ps=0
M8511 FAX1_9/a_70_6# FAX1_9/a_25_6# FAX1_9/a_46_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8512 FAX1_9/a_46_54# FAX1_9/C vdd vdd pfet w=36 l=2
+  ad=0 pd=0 as=0 ps=0
M8513 FAX1_8/C FAX1_9/a_25_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M8514 FAX1_9/a_2_6# FAX1_9/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8515 FAX1_9/a_33_54# FAX1_9/B FAX1_9/a_25_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8516 AOI22X1_74/A OAI21X1_146/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M8517 NAND2X1_119/a_9_6# OAI21X1_146/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M8518 vdd OAI21X1_145/Y AOI22X1_74/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8519 AOI22X1_74/A OAI21X1_145/Y NAND2X1_119/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8520 XOR2X1_0/A NOR2X1_6/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M8521 NAND2X1_6/a_9_6# NOR2X1_6/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M8522 vdd NAND2X1_6/B XOR2X1_0/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8523 XOR2X1_0/A NAND2X1_6/B NAND2X1_6/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8524 gnd OR2X1_10/B XNOR2X1_19/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M8525 INVX2_36/A OR2X1_10/B XNOR2X1_19/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M8526 XNOR2X1_19/a_12_41# out_temp_data_in[3] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8527 XNOR2X1_19/a_18_54# XNOR2X1_19/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M8528 XNOR2X1_19/a_35_6# XNOR2X1_19/a_2_6# INVX2_36/A Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M8529 XNOR2X1_19/a_18_6# XNOR2X1_19/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8530 vdd OR2X1_10/B XNOR2X1_19/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M8531 vdd out_temp_data_in[3] XNOR2X1_19/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8532 INVX2_36/A XNOR2X1_19/a_2_6# XNOR2X1_19/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M8533 XNOR2X1_19/a_35_54# OR2X1_10/B INVX2_36/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8534 XNOR2X1_19/a_12_41# out_temp_data_in[3] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M8535 gnd out_temp_data_in[3] XNOR2X1_19/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8536 vdd BUFX2_19/A BUFX2_18/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M8537 gnd BUFX2_19/A BUFX2_18/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M8538 BUFX2_18/Y BUFX2_18/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M8539 BUFX2_18/Y BUFX2_18/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8540 HAX1_30/B NOR2X1_9/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8541 HAX1_30/B INVX2_2/Y NOR2X1_9/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8542 NOR2X1_9/a_9_54# NOR2X1_9/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8543 gnd INVX2_2/Y HAX1_30/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8544 AOI21X1_19/a_2_54# NOR2X1_116/Y vdd vdd pfet w=40 l=2
+  ad=0.44n pd=0.182m as=0 ps=0
M8545 AOI21X1_19/a_12_6# INVX2_117/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M8546 gnd INVX2_128/Y AND2X2_17/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0.11n ps=52u
M8547 vdd INVX2_117/Y AOI21X1_19/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8548 AND2X2_17/A INVX2_128/Y AOI21X1_19/a_2_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M8549 AND2X2_17/A NOR2X1_116/Y AOI21X1_19/a_12_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8550 OR2X1_6/a_2_54# OR2X1_6/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8551 OR2X1_6/Y OR2X1_6/a_2_54# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8552 OR2X1_6/Y OR2X1_6/a_2_54# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M8553 vdd out_temp_data_in[0] OR2X1_6/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8554 OR2X1_6/a_9_54# OR2X1_6/A OR2X1_6/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M8555 gnd out_temp_data_in[0] OR2X1_6/a_2_54# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8556 gnd out_mines[19] OAI22X1_49/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M8557 OAI22X1_49/a_2_6# out_mines[18] OAI22X1_49/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M8558 OAI22X1_49/Y OAI22X1_51/D OAI22X1_49/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8559 OAI22X1_49/Y OAI22X1_51/B OAI22X1_49/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M8560 OAI22X1_49/a_28_54# OAI22X1_51/D OAI22X1_49/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M8561 OAI22X1_49/a_9_54# out_mines[19] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8562 OAI22X1_49/a_2_6# OAI22X1_51/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8563 vdd out_mines[18] OAI22X1_49/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8564 gnd BUFX2_25/Y OAI22X1_16/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M8565 OAI22X1_16/a_2_6# OR2X1_11/A OAI22X1_16/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M8566 OAI22X1_16/Y INVX2_69/Y OAI22X1_16/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8567 OAI22X1_16/Y INVX2_101/Y OAI22X1_16/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M8568 OAI22X1_16/a_28_54# INVX2_69/Y OAI22X1_16/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M8569 OAI22X1_16/a_9_54# BUFX2_25/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8570 OAI22X1_16/a_2_6# INVX2_101/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8571 vdd OR2X1_11/A OAI22X1_16/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8572 gnd INVX2_41/A OAI22X1_38/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M8573 OAI22X1_38/a_2_6# OAI22X1_38/C AOI21X1_8/C Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M8574 AOI21X1_8/C INVX2_22/Y OAI22X1_38/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8575 AOI21X1_8/C INVX2_16/Y OAI22X1_38/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M8576 OAI22X1_38/a_28_54# INVX2_22/Y AOI21X1_8/C vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M8577 OAI22X1_38/a_9_54# INVX2_41/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8578 OAI22X1_38/a_2_6# INVX2_16/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8579 vdd OAI22X1_38/C OAI22X1_38/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8580 gnd BUFX2_24/Y OAI22X1_27/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M8581 OAI22X1_27/a_2_6# OAI22X1_5/C OAI22X1_27/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M8582 OAI22X1_27/Y INVX2_83/Y OAI22X1_27/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8583 OAI22X1_27/Y OAI22X1_3/B OAI22X1_27/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M8584 OAI22X1_27/a_28_54# INVX2_83/Y OAI22X1_27/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M8585 OAI22X1_27/a_9_54# BUFX2_24/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8586 OAI22X1_27/a_2_6# OAI22X1_3/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8587 vdd OAI22X1_5/C OAI22X1_27/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8588 gnd INVX2_7/Y OAI21X1_71/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M8589 vdd OAI21X1_71/C NOR2X1_85/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M8590 NOR2X1_85/B OAI21X1_71/C OAI21X1_71/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8591 NOR2X1_85/B INVX2_107/Y OAI21X1_71/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8592 OAI21X1_71/a_9_54# INVX2_7/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8593 OAI21X1_71/a_2_6# INVX2_107/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8594 gnd OAI21X1_60/A OAI21X1_60/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M8595 vdd OAI21X1_60/C OAI21X1_60/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M8596 OAI21X1_60/Y OAI21X1_60/C OAI21X1_60/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8597 OAI21X1_60/Y OAI21X1_62/B OAI21X1_60/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8598 OAI21X1_60/a_9_54# OAI21X1_60/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8599 OAI21X1_60/a_2_6# OAI21X1_62/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8600 gnd INVX2_70/Y OAI21X1_93/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M8601 vdd OAI21X1_93/C OAI21X1_93/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M8602 OAI21X1_93/Y OAI21X1_93/C OAI21X1_93/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8603 OAI21X1_93/Y BUFX2_22/Y OAI21X1_93/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8604 OAI21X1_93/a_9_54# INVX2_70/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8605 OAI21X1_93/a_2_6# BUFX2_22/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8606 gnd INVX2_85/Y OAI21X1_82/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M8607 vdd OAI21X1_82/C OAI21X1_82/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M8608 OAI21X1_82/Y OAI21X1_82/C OAI21X1_82/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8609 OAI21X1_82/Y BUFX2_23/A OAI21X1_82/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8610 OAI21X1_82/a_9_54# INVX2_85/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8611 OAI21X1_82/a_2_6# BUFX2_23/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8612 NOR2X1_91/A NAND3X1_41/A vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M8613 NAND3X1_41/a_9_6# NAND3X1_41/A gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M8614 NOR2X1_91/A NOR2X1_94/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8615 NOR2X1_91/A NOR2X1_94/Y NAND3X1_41/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M8616 vdd NAND3X1_41/B NOR2X1_91/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8617 NAND3X1_41/a_14_6# NAND3X1_41/B NAND3X1_41/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M8618 NOR2X1_83/A INVX2_80/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M8619 NAND3X1_30/a_9_6# INVX2_80/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M8620 NOR2X1_83/A NOR2X1_84/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8621 NOR2X1_83/A NOR2X1_84/Y NAND3X1_30/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M8622 vdd AOI21X1_4/Y NOR2X1_83/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8623 NAND3X1_30/a_14_6# AOI21X1_4/Y NAND3X1_30/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M8624 NAND3X1_52/Y INVX2_127/A vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M8625 NAND3X1_52/a_9_6# INVX2_127/A gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M8626 NAND3X1_52/Y NOR2X1_116/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8627 NAND3X1_52/Y NOR2X1_116/Y NAND3X1_52/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M8628 vdd INVX2_117/Y NAND3X1_52/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8629 NAND3X1_52/a_14_6# INVX2_117/Y NAND3X1_52/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M8630 FAX1_13/B INVX2_3/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8631 FAX1_13/B NOR2X1_32/B NOR2X1_30/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8632 NOR2X1_30/a_9_54# INVX2_3/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8633 gnd NOR2X1_32/B FAX1_13/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8634 NOR2X1_63/Y NOR2X1_66/B gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8635 NOR2X1_63/Y NOR2X1_63/B NOR2X1_63/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8636 NOR2X1_63/a_9_54# NOR2X1_66/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8637 gnd NOR2X1_63/B NOR2X1_63/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8638 NOR2X1_52/Y INVX2_54/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8639 NOR2X1_52/Y NOR2X1_52/B NOR2X1_52/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8640 NOR2X1_52/a_9_54# INVX2_54/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8641 gnd NOR2X1_52/B NOR2X1_52/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8642 NOR2X1_41/Y NOR2X1_57/B gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8643 NOR2X1_41/Y NOR2X1_59/B NOR2X1_41/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8644 NOR2X1_41/a_9_54# NOR2X1_57/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8645 gnd NOR2X1_59/B NOR2X1_41/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8646 NOR2X1_96/Y out_temp_decoded[12] gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8647 NOR2X1_96/Y out_temp_cleared[12] NOR2X1_96/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8648 NOR2X1_96/a_9_54# out_temp_decoded[12] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8649 gnd out_temp_cleared[12] NOR2X1_96/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8650 NOR2X1_85/Y NOR2X1_85/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8651 NOR2X1_85/Y NOR2X1_85/B NOR2X1_85/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8652 NOR2X1_85/a_9_54# NOR2X1_85/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8653 gnd NOR2X1_85/B NOR2X1_85/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8654 NOR2X1_74/Y out_temp_decoded[5] gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8655 NOR2X1_74/Y out_temp_decoded[20] NOR2X1_74/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8656 NOR2X1_74/a_9_54# out_temp_decoded[5] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8657 gnd out_temp_decoded[20] NOR2X1_74/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8658 INVX2_230/Y INVX2_230/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8659 INVX2_230/Y INVX2_230/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M8660 INVX2_241/Y INVX2_241/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8661 INVX2_241/Y INVX2_241/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M8662 OR2X1_6/A out_temp_data_in[1] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8663 OR2X1_6/A out_temp_data_in[1] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M8664 AOI22X1_72/A OAI21X1_130/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M8665 NAND2X1_109/a_9_6# OAI21X1_130/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M8666 vdd OAI21X1_129/Y AOI22X1_72/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8667 AOI22X1_72/A OAI21X1_129/Y NAND2X1_109/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8668 NOR2X1_7/B XOR2X1_5/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M8669 NAND2X1_7/a_9_6# XOR2X1_5/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M8670 vdd XOR2X1_0/A NOR2X1_7/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8671 NOR2X1_7/B XOR2X1_0/A NAND2X1_7/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8672 NOR2X1_120/Y out_state_main[2] gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8673 NOR2X1_120/Y out_state_main[1] NOR2X1_120/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8674 NOR2X1_120/a_9_54# out_state_main[2] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8675 gnd out_state_main[1] NOR2X1_120/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8676 vdd BUFX2_19/A BUFX2_19/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M8677 gnd BUFX2_19/A BUFX2_19/a_2_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M8678 BUFX2_19/Y BUFX2_19/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M8679 BUFX2_19/Y BUFX2_19/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8680 OR2X1_7/a_2_54# out_temp_data_in[3] gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8681 OR2X1_7/Y OR2X1_7/a_2_54# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8682 OR2X1_7/Y OR2X1_7/a_2_54# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M8683 vdd out_temp_data_in[2] OR2X1_7/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8684 OR2X1_7/a_9_54# out_temp_data_in[3] OR2X1_7/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M8685 gnd out_temp_data_in[2] OR2X1_7/a_2_54# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8686 gnd BUFX2_24/Y OAI22X1_17/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M8687 OAI22X1_17/a_2_6# OAI22X1_5/C OAI22X1_17/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M8688 OAI22X1_17/Y INVX2_70/Y OAI22X1_17/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8689 OAI22X1_17/Y INVX2_102/Y OAI22X1_17/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M8690 OAI22X1_17/a_28_54# INVX2_70/Y OAI22X1_17/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M8691 OAI22X1_17/a_9_54# BUFX2_24/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8692 OAI22X1_17/a_2_6# INVX2_102/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8693 vdd OAI22X1_5/C OAI22X1_17/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8694 gnd INVX2_14/Y OAI22X1_39/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M8695 OAI22X1_39/a_2_6# INVX2_8/Y OAI22X1_39/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M8696 OAI22X1_39/Y INVX2_32/A OAI22X1_39/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8697 OAI22X1_39/Y INVX2_31/A OAI22X1_39/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M8698 OAI22X1_39/a_28_54# INVX2_32/A OAI22X1_39/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M8699 OAI22X1_39/a_9_54# INVX2_14/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8700 OAI22X1_39/a_2_6# INVX2_31/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8701 vdd INVX2_8/Y OAI22X1_39/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8702 gnd BUFX2_24/Y OAI22X1_28/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M8703 OAI22X1_28/a_2_6# OR2X1_11/A OAI22X1_28/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M8704 OAI22X1_28/Y INVX2_85/Y OAI22X1_28/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8705 OAI22X1_28/Y OAI22X1_3/D OAI22X1_28/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M8706 OAI22X1_28/a_28_54# INVX2_85/Y OAI22X1_28/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M8707 OAI22X1_28/a_9_54# BUFX2_24/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8708 OAI22X1_28/a_2_6# OAI22X1_3/D gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8709 vdd OR2X1_11/A OAI22X1_28/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8710 gnd NAND3X1_8/Y OAI21X1_50/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M8711 vdd BUFX2_18/Y INVX2_222/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M8712 INVX2_222/A BUFX2_18/Y OAI21X1_50/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8713 INVX2_222/A INVX2_179/Y OAI21X1_50/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8714 OAI21X1_50/a_9_54# NAND3X1_8/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8715 OAI21X1_50/a_2_6# INVX2_179/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8716 gnd out_mines[7] OAI21X1_72/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M8717 vdd OAI21X1_72/C NOR2X1_85/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M8718 NOR2X1_85/A OAI21X1_72/C OAI21X1_72/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8719 NOR2X1_85/A OAI21X1_72/B OAI21X1_72/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8720 OAI21X1_72/a_9_54# out_mines[7] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8721 OAI21X1_72/a_2_6# OAI21X1_72/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8722 gnd XNOR2X1_20/Y OAI21X1_61/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M8723 vdd AOI22X1_0/Y OAI21X1_61/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M8724 OAI21X1_61/Y AOI22X1_0/Y OAI21X1_61/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8725 OAI21X1_61/Y OR2X1_14/Y OAI21X1_61/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8726 OAI21X1_61/a_9_54# XNOR2X1_20/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8727 OAI21X1_61/a_2_6# OR2X1_14/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8728 gnd INVX2_69/Y OAI21X1_94/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M8729 vdd OAI21X1_94/C OAI21X1_94/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M8730 OAI21X1_94/Y OAI21X1_94/C OAI21X1_94/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8731 OAI21X1_94/Y BUFX2_22/Y OAI21X1_94/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8732 OAI21X1_94/a_9_54# INVX2_69/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8733 OAI21X1_94/a_2_6# BUFX2_22/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8734 gnd INVX2_83/Y OAI21X1_83/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M8735 vdd OAI21X1_83/C OAI21X1_83/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M8736 OAI21X1_83/Y OAI21X1_83/C OAI21X1_83/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8737 OAI21X1_83/Y BUFX2_22/Y OAI21X1_83/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8738 OAI21X1_83/a_9_54# INVX2_83/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8739 OAI21X1_83/a_2_6# BUFX2_22/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8740 OR2X1_10/a_2_54# out_temp_data_in[3] gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8741 OR2X1_10/Y OR2X1_10/a_2_54# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8742 OR2X1_10/Y OR2X1_10/a_2_54# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M8743 vdd OR2X1_10/B OR2X1_10/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8744 OR2X1_10/a_9_54# out_temp_data_in[3] OR2X1_10/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M8745 gnd OR2X1_10/B OR2X1_10/a_2_54# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8746 OAI21X1_71/C OAI22X1_1/B vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M8747 NAND3X1_31/a_9_6# OAI22X1_1/B gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M8748 OAI21X1_71/C INVX2_15/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8749 OAI21X1_71/C INVX2_15/Y NAND3X1_31/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M8750 vdd INVX2_74/Y OAI21X1_71/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8751 NAND3X1_31/a_14_6# INVX2_74/Y NAND3X1_31/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M8752 INVX2_84/A INVX2_82/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M8753 NAND3X1_20/a_9_6# INVX2_82/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M8754 INVX2_84/A INVX2_83/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8755 INVX2_84/A INVX2_83/Y NAND3X1_20/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M8756 vdd INVX2_81/Y INVX2_84/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8757 NAND3X1_20/a_14_6# INVX2_81/Y NAND3X1_20/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M8758 INVX2_128/A OR2X1_15/B vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M8759 NAND3X1_53/a_9_6# OR2X1_15/B gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M8760 INVX2_128/A NOR2X1_125/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8761 INVX2_128/A NOR2X1_125/Y NAND3X1_53/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M8762 vdd INVX2_119/Y INVX2_128/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8763 NAND3X1_53/a_14_6# INVX2_119/Y NAND3X1_53/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M8764 OAI21X1_78/C INVX2_96/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M8765 NAND3X1_42/a_9_6# INVX2_96/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M8766 OAI21X1_78/C INVX2_22/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8767 OAI21X1_78/C INVX2_22/Y NAND3X1_42/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M8768 vdd INVX2_64/Y OAI21X1_78/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8769 NAND3X1_42/a_14_6# INVX2_64/Y NAND3X1_42/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M8770 FAX1_17/B INVX2_3/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8771 FAX1_17/B NOR2X1_22/B NOR2X1_20/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8772 NOR2X1_20/a_9_54# INVX2_3/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8773 gnd NOR2X1_22/B FAX1_17/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8774 NOR2X1_64/Y NOR2X1_64/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8775 NOR2X1_64/Y NOR2X1_64/B NOR2X1_64/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8776 NOR2X1_64/a_9_54# NOR2X1_64/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8777 gnd NOR2X1_64/B NOR2X1_64/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8778 FAX1_11/B INVX2_4/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8779 FAX1_11/B NOR2X1_32/B NOR2X1_31/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8780 NOR2X1_31/a_9_54# INVX2_4/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8781 gnd NOR2X1_32/B FAX1_11/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8782 NOR2X1_53/Y NOR2X1_57/B gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8783 NOR2X1_53/Y NOR2X1_56/B NOR2X1_53/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8784 NOR2X1_53/a_9_54# NOR2X1_57/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8785 gnd NOR2X1_56/B NOR2X1_53/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8786 NOR2X1_42/Y OR2X1_6/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8787 NOR2X1_42/Y NOR2X1_59/B NOR2X1_42/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8788 NOR2X1_42/a_9_54# OR2X1_6/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8789 gnd NOR2X1_59/B NOR2X1_42/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8790 NOR2X1_86/Y NOR2X1_86/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8791 NOR2X1_86/Y OAI22X1_1/Y NOR2X1_86/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8792 NOR2X1_86/a_9_54# NOR2X1_86/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8793 gnd OAI22X1_1/Y NOR2X1_86/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8794 NOR2X1_97/Y NOR2X1_97/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8795 NOR2X1_97/Y NOR2X1_97/B NOR2X1_97/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8796 NOR2X1_97/a_9_54# NOR2X1_97/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8797 gnd NOR2X1_97/B NOR2X1_97/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8798 NOR2X1_75/Y out_temp_decoded[4] gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8799 NOR2X1_75/Y NOR2X1_75/B NOR2X1_75/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8800 NOR2X1_75/a_9_54# out_temp_decoded[4] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8801 gnd NOR2X1_75/B NOR2X1_75/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8802 INVX2_220/Y INVX2_220/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8803 INVX2_220/Y INVX2_220/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M8804 INVX2_231/Y INVX2_231/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8805 INVX2_231/Y INVX2_231/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M8806 OAI21X1_9/B BUFX2_6/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8807 OAI21X1_9/B BUFX2_6/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M8808 INVX2_242/Y INVX2_242/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8809 INVX2_242/Y INVX2_242/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M8810 OAI21X1_0/C OAI21X1_0/A vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M8811 NAND2X1_8/a_9_6# OAI21X1_0/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M8812 vdd OAI21X1_1/B OAI21X1_0/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8813 OAI21X1_0/C OAI21X1_1/B NAND2X1_8/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8814 NOR2X1_121/Y INVX2_125/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8815 NOR2X1_121/Y out_state_main[2] NOR2X1_121/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8816 NOR2X1_121/a_9_54# INVX2_125/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8817 gnd out_state_main[2] NOR2X1_121/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8818 NOR2X1_110/Y INVX2_47/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8819 NOR2X1_110/Y NOR2X1_110/B NOR2X1_110/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8820 NOR2X1_110/a_9_54# INVX2_47/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8821 gnd NOR2X1_110/B NOR2X1_110/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8822 OR2X1_8/a_2_54# out_temp_data_in[3] gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8823 OR2X1_8/Y OR2X1_8/a_2_54# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8824 OR2X1_8/Y OR2X1_8/a_2_54# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M8825 vdd OR2X1_8/B OR2X1_8/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8826 OR2X1_8/a_9_54# out_temp_data_in[3] OR2X1_8/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M8827 gnd OR2X1_8/B OR2X1_8/a_2_54# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8828 gnd BUFX2_24/Y OAI22X1_18/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M8829 OAI22X1_18/a_2_6# OR2X1_11/A OAI22X1_18/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M8830 OAI22X1_18/Y INVX2_71/Y OAI22X1_18/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8831 OAI22X1_18/Y INVX2_103/Y OAI22X1_18/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M8832 OAI22X1_18/a_28_54# INVX2_71/Y OAI22X1_18/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M8833 OAI22X1_18/a_9_54# BUFX2_24/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8834 OAI22X1_18/a_2_6# INVX2_103/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8835 vdd OR2X1_11/A OAI22X1_18/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8836 gnd XOR2X1_19/Y OAI22X1_29/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M8837 OAI22X1_29/a_2_6# XOR2X1_25/B XNOR2X1_25/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M8838 XNOR2X1_25/A INVX2_40/A OAI22X1_29/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8839 XNOR2X1_25/A XOR2X1_28/A OAI22X1_29/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M8840 OAI22X1_29/a_28_54# INVX2_40/A XNOR2X1_25/A vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M8841 OAI22X1_29/a_9_54# XOR2X1_19/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8842 OAI22X1_29/a_2_6# XOR2X1_28/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8843 vdd XOR2X1_25/B OAI22X1_29/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8844 gnd INVX2_226/Y OAI21X1_51/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M8845 vdd OAI21X1_51/C OAI21X1_51/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M8846 OAI21X1_51/Y OAI21X1_51/C OAI21X1_51/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8847 OAI21X1_51/Y NOR2X1_66/B OAI21X1_51/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8848 OAI21X1_51/a_9_54# INVX2_226/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8849 OAI21X1_51/a_2_6# NOR2X1_66/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8850 gnd OAI21X1_8/A OAI21X1_40/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M8851 vdd BUFX2_18/Y INVX2_232/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M8852 INVX2_232/A BUFX2_18/Y OAI21X1_40/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8853 INVX2_232/A OAI21X1_48/B OAI21X1_40/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8854 OAI21X1_40/a_9_54# OAI21X1_8/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8855 OAI21X1_40/a_2_6# OAI21X1_48/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8856 gnd OAI21X1_63/Y OAI21X1_62/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M8857 vdd OAI21X1_62/C OAI21X1_62/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M8858 OAI21X1_62/Y OAI21X1_62/C OAI21X1_62/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8859 OAI21X1_62/Y OAI21X1_62/B OAI21X1_62/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8860 OAI21X1_62/a_9_54# OAI21X1_63/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8861 OAI21X1_62/a_2_6# OAI21X1_62/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8862 gnd INVX2_13/Y OAI21X1_73/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M8863 vdd OAI21X1_73/C NOR2X1_86/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M8864 NOR2X1_86/A OAI21X1_73/C OAI21X1_73/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8865 NOR2X1_86/A INVX2_67/Y OAI21X1_73/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8866 OAI21X1_73/a_9_54# INVX2_13/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8867 OAI21X1_73/a_2_6# INVX2_67/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8868 gnd INVX2_68/Y OAI21X1_95/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M8869 vdd OAI21X1_95/C OAI21X1_95/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M8870 OAI21X1_95/Y OAI21X1_95/C OAI21X1_95/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8871 OAI21X1_95/Y BUFX2_23/Y OAI21X1_95/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8872 OAI21X1_95/a_9_54# INVX2_68/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8873 OAI21X1_95/a_2_6# BUFX2_23/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8874 gnd INVX2_82/Y OAI21X1_84/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M8875 vdd OAI21X1_84/C OAI21X1_84/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M8876 OAI21X1_84/Y OAI21X1_84/C OAI21X1_84/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8877 OAI21X1_84/Y BUFX2_22/Y OAI21X1_84/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8878 OAI21X1_84/a_9_54# INVX2_82/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8879 OAI21X1_84/a_2_6# BUFX2_22/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8880 OR2X1_11/a_2_54# OR2X1_11/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8881 OR2X1_11/Y OR2X1_11/a_2_54# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8882 OR2X1_11/Y OR2X1_11/a_2_54# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M8883 vdd OR2X1_11/B OR2X1_11/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8884 OR2X1_11/a_9_54# OR2X1_11/A OR2X1_11/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M8885 gnd OR2X1_11/B OR2X1_11/a_2_54# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8886 AND2X2_10/a_2_6# HAX1_35/YS vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M8887 AND2X2_10/a_9_6# HAX1_35/YS AND2X2_10/a_2_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=100p ps=50u
M8888 AND2X2_10/Y AND2X2_10/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8889 AND2X2_10/Y AND2X2_10/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M8890 vdd BUFX2_8/Y AND2X2_10/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8891 gnd BUFX2_8/Y AND2X2_10/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8892 OR2X1_13/B XNOR2X1_23/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M8893 NAND3X1_10/a_9_6# XNOR2X1_23/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M8894 OR2X1_13/B NOR2X1_68/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8895 OR2X1_13/B NOR2X1_68/Y NAND3X1_10/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M8896 vdd XNOR2X1_22/Y OR2X1_13/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8897 NAND3X1_10/a_14_6# XNOR2X1_22/Y NAND3X1_10/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M8898 NOR2X1_77/B INVX2_57/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M8899 NAND3X1_21/a_9_6# INVX2_57/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M8900 NOR2X1_77/B INVX2_59/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8901 NOR2X1_77/B INVX2_59/Y NAND3X1_21/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M8902 vdd INVX2_56/Y NOR2X1_77/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8903 NAND3X1_21/a_14_6# INVX2_56/Y NAND3X1_21/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M8904 OAI21X1_72/C INVX2_107/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M8905 NAND3X1_32/a_9_6# INVX2_107/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M8906 OAI21X1_72/C INVX2_7/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8907 OAI21X1_72/C INVX2_7/Y NAND3X1_32/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M8908 vdd INVX2_77/Y OAI21X1_72/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8909 NAND3X1_32/a_14_6# INVX2_77/Y NAND3X1_32/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M8910 OAI21X1_79/C INVX2_98/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M8911 NAND3X1_43/a_9_6# INVX2_98/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M8912 OAI21X1_79/C INVX2_11/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8913 OAI21X1_79/C INVX2_11/Y NAND3X1_43/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M8914 vdd INVX2_66/Y OAI21X1_79/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8915 NAND3X1_43/a_14_6# INVX2_66/Y NAND3X1_43/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M8916 AND2X2_19/B out_display_done vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M8917 NAND3X1_54/a_9_6# out_display_done gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M8918 AND2X2_19/B INVX2_122/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8919 AND2X2_19/B INVX2_122/Y NAND3X1_54/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M8920 vdd in_data_in AND2X2_19/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8921 NAND3X1_54/a_14_6# in_data_in NAND3X1_54/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M8922 HAX1_34/A NOR2X1_9/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8923 HAX1_34/A INVX2_3/Y NOR2X1_10/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8924 NOR2X1_10/a_9_54# NOR2X1_9/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8925 gnd INVX2_3/Y HAX1_34/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8926 FAX1_15/B INVX2_4/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8927 FAX1_15/B NOR2X1_22/B NOR2X1_21/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8928 NOR2X1_21/a_9_54# INVX2_4/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8929 gnd NOR2X1_22/B FAX1_15/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8930 FAX1_4/A INVX2_17/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8931 FAX1_4/A NOR2X1_32/B NOR2X1_32/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8932 NOR2X1_32/a_9_54# INVX2_17/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8933 gnd NOR2X1_32/B FAX1_4/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8934 NOR2X1_54/Y OR2X1_6/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8935 NOR2X1_54/Y NOR2X1_56/B NOR2X1_54/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8936 NOR2X1_54/a_9_54# OR2X1_6/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8937 gnd NOR2X1_56/B NOR2X1_54/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8938 NOR2X1_43/Y NOR2X1_43/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8939 NOR2X1_43/Y NOR2X1_43/B NOR2X1_43/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8940 NOR2X1_43/a_9_54# NOR2X1_43/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8941 gnd NOR2X1_43/B NOR2X1_43/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8942 NOR2X1_65/Y NOR2X1_65/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8943 NOR2X1_65/Y NOR2X1_66/B NOR2X1_65/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8944 NOR2X1_65/a_9_54# NOR2X1_65/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8945 gnd NOR2X1_66/B NOR2X1_65/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8946 NOR2X1_87/Y NOR2X1_87/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8947 NOR2X1_87/Y NOR2X1_87/B NOR2X1_87/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8948 NOR2X1_87/a_9_54# NOR2X1_87/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8949 gnd NOR2X1_87/B NOR2X1_87/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8950 NOR2X1_76/Y out_temp_decoded[9] gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8951 NOR2X1_76/Y out_temp_decoded[24] NOR2X1_76/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8952 NOR2X1_76/a_9_54# out_temp_decoded[9] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8953 gnd out_temp_decoded[24] NOR2X1_76/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8954 NOR2X1_98/Y out_temp_decoded[5] gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8955 NOR2X1_98/Y out_temp_cleared[5] NOR2X1_98/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8956 NOR2X1_98/a_9_54# out_temp_decoded[5] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8957 gnd out_temp_cleared[5] NOR2X1_98/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8958 INVX2_210/Y INVX2_210/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8959 INVX2_210/Y INVX2_210/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M8960 INVX2_221/Y INVX2_221/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8961 INVX2_221/Y INVX2_221/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M8962 INVX2_232/Y INVX2_232/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8963 INVX2_232/Y INVX2_232/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M8964 INVX2_243/Y INVX2_243/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8965 INVX2_243/Y INVX2_243/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M8966 OAI21X1_1/B out_temp_data_in[2] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8967 OAI21X1_1/B out_temp_data_in[2] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M8968 NOR2X1_43/B out_temp_data_in[4] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M8969 NAND2X1_9/a_9_6# out_temp_data_in[4] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M8970 vdd INVX2_54/A NOR2X1_43/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8971 NOR2X1_43/B INVX2_54/A NAND2X1_9/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8972 AOI21X1_7/A out_temp_decoded[19] gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8973 AOI21X1_7/A out_temp_cleared[19] NOR2X1_100/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8974 NOR2X1_100/a_9_54# out_temp_decoded[19] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8975 gnd out_temp_cleared[19] AOI21X1_7/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8976 NOR2X1_122/Y out_state_main[3] gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8977 NOR2X1_122/Y out_state_main[0] NOR2X1_122/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8978 NOR2X1_122/a_9_54# out_state_main[3] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8979 gnd out_state_main[0] NOR2X1_122/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8980 NOR2X1_111/Y INVX2_251/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8981 NOR2X1_111/Y out_temp_data_in[1] NOR2X1_111/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M8982 NOR2X1_111/a_9_54# INVX2_251/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8983 gnd out_temp_data_in[1] NOR2X1_111/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8984 OR2X1_9/a_2_54# out_temp_data_in[1] gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M8985 OR2X1_9/Y OR2X1_9/a_2_54# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M8986 OR2X1_9/Y OR2X1_9/a_2_54# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M8987 vdd out_temp_data_in[0] OR2X1_9/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M8988 OR2X1_9/a_9_54# out_temp_data_in[1] OR2X1_9/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M8989 gnd out_temp_data_in[0] OR2X1_9/a_2_54# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M8990 gnd BUFX2_24/Y OAI22X1_19/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M8991 OAI22X1_19/a_2_6# OAI22X1_5/C OAI22X1_19/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M8992 OAI22X1_19/Y INVX2_72/Y OAI22X1_19/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8993 OAI22X1_19/Y INVX2_104/Y OAI22X1_19/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M8994 OAI22X1_19/a_28_54# INVX2_72/Y OAI22X1_19/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M8995 OAI22X1_19/a_9_54# BUFX2_24/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8996 OAI22X1_19/a_2_6# INVX2_104/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M8997 vdd OAI22X1_5/C OAI22X1_19/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M8998 gnd OR2X1_12/B OAI21X1_52/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M8999 vdd BUFX2_19/A INVX2_226/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9000 INVX2_226/A BUFX2_19/A OAI21X1_52/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9001 INVX2_226/A INVX2_179/Y OAI21X1_52/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9002 OAI21X1_52/a_9_54# OR2X1_12/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9003 OAI21X1_52/a_2_6# INVX2_179/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9004 gnd NAND3X1_7/Y OAI21X1_30/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9005 vdd BUFX2_18/Y INVX2_241/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9006 INVX2_241/A BUFX2_18/Y OAI21X1_30/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9007 INVX2_241/A OAI21X1_30/B OAI21X1_30/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9008 OAI21X1_30/a_9_54# NAND3X1_7/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9009 OAI21X1_30/a_2_6# OAI21X1_30/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9010 gnd INVX2_237/Y OAI21X1_41/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9011 vdd OAI21X1_41/C OAI21X1_41/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9012 OAI21X1_41/Y OAI21X1_41/C OAI21X1_41/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9013 OAI21X1_41/Y OAI21X1_9/B OAI21X1_41/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9014 OAI21X1_41/a_9_54# INVX2_237/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9015 OAI21X1_41/a_2_6# OAI21X1_9/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9016 gnd NOR2X1_72/Y OAI21X1_63/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9017 vdd AOI21X1_3/A OAI21X1_63/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9018 OAI21X1_63/Y AOI21X1_3/A OAI21X1_63/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9019 OAI21X1_63/Y INVX2_88/Y OAI21X1_63/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9020 OAI21X1_63/a_9_54# NOR2X1_72/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9021 OAI21X1_63/a_2_6# INVX2_88/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9022 gnd INVX2_16/Y OAI21X1_74/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9023 vdd OAI21X1_74/C NOR2X1_87/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9024 NOR2X1_87/B OAI21X1_74/C OAI21X1_74/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9025 NOR2X1_87/B INVX2_104/Y OAI21X1_74/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9026 OAI21X1_74/a_9_54# INVX2_16/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9027 OAI21X1_74/a_2_6# INVX2_104/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9028 gnd INVX2_67/Y OAI21X1_96/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9029 vdd OAI21X1_96/C OAI21X1_96/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9030 OAI21X1_96/Y OAI21X1_96/C OAI21X1_96/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9031 OAI21X1_96/Y BUFX2_23/Y OAI21X1_96/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9032 OAI21X1_96/a_9_54# INVX2_67/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9033 OAI21X1_96/a_2_6# BUFX2_23/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9034 gnd INVX2_81/Y OAI21X1_85/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9035 vdd OAI21X1_85/C OAI21X1_85/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9036 OAI21X1_85/Y OAI21X1_85/C OAI21X1_85/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9037 OAI21X1_85/Y BUFX2_22/Y OAI21X1_85/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9038 OAI21X1_85/a_9_54# INVX2_81/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9039 OAI21X1_85/a_2_6# BUFX2_22/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9040 OR2X1_12/a_2_54# OR2X1_12/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9041 OR2X1_12/Y OR2X1_12/a_2_54# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9042 OR2X1_12/Y OR2X1_12/a_2_54# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M9043 vdd OR2X1_12/B OR2X1_12/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9044 OR2X1_12/a_9_54# OR2X1_12/A OR2X1_12/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M9045 gnd OR2X1_12/B OR2X1_12/a_2_54# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9046 AND2X2_11/a_2_6# HAX1_36/YS vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M9047 AND2X2_11/a_9_6# HAX1_36/YS AND2X2_11/a_2_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=100p ps=50u
M9048 AND2X2_11/Y AND2X2_11/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9049 AND2X2_11/Y AND2X2_11/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9050 vdd BUFX2_8/Y AND2X2_11/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9051 gnd BUFX2_8/Y AND2X2_11/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9052 NOR2X1_77/A INVX2_75/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M9053 NAND3X1_22/a_9_6# INVX2_75/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M9054 NOR2X1_77/A INVX2_77/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9055 NOR2X1_77/A INVX2_77/Y NAND3X1_22/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M9056 vdd INVX2_74/Y NOR2X1_77/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9057 NAND3X1_22/a_14_6# INVX2_74/Y NAND3X1_22/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M9058 OR2X1_13/A XNOR2X1_24/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M9059 NAND3X1_11/a_9_6# XNOR2X1_24/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M9060 OR2X1_13/A NOR2X1_69/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9061 OR2X1_13/A NOR2X1_69/Y NAND3X1_11/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M9062 vdd INVX2_0/A OR2X1_13/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9063 NAND3X1_11/a_14_6# INVX2_0/A NAND3X1_11/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M9064 NOR2X1_97/B NAND3X1_44/A vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M9065 NAND3X1_44/a_9_6# NAND3X1_44/A gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M9066 NOR2X1_97/B AOI21X1_6/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9067 NOR2X1_97/B AOI21X1_6/Y NAND3X1_44/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M9068 vdd NAND3X1_44/B NOR2X1_97/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9069 NAND3X1_44/a_14_6# NAND3X1_44/B NAND3X1_44/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M9070 NOR2X1_82/A NOR2X1_90/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M9071 NAND3X1_33/a_9_6# NOR2X1_90/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M9072 NOR2X1_82/A NOR2X1_87/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9073 NOR2X1_82/A NOR2X1_87/Y NAND3X1_33/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M9074 vdd NOR2X1_89/Y NOR2X1_82/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9075 NAND3X1_33/a_14_6# NOR2X1_89/Y NAND3X1_33/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M9076 INVX2_122/A out_state_main[3] vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M9077 NAND3X1_55/a_9_6# out_state_main[3] gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M9078 INVX2_122/A NOR2X1_120/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9079 INVX2_122/A NOR2X1_120/Y NAND3X1_55/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M9080 vdd INVX2_116/Y INVX2_122/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9081 NAND3X1_55/a_14_6# INVX2_116/Y NAND3X1_55/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M9082 FAX1_18/A NOR2X1_9/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9083 FAX1_18/A INVX2_4/Y NOR2X1_11/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9084 NOR2X1_11/a_9_54# NOR2X1_9/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9085 gnd INVX2_4/Y FAX1_18/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9086 FAX1_13/A INVX2_17/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9087 FAX1_13/A NOR2X1_22/B NOR2X1_22/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9088 NOR2X1_22/a_9_54# INVX2_17/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9089 gnd NOR2X1_22/B FAX1_13/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9090 NOR2X1_44/Y NOR2X1_57/B gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9091 NOR2X1_44/Y NOR2X1_47/B NOR2X1_44/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9092 NOR2X1_44/a_9_54# NOR2X1_57/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9093 gnd NOR2X1_47/B NOR2X1_44/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9094 NOR2X1_55/Y NOR2X1_55/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9095 NOR2X1_55/Y NOR2X1_56/B NOR2X1_55/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9096 NOR2X1_55/a_9_54# NOR2X1_55/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9097 gnd NOR2X1_56/B NOR2X1_55/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9098 NOR2X1_33/Y out_temp_data_in[3] gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9099 NOR2X1_33/Y OAI21X1_0/C NOR2X1_33/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9100 NOR2X1_33/a_9_54# out_temp_data_in[3] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9101 gnd OAI21X1_0/C NOR2X1_33/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9102 NOR2X1_66/Y NOR2X1_66/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9103 NOR2X1_66/Y NOR2X1_66/B NOR2X1_66/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9104 NOR2X1_66/a_9_54# NOR2X1_66/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9105 gnd NOR2X1_66/B NOR2X1_66/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9106 NOR2X1_88/Y out_temp_decoded[10] gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9107 NOR2X1_88/Y out_temp_cleared[10] NOR2X1_88/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9108 NOR2X1_88/a_9_54# out_temp_decoded[10] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9109 gnd out_temp_cleared[10] NOR2X1_88/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9110 NOR2X1_77/Y NOR2X1_77/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9111 NOR2X1_77/Y NOR2X1_77/B NOR2X1_77/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9112 NOR2X1_77/a_9_54# NOR2X1_77/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9113 gnd NOR2X1_77/B NOR2X1_77/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9114 NOR2X1_99/Y out_temp_decoded[20] gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9115 NOR2X1_99/Y out_temp_cleared[20] NOR2X1_99/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9116 NOR2X1_99/a_9_54# out_temp_decoded[20] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9117 gnd out_temp_cleared[20] NOR2X1_99/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9118 INVX2_200/Y INVX2_200/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9119 INVX2_200/Y INVX2_200/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9120 INVX2_211/Y INVX2_211/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9121 INVX2_211/Y INVX2_211/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9122 INVX2_222/Y INVX2_222/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9123 INVX2_222/Y INVX2_222/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9124 OAI21X1_9/A INVX2_233/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9125 OAI21X1_9/A INVX2_233/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9126 INVX2_244/Y INVX2_244/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9127 INVX2_244/Y INVX2_244/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9128 INVX2_255/Y INVX2_256/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9129 INVX2_255/Y INVX2_256/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9130 NOR2X1_101/Y out_temp_decoded[24] gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9131 NOR2X1_101/Y out_temp_cleared[24] NOR2X1_101/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9132 NOR2X1_101/a_9_54# out_temp_decoded[24] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9133 gnd out_temp_cleared[24] NOR2X1_101/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9134 OR2X1_16/B OR2X1_16/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9135 OR2X1_16/B out_gameover NOR2X1_123/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9136 NOR2X1_123/a_9_54# OR2X1_16/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9137 gnd out_gameover OR2X1_16/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9138 NOR2X1_112/Y out_temp_data_in[0] gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9139 NOR2X1_112/Y out_temp_data_in[1] NOR2X1_112/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9140 NOR2X1_112/a_9_54# out_temp_data_in[0] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9141 gnd out_temp_data_in[1] NOR2X1_112/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9142 INVX2_90/Y out_temp_cleared[23] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9143 INVX2_90/Y out_temp_cleared[23] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9144 gnd OR2X1_12/B OAI21X1_20/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9145 vdd BUFX2_19/Y INVX2_224/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9146 INVX2_224/A BUFX2_19/Y OAI21X1_20/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9147 INVX2_224/A INVX2_180/Y OAI21X1_20/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9148 OAI21X1_20/a_9_54# OR2X1_12/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9149 OAI21X1_20/a_2_6# INVX2_180/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9150 gnd NOR2X1_66/B OAI21X1_53/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9151 vdd OAI21X1_53/C OAI21X1_53/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9152 OAI21X1_53/Y OAI21X1_53/C OAI21X1_53/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9153 OAI21X1_53/Y OAI21X1_4/A OAI21X1_53/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9154 OAI21X1_53/a_9_54# NOR2X1_66/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9155 OAI21X1_53/a_2_6# OAI21X1_4/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9156 gnd OAI21X1_44/A OAI21X1_42/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9157 vdd BUFX2_18/Y INVX2_237/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9158 INVX2_237/A BUFX2_18/Y OAI21X1_42/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9159 INVX2_237/A OAI21X1_46/B OAI21X1_42/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9160 OAI21X1_42/a_9_54# OAI21X1_44/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9161 OAI21X1_42/a_2_6# OAI21X1_46/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9162 gnd INVX2_242/Y OAI21X1_31/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9163 vdd OAI21X1_31/C OAI21X1_31/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9164 OAI21X1_31/Y OAI21X1_31/C OAI21X1_31/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9165 OAI21X1_31/Y OAI21X1_9/B OAI21X1_31/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9166 OAI21X1_31/a_9_54# INVX2_242/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9167 OAI21X1_31/a_2_6# OAI21X1_9/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9168 gnd INVX2_79/Y OAI21X1_86/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9169 vdd OAI21X1_86/C OAI21X1_86/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9170 OAI21X1_86/Y OAI21X1_86/C OAI21X1_86/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9171 OAI21X1_86/Y BUFX2_22/Y OAI21X1_86/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9172 OAI21X1_86/a_9_54# INVX2_79/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9173 OAI21X1_86/a_2_6# BUFX2_22/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9174 gnd INVX2_6/Y OAI21X1_75/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9175 vdd OAI21X1_75/C NOR2X1_89/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9176 NOR2X1_89/B OAI21X1_75/C OAI21X1_75/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9177 NOR2X1_89/B INVX2_108/Y OAI21X1_75/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9178 OAI21X1_75/a_9_54# INVX2_6/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9179 OAI21X1_75/a_2_6# INVX2_108/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9180 gnd OR2X1_11/A OAI21X1_64/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9181 vdd INVX2_217/A INVX2_256/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9182 INVX2_256/A INVX2_217/A OAI21X1_64/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9183 INVX2_256/A AOI21X1_3/A OAI21X1_64/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9184 OAI21X1_64/a_9_54# OR2X1_11/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9185 OAI21X1_64/a_2_6# AOI21X1_3/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9186 gnd INVX2_66/Y OAI21X1_97/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9187 vdd OAI21X1_97/C OAI21X1_97/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9188 OAI21X1_97/Y OAI21X1_97/C OAI21X1_97/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9189 OAI21X1_97/Y BUFX2_23/Y OAI21X1_97/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9190 OAI21X1_97/a_9_54# INVX2_66/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9191 OAI21X1_97/a_2_6# BUFX2_23/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9192 OR2X1_13/a_2_54# OR2X1_13/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9193 OR2X1_13/Y OR2X1_13/a_2_54# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9194 OR2X1_13/Y OR2X1_13/a_2_54# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M9195 vdd OR2X1_13/B OR2X1_13/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9196 OR2X1_13/a_9_54# OR2X1_13/A OR2X1_13/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M9197 gnd OR2X1_13/B OR2X1_13/a_2_54# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9198 AND2X2_12/a_2_6# HAX1_37/YS vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M9199 AND2X2_12/a_9_6# HAX1_37/YS AND2X2_12/a_2_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=100p ps=50u
M9200 AND2X2_12/Y AND2X2_12/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9201 AND2X2_12/Y AND2X2_12/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9202 vdd BUFX2_6/Y AND2X2_12/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9203 gnd BUFX2_6/Y AND2X2_12/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9204 vdd out_global_score[30] HAX1_0/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M9205 HAX1_0/a_41_74# HAX1_0/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M9206 HAX1_0/a_9_6# out_global_score[30] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M9207 HAX1_0/a_41_74# HAX1_0/B HAX1_0/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M9208 vdd out_global_score[30] HAX1_0/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9209 vdd HAX1_0/a_2_74# HAX1_0/YC vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M9210 HAX1_0/a_38_6# HAX1_0/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9211 HAX1_0/YS HAX1_0/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9212 HAX1_0/a_38_6# out_global_score[30] HAX1_0/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9213 HAX1_0/YS HAX1_0/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M9214 HAX1_0/a_2_74# HAX1_0/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9215 HAX1_0/a_2_74# HAX1_0/B HAX1_0/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9216 HAX1_0/a_49_54# HAX1_0/B HAX1_0/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9217 gnd HAX1_0/a_2_74# HAX1_0/YC Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M9218 NOR2X1_78/B INVX2_69/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M9219 NAND3X1_23/a_9_6# INVX2_69/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M9220 NOR2X1_78/B INVX2_70/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9221 NOR2X1_78/B INVX2_70/Y NAND3X1_23/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M9222 vdd INVX2_68/Y NOR2X1_78/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9223 NAND3X1_23/a_14_6# INVX2_68/Y NAND3X1_23/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M9224 NOR2X1_66/B AND2X2_8/A vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M9225 NAND3X1_12/a_9_6# AND2X2_8/A gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M9226 NOR2X1_66/B INVX2_0/A vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9227 NOR2X1_66/B INVX2_0/A NAND3X1_12/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M9228 vdd INVX2_130/Y NOR2X1_66/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9229 NAND3X1_12/a_14_6# INVX2_130/Y NAND3X1_12/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M9230 NOR2X1_87/A NAND3X1_36/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M9231 NAND3X1_34/a_9_6# NAND3X1_36/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M9232 NOR2X1_87/A NAND3X1_34/C vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9233 NOR2X1_87/A NAND3X1_34/C NAND3X1_34/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M9234 vdd NAND3X1_35/Y NOR2X1_87/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9235 NAND3X1_34/a_14_6# NAND3X1_35/Y NAND3X1_34/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M9236 INVX2_124/A out_alu_done vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M9237 NAND3X1_56/a_9_6# out_alu_done gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M9238 INVX2_124/A out_gameover vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9239 INVX2_124/A out_gameover NAND3X1_56/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M9240 vdd INVX2_123/Y INVX2_124/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9241 NAND3X1_56/a_14_6# INVX2_123/Y NAND3X1_56/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M9242 OAI21X1_80/C OAI22X1_2/D vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M9243 NAND3X1_45/a_9_6# OAI22X1_2/D gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M9244 OAI21X1_80/C INVX2_28/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9245 OAI21X1_80/C INVX2_28/Y NAND3X1_45/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M9246 vdd INVX2_81/Y OAI21X1_80/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9247 NAND3X1_45/a_14_6# INVX2_81/Y NAND3X1_45/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M9248 FAX1_17/A NOR2X1_9/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9249 FAX1_17/A INVX2_17/Y NOR2X1_12/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9250 NOR2X1_12/a_9_54# NOR2X1_9/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9251 gnd INVX2_17/Y FAX1_17/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9252 HAX1_33/B INVX2_1/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9253 HAX1_33/B NOR2X1_27/B NOR2X1_23/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9254 NOR2X1_23/a_9_54# INVX2_1/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9255 gnd NOR2X1_27/B HAX1_33/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9256 NOR2X1_45/Y OR2X1_6/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9257 NOR2X1_45/Y NOR2X1_47/B NOR2X1_45/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9258 NOR2X1_45/a_9_54# OR2X1_6/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9259 gnd NOR2X1_47/B NOR2X1_45/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9260 OAI21X1_0/A out_temp_data_in[1] gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9261 OAI21X1_0/A out_temp_data_in[0] NOR2X1_34/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9262 NOR2X1_34/a_9_54# out_temp_data_in[1] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9263 gnd out_temp_data_in[0] OAI21X1_0/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9264 NOR2X1_67/Y BUFX2_3/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9265 NOR2X1_67/Y BUFX2_8/Y NOR2X1_67/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9266 NOR2X1_67/a_9_54# BUFX2_3/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9267 gnd BUFX2_8/Y NOR2X1_67/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9268 NOR2X1_56/Y INVX2_54/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9269 NOR2X1_56/Y NOR2X1_56/B NOR2X1_56/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9270 NOR2X1_56/a_9_54# INVX2_54/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9271 gnd NOR2X1_56/B NOR2X1_56/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9272 NOR2X1_78/Y NOR2X1_78/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9273 NOR2X1_78/Y NOR2X1_78/B NOR2X1_78/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9274 NOR2X1_78/a_9_54# NOR2X1_78/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9275 gnd NOR2X1_78/B NOR2X1_78/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9276 NOR2X1_89/Y OAI22X1_2/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9277 NOR2X1_89/Y NOR2X1_89/B NOR2X1_89/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9278 NOR2X1_89/a_9_54# OAI22X1_2/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9279 gnd NOR2X1_89/B NOR2X1_89/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9280 INVX2_201/Y INVX2_201/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9281 INVX2_201/Y INVX2_201/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9282 INVX2_212/Y INVX2_212/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9283 INVX2_212/Y INVX2_212/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9284 OAI21X1_3/A OAI21X1_4/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9285 OAI21X1_3/A OAI21X1_4/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9286 INVX2_245/Y INVX2_245/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9287 INVX2_245/Y INVX2_245/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9288 INVX2_234/Y INVX2_234/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9289 INVX2_234/Y INVX2_234/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9290 OR2X1_11/B INVX2_256/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9291 OR2X1_11/B INVX2_256/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9292 gnd HAX1_49/YS MUX2X1_30/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M9293 MUX2X1_30/a_17_50# HAX1_49/A vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M9294 OAI21X1_4/A OR2X1_0/Y MUX2X1_30/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M9295 MUX2X1_30/a_30_54# MUX2X1_30/a_2_10# OAI21X1_4/A vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M9296 MUX2X1_30/a_17_10# HAX1_49/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M9297 vdd OR2X1_0/Y MUX2X1_30/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M9298 MUX2X1_30/a_30_10# OR2X1_0/Y OAI21X1_4/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M9299 gnd OR2X1_0/Y MUX2X1_30/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M9300 vdd HAX1_49/YS MUX2X1_30/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9301 OAI21X1_4/A MUX2X1_30/a_2_10# MUX2X1_30/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9302 NOR2X1_124/Y OR2X1_15/B gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9303 NOR2X1_124/Y NOR2X1_124/B NOR2X1_124/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9304 NOR2X1_124/a_9_54# OR2X1_15/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9305 gnd NOR2X1_124/B NOR2X1_124/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9306 BUFX2_25/A BUFX2_7/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9307 BUFX2_25/A AOI21X1_2/A NOR2X1_102/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9308 NOR2X1_102/a_9_54# BUFX2_7/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9309 gnd AOI21X1_2/A BUFX2_25/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9310 NOR2X1_113/Y OR2X1_6/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9311 NOR2X1_113/Y INVX2_251/Y NOR2X1_113/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9312 NOR2X1_113/a_9_54# OR2X1_6/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9313 gnd INVX2_251/Y NOR2X1_113/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9314 INVX2_91/Y out_temp_cleared[22] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9315 INVX2_91/Y out_temp_cleared[22] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9316 INVX2_80/Y INVX2_80/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9317 INVX2_80/Y INVX2_80/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9318 gnd OAI21X1_6/A OAI21X1_10/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9319 vdd BUFX2_19/Y INVX2_233/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9320 INVX2_233/A BUFX2_19/Y OAI21X1_10/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9321 INVX2_233/A OAI21X1_44/A OAI21X1_10/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9322 OAI21X1_10/a_9_54# OAI21X1_6/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9323 OAI21X1_10/a_2_6# OAI21X1_44/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9324 gnd NOR2X1_66/B OAI21X1_54/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9325 vdd OAI21X1_54/C OAI21X1_54/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9326 OAI21X1_54/Y OAI21X1_54/C OAI21X1_54/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9327 OAI21X1_54/Y OR2X1_12/A OAI21X1_54/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9328 OAI21X1_54/a_9_54# NOR2X1_66/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9329 OAI21X1_54/a_2_6# OR2X1_12/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9330 gnd NAND3X1_7/Y OAI21X1_32/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9331 vdd BUFX2_18/Y INVX2_242/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9332 INVX2_242/A BUFX2_18/Y OAI21X1_32/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9333 INVX2_242/A OAI21X1_32/B OAI21X1_32/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9334 OAI21X1_32/a_9_54# NAND3X1_7/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9335 OAI21X1_32/a_2_6# OAI21X1_32/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9336 gnd INVX2_238/Y OAI21X1_43/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9337 vdd OAI21X1_43/C OAI21X1_43/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9338 OAI21X1_43/Y OAI21X1_43/C OAI21X1_43/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9339 OAI21X1_43/Y OAI21X1_9/B OAI21X1_43/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9340 OAI21X1_43/a_9_54# INVX2_238/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9341 OAI21X1_43/a_2_6# OAI21X1_9/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9342 gnd INVX2_229/Y OAI21X1_21/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9343 vdd OAI21X1_21/C OAI21X1_21/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9344 OAI21X1_21/Y OAI21X1_21/C OAI21X1_21/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9345 OAI21X1_21/Y NOR2X1_66/B OAI21X1_21/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9346 OAI21X1_21/a_9_54# INVX2_229/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9347 OAI21X1_21/a_2_6# NOR2X1_66/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9348 gnd INVX2_78/Y OAI21X1_87/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9349 vdd OAI21X1_87/C OAI21X1_87/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9350 OAI21X1_87/Y OAI21X1_87/C OAI21X1_87/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9351 OAI21X1_87/Y BUFX2_22/Y OAI21X1_87/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9352 OAI21X1_87/a_9_54# INVX2_78/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9353 OAI21X1_87/a_2_6# BUFX2_22/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9354 gnd out_mines[2] OAI21X1_76/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9355 vdd OAI21X1_76/C NOR2X1_90/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9356 NOR2X1_90/A OAI21X1_76/C OAI21X1_76/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9357 NOR2X1_90/A OAI21X1_76/B OAI21X1_76/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9358 OAI21X1_76/a_9_54# out_mines[2] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9359 OAI21X1_76/a_2_6# OAI21X1_76/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9360 gnd OR2X1_11/A OAI21X1_65/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9361 vdd OAI21X1_65/C OAI21X1_65/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9362 OAI21X1_65/Y OAI21X1_65/C OAI21X1_65/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9363 OAI21X1_65/Y AOI21X1_3/A OAI21X1_65/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9364 OAI21X1_65/a_9_54# OR2X1_11/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9365 OAI21X1_65/a_2_6# AOI21X1_3/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9366 gnd INVX2_65/Y OAI21X1_98/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9367 vdd OAI21X1_98/C OAI21X1_98/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9368 OAI21X1_98/Y OAI21X1_98/C OAI21X1_98/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9369 OAI21X1_98/Y BUFX2_23/Y OAI21X1_98/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9370 OAI21X1_98/a_9_54# INVX2_65/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9371 OAI21X1_98/a_2_6# BUFX2_23/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9372 OR2X1_14/a_2_54# OR2X1_14/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9373 OR2X1_14/Y OR2X1_14/a_2_54# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9374 OR2X1_14/Y OR2X1_14/a_2_54# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M9375 vdd OR2X1_14/B OR2X1_14/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9376 OR2X1_14/a_9_54# OR2X1_14/A OR2X1_14/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M9377 gnd OR2X1_14/B OR2X1_14/a_2_54# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9378 AND2X2_13/a_2_6# INVX2_29/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M9379 AND2X2_13/a_9_6# INVX2_29/Y AND2X2_13/a_2_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=100p ps=50u
M9380 AND2X2_13/Y AND2X2_13/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9381 AND2X2_13/Y AND2X2_13/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9382 vdd BUFX2_6/Y AND2X2_13/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9383 gnd BUFX2_6/Y AND2X2_13/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9384 vdd out_global_score[29] HAX1_1/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M9385 HAX1_1/a_41_74# HAX1_1/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M9386 HAX1_1/a_9_6# out_global_score[29] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M9387 HAX1_1/a_41_74# HAX1_1/B HAX1_1/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M9388 vdd out_global_score[29] HAX1_1/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9389 vdd HAX1_1/a_2_74# HAX1_0/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M9390 HAX1_1/a_38_6# HAX1_1/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9391 HAX1_1/YS HAX1_1/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9392 HAX1_1/a_38_6# out_global_score[29] HAX1_1/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9393 HAX1_1/YS HAX1_1/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M9394 HAX1_1/a_2_74# HAX1_1/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9395 HAX1_1/a_2_74# HAX1_1/B HAX1_1/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9396 HAX1_1/a_49_54# HAX1_1/B HAX1_1/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9397 gnd HAX1_1/a_2_74# HAX1_0/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M9398 INVX2_184/A NOR2X1_70/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M9399 NAND3X1_13/a_9_6# NOR2X1_70/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M9400 INVX2_184/A AND2X2_14/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9401 INVX2_184/A AND2X2_14/Y NAND3X1_13/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M9402 vdd INVX2_131/Y INVX2_184/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9403 NAND3X1_13/a_14_6# INVX2_131/Y NAND3X1_13/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M9404 NAND3X1_35/Y INVX2_102/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M9405 NAND3X1_35/a_9_6# INVX2_102/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M9406 NAND3X1_35/Y INVX2_26/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9407 NAND3X1_35/Y INVX2_26/Y NAND3X1_35/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M9408 vdd INVX2_70/Y NAND3X1_35/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9409 NAND3X1_35/a_14_6# INVX2_70/Y NAND3X1_35/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M9410 NOR2X1_78/A INVX2_64/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M9411 NAND3X1_24/a_9_6# INVX2_64/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M9412 NOR2X1_78/A INVX2_65/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9413 NOR2X1_78/A INVX2_65/Y NAND3X1_24/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M9414 vdd INVX2_63/Y NOR2X1_78/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9415 NAND3X1_24/a_14_6# INVX2_63/Y NAND3X1_24/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M9416 NOR2X1_97/A NAND3X1_46/A vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M9417 NAND3X1_46/a_9_6# NAND3X1_46/A gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M9418 NOR2X1_97/A AOI21X1_7/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9419 NOR2X1_97/A AOI21X1_7/Y NAND3X1_46/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M9420 vdd NAND3X1_46/B NOR2X1_97/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9421 NAND3X1_46/a_14_6# NAND3X1_46/B NAND3X1_46/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M9422 NAND3X1_57/Y NOR2X1_121/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M9423 NAND3X1_57/a_9_6# NOR2X1_121/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M9424 NAND3X1_57/Y out_place_done vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9425 NAND3X1_57/Y out_place_done NAND3X1_57/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M9426 vdd in_data_in NAND3X1_57/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9427 NAND3X1_57/a_14_6# in_data_in NAND3X1_57/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M9428 HAX1_30/A INVX2_1/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9429 HAX1_30/A NOR2X1_17/B NOR2X1_13/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9430 NOR2X1_13/a_9_54# INVX2_1/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9431 gnd NOR2X1_17/B HAX1_30/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9432 HAX1_32/A INVX2_2/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9433 HAX1_32/A NOR2X1_27/B NOR2X1_24/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9434 NOR2X1_24/a_9_54# INVX2_2/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9435 gnd NOR2X1_27/B HAX1_32/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9436 NOR2X1_46/Y NOR2X1_55/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9437 NOR2X1_46/Y NOR2X1_47/B NOR2X1_46/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9438 NOR2X1_46/a_9_54# NOR2X1_55/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9439 gnd NOR2X1_47/B NOR2X1_46/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9440 NOR2X1_35/Y NOR2X1_55/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9441 NOR2X1_35/Y NOR2X1_58/A NOR2X1_35/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9442 NOR2X1_35/a_9_54# NOR2X1_55/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9443 gnd NOR2X1_58/A NOR2X1_35/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9444 NOR2X1_68/Y XOR2X1_15/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9445 NOR2X1_68/Y XOR2X1_14/Y NOR2X1_68/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9446 NOR2X1_68/a_9_54# XOR2X1_15/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9447 gnd XOR2X1_14/Y NOR2X1_68/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9448 NOR2X1_57/Y NOR2X1_58/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9449 NOR2X1_57/Y NOR2X1_57/B NOR2X1_57/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9450 NOR2X1_57/a_9_54# NOR2X1_58/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9451 gnd NOR2X1_57/B NOR2X1_57/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9452 NOR2X1_79/Y NOR2X1_79/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9453 NOR2X1_79/Y NOR2X1_79/B NOR2X1_79/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9454 NOR2X1_79/a_9_54# NOR2X1_79/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9455 gnd NOR2X1_79/B NOR2X1_79/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9456 INVX2_202/Y INVX2_202/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9457 INVX2_202/Y INVX2_202/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9458 INVX2_213/Y INVX2_213/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9459 INVX2_213/Y INVX2_213/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9460 MUX2X1_0/B NOR2X1_7/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9461 MUX2X1_0/B NOR2X1_7/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9462 INVX2_224/Y INVX2_224/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9463 INVX2_224/Y INVX2_224/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9464 INVX2_235/Y INVX2_235/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9465 INVX2_235/Y INVX2_235/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9466 INVX2_257/Y OR2X1_11/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9467 INVX2_257/Y OR2X1_11/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9468 gnd HAX1_45/YS MUX2X1_20/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M9469 MUX2X1_20/a_17_50# HAX1_45/A vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M9470 MUX2X1_20/Y OR2X1_2/Y MUX2X1_20/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M9471 MUX2X1_20/a_30_54# MUX2X1_20/a_2_10# MUX2X1_20/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M9472 MUX2X1_20/a_17_10# HAX1_45/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M9473 vdd OR2X1_2/Y MUX2X1_20/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M9474 MUX2X1_20/a_30_10# OR2X1_2/Y MUX2X1_20/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M9475 gnd OR2X1_2/Y MUX2X1_20/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M9476 vdd HAX1_45/YS MUX2X1_20/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9477 MUX2X1_20/Y MUX2X1_20/a_2_10# MUX2X1_20/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9478 gnd HAX1_48/YS MUX2X1_31/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M9479 MUX2X1_31/a_17_50# HAX1_48/A vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M9480 OR2X1_12/A OR2X1_0/Y MUX2X1_31/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M9481 MUX2X1_31/a_30_54# MUX2X1_31/a_2_10# OR2X1_12/A vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M9482 MUX2X1_31/a_17_10# HAX1_48/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M9483 vdd OR2X1_0/Y MUX2X1_31/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M9484 MUX2X1_31/a_30_10# OR2X1_0/Y OR2X1_12/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M9485 gnd OR2X1_0/Y MUX2X1_31/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M9486 vdd HAX1_48/YS MUX2X1_31/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9487 OR2X1_12/A MUX2X1_31/a_2_10# MUX2X1_31/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9488 AOI21X1_2/A INVX2_217/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9489 AOI21X1_2/A BUFX2_7/Y NOR2X1_103/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9490 NOR2X1_103/a_9_54# INVX2_217/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9491 gnd BUFX2_7/Y AOI21X1_2/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9492 NOR2X1_114/Y OR2X1_6/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9493 NOR2X1_114/Y out_temp_data_in[0] NOR2X1_114/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9494 NOR2X1_114/a_9_54# OR2X1_6/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9495 gnd out_temp_data_in[0] NOR2X1_114/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9496 NOR2X1_125/Y INVX2_120/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9497 NOR2X1_125/Y INVX2_117/A NOR2X1_125/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9498 NOR2X1_125/a_9_54# INVX2_120/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9499 gnd INVX2_117/A NOR2X1_125/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9500 NAND2X1_90/Y NOR2X1_46/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M9501 NAND2X1_90/a_9_6# NOR2X1_46/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M9502 vdd BUFX2_21/Y NAND2X1_90/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9503 NAND2X1_90/Y BUFX2_21/Y NAND2X1_90/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9504 INVX2_70/Y out_temp_decoded[11] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9505 INVX2_70/Y out_temp_decoded[11] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9506 INVX2_81/Y out_temp_decoded[3] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9507 INVX2_81/Y out_temp_decoded[3] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9508 INVX2_92/Y out_temp_cleared[21] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9509 INVX2_92/Y out_temp_cleared[21] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9510 gnd INVX2_234/Y OAI21X1_11/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9511 vdd OAI21X1_11/C OAI21X1_11/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9512 OAI21X1_11/Y OAI21X1_11/C OAI21X1_11/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9513 OAI21X1_11/Y OAI21X1_9/B OAI21X1_11/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9514 OAI21X1_11/a_9_54# INVX2_234/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9515 OAI21X1_11/a_2_6# OAI21X1_9/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9516 gnd OAI21X1_44/A OAI21X1_44/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9517 vdd BUFX2_18/Y INVX2_238/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9518 INVX2_238/A BUFX2_18/Y OAI21X1_44/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9519 INVX2_238/A OAI21X1_48/B OAI21X1_44/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9520 OAI21X1_44/a_9_54# OAI21X1_44/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9521 OAI21X1_44/a_2_6# OAI21X1_48/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9522 gnd OAI21X1_8/A OAI21X1_22/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9523 vdd BUFX2_19/Y INVX2_229/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9524 INVX2_229/A BUFX2_19/Y OAI21X1_22/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9525 INVX2_229/A OAI21X1_30/B OAI21X1_22/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9526 OAI21X1_22/a_9_54# OAI21X1_8/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9527 OAI21X1_22/a_2_6# OAI21X1_30/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9528 gnd INVX2_221/Y OAI21X1_33/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9529 vdd OAI21X1_33/C OAI21X1_33/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9530 OAI21X1_33/Y OAI21X1_33/C OAI21X1_33/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9531 OAI21X1_33/Y OAI21X1_9/B OAI21X1_33/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9532 OAI21X1_33/a_9_54# INVX2_221/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9533 OAI21X1_33/a_2_6# OAI21X1_9/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9534 gnd NOR2X1_66/B OAI21X1_55/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9535 vdd OAI21X1_55/C OAI21X1_55/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9536 OAI21X1_55/Y OAI21X1_55/C OAI21X1_55/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9537 OAI21X1_55/Y NAND3X1_9/A OAI21X1_55/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9538 OAI21X1_55/a_9_54# NOR2X1_66/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9539 OAI21X1_55/a_2_6# NAND3X1_9/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9540 gnd INVX2_15/Y OAI21X1_66/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9541 vdd OAI21X1_66/C INVX2_76/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9542 INVX2_76/A OAI21X1_66/C OAI21X1_66/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9543 INVX2_76/A INVX2_74/Y OAI21X1_66/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9544 OAI21X1_66/a_9_54# INVX2_15/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9545 OAI21X1_66/a_2_6# INVX2_74/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9546 gnd out_mines[22] OAI21X1_77/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9547 vdd OAI21X1_77/C AOI21X1_5/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9548 AOI21X1_5/C OAI21X1_77/C OAI21X1_77/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9549 AOI21X1_5/C OAI21X1_77/B OAI21X1_77/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9550 OAI21X1_77/a_9_54# out_mines[22] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9551 OAI21X1_77/a_2_6# OAI21X1_77/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9552 gnd INVX2_77/Y OAI21X1_88/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9553 vdd OAI21X1_88/C OAI21X1_88/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9554 OAI21X1_88/Y OAI21X1_88/C OAI21X1_88/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9555 OAI21X1_88/Y BUFX2_22/Y OAI21X1_88/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9556 OAI21X1_88/a_9_54# INVX2_77/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9557 OAI21X1_88/a_2_6# BUFX2_22/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9558 gnd INVX2_64/Y OAI21X1_99/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9559 vdd OAI21X1_99/C OAI21X1_99/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9560 OAI21X1_99/Y OAI21X1_99/C OAI21X1_99/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9561 OAI21X1_99/Y BUFX2_23/Y OAI21X1_99/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9562 OAI21X1_99/a_9_54# INVX2_64/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9563 OAI21X1_99/a_2_6# BUFX2_23/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9564 OR2X1_15/a_2_54# OR2X1_15/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9565 OR2X1_15/Y OR2X1_15/a_2_54# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9566 OR2X1_15/Y OR2X1_15/a_2_54# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M9567 vdd OR2X1_15/B OR2X1_15/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9568 OR2X1_15/a_9_54# OR2X1_15/A OR2X1_15/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M9569 gnd OR2X1_15/B OR2X1_15/a_2_54# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9570 AND2X2_14/a_2_6# INVX2_132/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M9571 AND2X2_14/a_9_6# INVX2_132/Y AND2X2_14/a_2_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=100p ps=50u
M9572 AND2X2_14/Y AND2X2_14/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9573 AND2X2_14/Y AND2X2_14/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9574 vdd AND2X2_14/B AND2X2_14/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9575 gnd AND2X2_14/B AND2X2_14/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9576 vdd out_global_score[28] HAX1_2/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M9577 HAX1_2/a_41_74# HAX1_2/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M9578 HAX1_2/a_9_6# out_global_score[28] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M9579 HAX1_2/a_41_74# HAX1_2/B HAX1_2/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M9580 vdd out_global_score[28] HAX1_2/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9581 vdd HAX1_2/a_2_74# HAX1_1/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M9582 HAX1_2/a_38_6# HAX1_2/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9583 HAX1_2/YS HAX1_2/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9584 HAX1_2/a_38_6# out_global_score[28] HAX1_2/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9585 HAX1_2/YS HAX1_2/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M9586 HAX1_2/a_2_74# HAX1_2/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9587 HAX1_2/a_2_74# HAX1_2/B HAX1_2/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9588 HAX1_2/a_49_54# HAX1_2/B HAX1_2/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9589 gnd HAX1_2/a_2_74# HAX1_1/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M9590 OAI21X1_59/A INVX2_131/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M9591 NAND3X1_14/a_9_6# INVX2_131/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M9592 OAI21X1_59/A INVX2_132/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9593 OAI21X1_59/A INVX2_132/Y NAND3X1_14/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M9594 vdd INVX2_130/Y OAI21X1_59/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9595 NAND3X1_14/a_14_6# INVX2_130/Y NAND3X1_14/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M9596 NAND3X1_36/Y INVX2_104/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M9597 NAND3X1_36/a_9_6# INVX2_104/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M9598 NAND3X1_36/Y INVX2_16/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9599 NAND3X1_36/Y INVX2_16/Y NAND3X1_36/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M9600 vdd INVX2_72/Y NAND3X1_36/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9601 NAND3X1_36/a_14_6# INVX2_72/Y NAND3X1_36/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M9602 OAI21X1_81/C INVX2_95/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M9603 NAND3X1_47/a_9_6# INVX2_95/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M9604 OAI21X1_81/C INVX2_25/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9605 OAI21X1_81/C INVX2_25/Y NAND3X1_47/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M9606 vdd INVX2_63/Y OAI21X1_81/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9607 NAND3X1_47/a_14_6# INVX2_63/Y NAND3X1_47/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M9608 NOR2X1_79/B INVX2_76/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M9609 NAND3X1_25/a_9_6# INVX2_76/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M9610 NOR2X1_79/B NOR2X1_80/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9611 NOR2X1_79/B NOR2X1_80/Y NAND3X1_25/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M9612 vdd INVX2_80/Y NOR2X1_79/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9613 NAND3X1_25/a_14_6# INVX2_80/Y NAND3X1_25/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M9614 INVX2_123/A out_state_main[2] vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M9615 NAND3X1_58/a_9_6# out_state_main[2] gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M9616 INVX2_123/A NOR2X1_122/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9617 INVX2_123/A NOR2X1_122/Y NAND3X1_58/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M9618 vdd out_state_main[1] INVX2_123/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9619 NAND3X1_58/a_14_6# out_state_main[1] NAND3X1_58/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M9620 HAX1_34/B INVX2_2/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9621 HAX1_34/B NOR2X1_17/B NOR2X1_14/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9622 NOR2X1_14/a_9_54# INVX2_2/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9623 gnd NOR2X1_17/B HAX1_34/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9624 HAX1_31/A INVX2_3/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9625 HAX1_31/A NOR2X1_27/B NOR2X1_25/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9626 NOR2X1_25/a_9_54# INVX2_3/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9627 gnd NOR2X1_27/B HAX1_31/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9628 NOR2X1_36/Y NOR2X1_58/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9629 NOR2X1_36/Y INVX2_54/Y NOR2X1_36/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9630 NOR2X1_36/a_9_54# NOR2X1_58/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9631 gnd INVX2_54/Y NOR2X1_36/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9632 NOR2X1_47/Y INVX2_54/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9633 NOR2X1_47/Y NOR2X1_47/B NOR2X1_47/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9634 NOR2X1_47/a_9_54# INVX2_54/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9635 gnd NOR2X1_47/B NOR2X1_47/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9636 NOR2X1_58/Y NOR2X1_58/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9637 NOR2X1_58/Y OR2X1_6/Y NOR2X1_58/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9638 NOR2X1_58/a_9_54# NOR2X1_58/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9639 gnd OR2X1_6/Y NOR2X1_58/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9640 NOR2X1_69/Y out_start gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9641 NOR2X1_69/Y BUFX2_3/Y NOR2X1_69/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9642 NOR2X1_69/a_9_54# out_start vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9643 gnd BUFX2_3/Y NOR2X1_69/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9644 INVX2_203/Y INVX2_203/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9645 INVX2_203/Y INVX2_203/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9646 INVX2_214/Y INVX2_214/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9647 INVX2_214/Y INVX2_214/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9648 INVX2_225/Y INVX2_225/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9649 INVX2_225/Y INVX2_225/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9650 INVX2_236/Y INVX2_236/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9651 INVX2_236/Y INVX2_236/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9652 OAI21X1_1/A out_temp_data_in[3] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9653 OAI21X1_1/A out_temp_data_in[3] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9654 INVX2_258/Y OR2X1_11/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9655 INVX2_258/Y OR2X1_11/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9656 gnd HAX1_41/YS MUX2X1_10/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M9657 MUX2X1_10/a_17_50# HAX1_41/A vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M9658 MUX2X1_10/Y OR2X1_4/Y MUX2X1_10/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M9659 MUX2X1_10/a_30_54# MUX2X1_10/a_2_10# MUX2X1_10/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M9660 MUX2X1_10/a_17_10# HAX1_41/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M9661 vdd OR2X1_4/Y MUX2X1_10/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M9662 MUX2X1_10/a_30_10# OR2X1_4/Y MUX2X1_10/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M9663 gnd OR2X1_4/Y MUX2X1_10/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M9664 vdd HAX1_41/YS MUX2X1_10/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9665 MUX2X1_10/Y MUX2X1_10/a_2_10# MUX2X1_10/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9666 gnd HAX1_44/YS MUX2X1_21/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M9667 MUX2X1_21/a_17_50# HAX1_44/A vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M9668 MUX2X1_21/Y OR2X1_2/Y MUX2X1_21/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M9669 MUX2X1_21/a_30_54# MUX2X1_21/a_2_10# MUX2X1_21/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M9670 MUX2X1_21/a_17_10# HAX1_44/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M9671 vdd OR2X1_2/Y MUX2X1_21/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M9672 MUX2X1_21/a_30_10# OR2X1_2/Y MUX2X1_21/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M9673 gnd OR2X1_2/Y MUX2X1_21/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M9674 vdd HAX1_44/YS MUX2X1_21/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9675 MUX2X1_21/Y MUX2X1_21/a_2_10# MUX2X1_21/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9676 gnd XNOR2X1_1/Y MUX2X1_32/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M9677 MUX2X1_32/a_17_50# MUX2X1_32/B vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M9678 NOR2X1_66/A OR2X1_0/Y MUX2X1_32/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M9679 MUX2X1_32/a_30_54# MUX2X1_32/a_2_10# NOR2X1_66/A vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M9680 MUX2X1_32/a_17_10# MUX2X1_32/B gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M9681 vdd OR2X1_0/Y MUX2X1_32/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M9682 MUX2X1_32/a_30_10# OR2X1_0/Y NOR2X1_66/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M9683 gnd OR2X1_0/Y MUX2X1_32/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M9684 vdd XNOR2X1_1/Y MUX2X1_32/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9685 NOR2X1_66/A MUX2X1_32/a_2_10# MUX2X1_32/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9686 NOR2X1_115/Y NOR2X1_125/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9687 NOR2X1_115/Y NOR2X1_116/Y NOR2X1_115/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9688 NOR2X1_115/a_9_54# NOR2X1_125/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9689 gnd NOR2X1_116/Y NOR2X1_115/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9690 BUFX2_21/A AND2X2_6/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9691 BUFX2_21/A NOR2X1_104/B NOR2X1_104/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9692 NOR2X1_104/a_9_54# AND2X2_6/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9693 gnd NOR2X1_104/B BUFX2_21/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9694 NAND2X1_91/Y NOR2X1_45/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M9695 NAND2X1_91/a_9_6# NOR2X1_45/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M9696 vdd BUFX2_21/Y NAND2X1_91/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9697 NAND2X1_91/Y BUFX2_21/Y NAND2X1_91/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9698 OAI21X1_93/C NOR2X1_57/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M9699 NAND2X1_80/a_9_6# NOR2X1_57/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M9700 vdd BUFX2_20/Y OAI21X1_93/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9701 OAI21X1_93/C BUFX2_20/Y NAND2X1_80/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9702 INVX2_71/Y out_temp_decoded[10] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9703 INVX2_71/Y out_temp_decoded[10] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9704 INVX2_60/Y out_temp_decoded[20] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9705 INVX2_60/Y out_temp_decoded[20] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9706 INVX2_82/Y out_temp_decoded[2] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9707 INVX2_82/Y out_temp_decoded[2] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9708 INVX2_93/Y out_temp_cleared[20] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9709 INVX2_93/Y out_temp_cleared[20] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9710 gnd OAI21X1_8/B OAI21X1_12/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9711 vdd BUFX2_19/Y INVX2_234/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9712 INVX2_234/A BUFX2_19/Y OAI21X1_12/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9713 INVX2_234/A OAI21X1_44/A OAI21X1_12/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9714 OAI21X1_12/a_9_54# OAI21X1_8/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9715 OAI21X1_12/a_2_6# OAI21X1_44/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9716 gnd NAND3X1_8/Y OAI21X1_34/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9717 vdd BUFX2_18/Y INVX2_221/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9718 INVX2_221/A BUFX2_18/Y OAI21X1_34/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9719 INVX2_221/A INVX2_181/Y OAI21X1_34/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9720 OAI21X1_34/a_9_54# NAND3X1_8/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9721 OAI21X1_34/a_2_6# INVX2_181/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9722 gnd INVX2_243/Y OAI21X1_45/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9723 vdd OAI21X1_45/C OAI21X1_45/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9724 OAI21X1_45/Y OAI21X1_45/C OAI21X1_45/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9725 OAI21X1_45/Y OAI21X1_9/B OAI21X1_45/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9726 OAI21X1_45/a_9_54# INVX2_243/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9727 OAI21X1_45/a_2_6# OAI21X1_9/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9728 gnd INVX2_230/Y OAI21X1_23/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9729 vdd OAI21X1_23/C OAI21X1_23/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9730 OAI21X1_23/Y OAI21X1_23/C OAI21X1_23/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9731 OAI21X1_23/Y NOR2X1_66/B OAI21X1_23/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9732 OAI21X1_23/a_9_54# INVX2_230/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9733 OAI21X1_23/a_2_6# NOR2X1_66/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9734 gnd NOR2X1_66/B OAI21X1_56/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9735 vdd OAI21X1_56/C OAI21X1_56/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9736 OAI21X1_56/Y OAI21X1_56/C OAI21X1_56/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9737 OAI21X1_56/Y NOR2X1_63/B OAI21X1_56/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9738 OAI21X1_56/a_9_54# NOR2X1_66/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9739 OAI21X1_56/a_2_6# NOR2X1_63/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9740 gnd INVX2_16/Y OAI21X1_67/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9741 vdd OAI21X1_67/C INVX2_73/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9742 INVX2_73/A OAI21X1_67/C OAI21X1_67/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9743 INVX2_73/A INVX2_72/Y OAI21X1_67/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9744 OAI21X1_67/a_9_54# INVX2_16/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9745 OAI21X1_67/a_2_6# INVX2_72/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9746 gnd INVX2_11/Y OAI21X1_78/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9747 vdd OAI21X1_78/C NOR2X1_94/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9748 NOR2X1_94/B OAI21X1_78/C OAI21X1_78/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9749 NOR2X1_94/B INVX2_98/Y OAI21X1_78/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9750 OAI21X1_78/a_9_54# INVX2_11/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9751 OAI21X1_78/a_2_6# INVX2_98/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9752 gnd INVX2_75/Y OAI21X1_89/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9753 vdd OAI21X1_89/C OAI21X1_89/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9754 OAI21X1_89/Y OAI21X1_89/C OAI21X1_89/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9755 OAI21X1_89/Y BUFX2_22/Y OAI21X1_89/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9756 OAI21X1_89/a_9_54# INVX2_75/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9757 OAI21X1_89/a_2_6# BUFX2_22/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9758 OR2X1_16/a_2_54# OR2X1_16/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9759 OR2X1_16/Y OR2X1_16/a_2_54# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9760 OR2X1_16/Y OR2X1_16/a_2_54# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M9761 vdd OR2X1_16/B OR2X1_16/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9762 OR2X1_16/a_9_54# OR2X1_16/A OR2X1_16/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M9763 gnd OR2X1_16/B OR2X1_16/a_2_54# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9764 AND2X2_15/a_2_6# NOR2X1_78/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M9765 AND2X2_15/a_9_6# NOR2X1_78/Y AND2X2_15/a_2_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=100p ps=50u
M9766 AND2X2_15/Y AND2X2_15/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9767 AND2X2_15/Y AND2X2_15/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9768 vdd NOR2X1_77/Y AND2X2_15/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9769 gnd NOR2X1_77/Y AND2X2_15/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9770 vdd out_global_score[27] HAX1_3/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M9771 HAX1_3/a_41_74# HAX1_3/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M9772 HAX1_3/a_9_6# out_global_score[27] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M9773 HAX1_3/a_41_74# HAX1_3/B HAX1_3/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M9774 vdd out_global_score[27] HAX1_3/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9775 vdd HAX1_3/a_2_74# HAX1_2/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M9776 HAX1_3/a_38_6# HAX1_3/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9777 HAX1_3/YS HAX1_3/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9778 HAX1_3/a_38_6# out_global_score[27] HAX1_3/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9779 HAX1_3/YS HAX1_3/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M9780 HAX1_3/a_2_74# HAX1_3/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9781 HAX1_3/a_2_74# HAX1_3/B HAX1_3/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9782 HAX1_3/a_49_54# HAX1_3/B HAX1_3/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9783 gnd HAX1_3/a_2_74# HAX1_2/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M9784 NOR2X1_79/A AOI21X1_4/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M9785 NAND3X1_26/a_9_6# AOI21X1_4/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M9786 NOR2X1_79/A NOR2X1_81/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9787 NOR2X1_79/A NOR2X1_81/Y NAND3X1_26/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M9788 vdd INVX2_62/Y NOR2X1_79/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9789 NAND3X1_26/a_14_6# INVX2_62/Y NAND3X1_26/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M9790 OAI22X1_5/C AND2X2_14/B vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M9791 NAND3X1_48/a_9_6# AND2X2_14/B gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M9792 OAI22X1_5/C out_alu vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9793 OAI22X1_5/C out_alu NAND3X1_48/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M9794 vdd INVX2_131/Y OAI22X1_5/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9795 NAND3X1_48/a_14_6# INVX2_131/Y NAND3X1_48/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M9796 INVX2_86/A AND2X2_15/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M9797 NAND3X1_15/a_9_6# AND2X2_15/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M9798 INVX2_86/A NOR2X1_71/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9799 INVX2_86/A NOR2X1_71/Y NAND3X1_15/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M9800 vdd INVX2_84/Y INVX2_86/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9801 NAND3X1_15/a_14_6# INVX2_84/Y NAND3X1_15/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M9802 OAI21X1_75/C OAI22X1_3/D vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M9803 NAND3X1_37/a_9_6# OAI22X1_3/D gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M9804 OAI21X1_75/C INVX2_9/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9805 OAI21X1_75/C INVX2_9/Y NAND3X1_37/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M9806 vdd INVX2_85/Y OAI21X1_75/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9807 NAND3X1_37/a_14_6# INVX2_85/Y NAND3X1_37/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M9808 FAX1_18/B INVX2_3/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9809 FAX1_18/B NOR2X1_17/B NOR2X1_15/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9810 NOR2X1_15/a_9_54# INVX2_3/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9811 gnd NOR2X1_17/B FAX1_18/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9812 FAX1_13/C INVX2_4/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9813 FAX1_13/C NOR2X1_27/B NOR2X1_26/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9814 NOR2X1_26/a_9_54# INVX2_4/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9815 gnd NOR2X1_27/B FAX1_13/C Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9816 NOR2X1_37/Y NOR2X1_40/B gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9817 NOR2X1_37/Y NOR2X1_57/B NOR2X1_37/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9818 NOR2X1_37/a_9_54# NOR2X1_40/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9819 gnd NOR2X1_57/B NOR2X1_37/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9820 NOR2X1_59/Y INVX2_54/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9821 NOR2X1_59/Y NOR2X1_59/B NOR2X1_59/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9822 NOR2X1_59/a_9_54# INVX2_54/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9823 gnd NOR2X1_59/B NOR2X1_59/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9824 NOR2X1_48/Y NOR2X1_55/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9825 NOR2X1_48/Y NOR2X1_59/B NOR2X1_48/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9826 NOR2X1_48/a_9_54# NOR2X1_55/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9827 gnd NOR2X1_59/B NOR2X1_48/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9828 INVX2_204/Y INVX2_204/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9829 INVX2_204/Y INVX2_204/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9830 INVX2_215/Y INVX2_215/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9831 INVX2_215/Y INVX2_215/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9832 BUFX2_8/A NOR2X1_66/B gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9833 BUFX2_8/A NOR2X1_66/B vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9834 INVX2_226/Y INVX2_226/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9835 INVX2_226/Y INVX2_226/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9836 INVX2_237/Y INVX2_237/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9837 INVX2_237/Y INVX2_237/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9838 INVX2_259/Y INVX1_0/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9839 INVX2_259/Y INVX1_0/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9840 gnd HAX1_40/YS MUX2X1_11/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M9841 MUX2X1_11/a_17_50# HAX1_40/A vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M9842 MUX2X1_11/Y OR2X1_4/Y MUX2X1_11/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M9843 MUX2X1_11/a_30_54# MUX2X1_11/a_2_10# MUX2X1_11/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M9844 MUX2X1_11/a_17_10# HAX1_40/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M9845 vdd OR2X1_4/Y MUX2X1_11/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M9846 MUX2X1_11/a_30_10# OR2X1_4/Y MUX2X1_11/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M9847 gnd OR2X1_4/Y MUX2X1_11/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M9848 vdd HAX1_40/YS MUX2X1_11/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9849 MUX2X1_11/Y MUX2X1_11/a_2_10# MUX2X1_11/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9850 gnd XNOR2X1_5/Y MUX2X1_22/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M9851 MUX2X1_22/a_17_50# MUX2X1_22/B vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M9852 MUX2X1_22/Y OR2X1_2/Y MUX2X1_22/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M9853 MUX2X1_22/a_30_54# MUX2X1_22/a_2_10# MUX2X1_22/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M9854 MUX2X1_22/a_17_10# MUX2X1_22/B gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M9855 vdd OR2X1_2/Y MUX2X1_22/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M9856 MUX2X1_22/a_30_10# OR2X1_2/Y MUX2X1_22/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M9857 gnd OR2X1_2/Y MUX2X1_22/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M9858 vdd XNOR2X1_5/Y MUX2X1_22/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9859 MUX2X1_22/Y MUX2X1_22/a_2_10# MUX2X1_22/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9860 gnd XNOR2X1_0/Y MUX2X1_33/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M9861 MUX2X1_33/a_17_50# NOR2X1_0/A vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M9862 NAND3X1_9/A OR2X1_0/Y MUX2X1_33/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M9863 MUX2X1_33/a_30_54# MUX2X1_33/a_2_10# NAND3X1_9/A vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M9864 MUX2X1_33/a_17_10# NOR2X1_0/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M9865 vdd OR2X1_0/Y MUX2X1_33/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M9866 MUX2X1_33/a_30_10# OR2X1_0/Y NAND3X1_9/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M9867 gnd OR2X1_0/Y MUX2X1_33/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M9868 vdd XNOR2X1_0/Y MUX2X1_33/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9869 NAND3X1_9/A MUX2X1_33/a_2_10# MUX2X1_33/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9870 AND2X2_14/B out_load gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9871 AND2X2_14/B BUFX2_3/Y NOR2X1_105/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9872 NOR2X1_105/a_9_54# out_load vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9873 gnd BUFX2_3/Y AND2X2_14/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9874 NOR2X1_116/Y INVX2_119/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M9875 NOR2X1_116/Y INVX2_120/A NOR2X1_116/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M9876 NOR2X1_116/a_9_54# INVX2_119/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9877 gnd INVX2_120/A NOR2X1_116/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9878 OAI21X1_83/C NOR2X1_48/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M9879 NAND2X1_70/a_9_6# NOR2X1_48/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M9880 vdd BUFX2_20/Y OAI21X1_83/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9881 OAI21X1_83/C BUFX2_20/Y NAND2X1_70/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9882 NAND2X1_92/Y NOR2X1_44/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M9883 NAND2X1_92/a_9_6# NOR2X1_44/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M9884 vdd BUFX2_21/Y NAND2X1_92/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9885 NAND2X1_92/Y BUFX2_21/Y NAND2X1_92/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9886 OAI21X1_94/C NOR2X1_56/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M9887 NAND2X1_81/a_9_6# NOR2X1_56/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M9888 vdd BUFX2_20/Y OAI21X1_94/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9889 OAI21X1_94/C BUFX2_20/Y NAND2X1_81/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9890 INVX2_72/Y out_temp_decoded[9] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9891 INVX2_72/Y out_temp_decoded[9] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9892 INVX2_61/Y out_temp_decoded[19] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9893 INVX2_61/Y out_temp_decoded[19] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9894 INVX2_50/Y INVX2_50/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9895 INVX2_50/Y INVX2_50/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9896 INVX2_94/Y out_temp_cleared[19] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9897 INVX2_94/Y out_temp_cleared[19] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9898 INVX2_83/Y out_temp_decoded[1] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9899 INVX2_83/Y out_temp_decoded[1] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9900 gnd INVX2_239/Y OAI21X1_13/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9901 vdd OAI21X1_13/C OAI21X1_13/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9902 OAI21X1_13/Y OAI21X1_13/C OAI21X1_13/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9903 OAI21X1_13/Y OAI21X1_9/B OAI21X1_13/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9904 OAI21X1_13/a_9_54# INVX2_239/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9905 OAI21X1_13/a_2_6# OAI21X1_9/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9906 gnd INVX2_225/Y OAI21X1_35/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9907 vdd OAI21X1_35/C OAI21X1_35/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9908 OAI21X1_35/Y OAI21X1_35/C OAI21X1_35/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9909 OAI21X1_35/Y OAI21X1_9/B OAI21X1_35/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9910 OAI21X1_35/a_9_54# INVX2_225/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9911 OAI21X1_35/a_2_6# OAI21X1_9/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9912 gnd OAI21X1_8/A OAI21X1_24/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9913 vdd BUFX2_19/Y INVX2_230/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9914 INVX2_230/A BUFX2_19/Y OAI21X1_24/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9915 INVX2_230/A OAI21X1_32/B OAI21X1_24/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9916 OAI21X1_24/a_9_54# OAI21X1_8/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9917 OAI21X1_24/a_2_6# OAI21X1_32/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9918 gnd NAND3X1_7/Y OAI21X1_46/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9919 vdd BUFX2_18/Y INVX2_243/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9920 INVX2_243/A BUFX2_18/Y OAI21X1_46/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9921 INVX2_243/A OAI21X1_46/B OAI21X1_46/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9922 OAI21X1_46/a_9_54# NAND3X1_7/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9923 OAI21X1_46/a_2_6# OAI21X1_46/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9924 gnd INVX2_21/Y OAI21X1_68/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9925 vdd OAI21X1_68/C INVX2_62/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9926 INVX2_62/A OAI21X1_68/C OAI21X1_68/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9927 INVX2_62/A INVX2_60/Y OAI21X1_68/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9928 OAI21X1_68/a_9_54# INVX2_21/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9929 OAI21X1_68/a_2_6# INVX2_60/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9930 gnd INVX2_0/Y OAI21X1_57/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9931 vdd AND2X2_8/B OAI21X1_57/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9932 OAI21X1_57/Y AND2X2_8/B OAI21X1_57/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9933 OAI21X1_57/Y OAI21X1_57/B OAI21X1_57/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9934 OAI21X1_57/a_9_54# INVX2_0/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9935 OAI21X1_57/a_2_6# OAI21X1_57/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9936 gnd out_mines[16] OAI21X1_79/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M9937 vdd OAI21X1_79/C NOR2X1_94/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M9938 NOR2X1_94/A OAI21X1_79/C OAI21X1_79/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9939 NOR2X1_94/A OAI21X1_79/B OAI21X1_79/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9940 OAI21X1_79/a_9_54# out_mines[16] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9941 OAI21X1_79/a_2_6# OAI21X1_79/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9942 AND2X2_16/a_2_6# AND2X2_16/A vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M9943 AND2X2_16/a_9_6# AND2X2_16/A AND2X2_16/a_2_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=100p ps=50u
M9944 AND2X2_16/Y AND2X2_16/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9945 AND2X2_16/Y AND2X2_16/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9946 vdd AND2X2_16/B AND2X2_16/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9947 gnd AND2X2_16/B AND2X2_16/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9948 gnd NOR2X1_0/A XNOR2X1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M9949 XNOR2X1_0/Y NOR2X1_0/A XNOR2X1_0/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M9950 XNOR2X1_0/a_12_41# NOR2X1_0/B gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9951 XNOR2X1_0/a_18_54# XNOR2X1_0/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M9952 XNOR2X1_0/a_35_6# XNOR2X1_0/a_2_6# XNOR2X1_0/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M9953 XNOR2X1_0/a_18_6# XNOR2X1_0/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9954 vdd NOR2X1_0/A XNOR2X1_0/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M9955 vdd NOR2X1_0/B XNOR2X1_0/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9956 XNOR2X1_0/Y XNOR2X1_0/a_2_6# XNOR2X1_0/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M9957 XNOR2X1_0/a_35_54# NOR2X1_0/A XNOR2X1_0/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9958 XNOR2X1_0/a_12_41# NOR2X1_0/B vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9959 gnd NOR2X1_0/B XNOR2X1_0/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9960 INVX1_0/Y in_clkb vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=100p ps=50u
M9961 INVX1_0/Y in_clkb gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=50p ps=30u
M9962 DFFNEGX1_90/a_76_6# BUFX2_11/Y DFFNEGX1_90/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M9963 gnd BUFX2_11/Y DFFNEGX1_90/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M9964 DFFNEGX1_90/a_66_6# DFFNEGX1_90/a_2_6# DFFNEGX1_90/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M9965 out_temp_cleared[1] DFFNEGX1_90/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9966 DFFNEGX1_90/a_23_6# BUFX2_11/Y DFFNEGX1_90/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M9967 DFFNEGX1_90/a_23_6# DFFNEGX1_90/a_2_6# DFFNEGX1_90/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M9968 gnd DFFNEGX1_90/a_34_4# DFFNEGX1_90/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M9969 vdd DFFNEGX1_90/a_34_4# DFFNEGX1_90/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M9970 DFFNEGX1_90/a_61_74# DFFNEGX1_90/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M9971 DFFNEGX1_90/a_34_4# DFFNEGX1_90/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9972 DFFNEGX1_90/a_34_4# DFFNEGX1_90/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M9973 vdd out_temp_cleared[1] DFFNEGX1_90/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M9974 gnd out_temp_cleared[1] DFFNEGX1_90/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9975 DFFNEGX1_90/a_61_6# DFFNEGX1_90/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9976 DFFNEGX1_90/a_76_84# DFFNEGX1_90/a_2_6# DFFNEGX1_90/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M9977 out_temp_cleared[1] DFFNEGX1_90/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M9978 vdd BUFX2_11/Y DFFNEGX1_90/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M9979 DFFNEGX1_90/a_31_6# DFFNEGX1_90/a_2_6# DFFNEGX1_90/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9980 DFFNEGX1_90/a_66_6# BUFX2_11/Y DFFNEGX1_90/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9981 DFFNEGX1_90/a_17_74# OAI22X1_27/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9982 DFFNEGX1_90/a_31_74# BUFX2_11/Y DFFNEGX1_90/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9983 DFFNEGX1_90/a_17_6# OAI22X1_27/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M9984 vdd out_global_score[26] HAX1_4/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M9985 HAX1_4/a_41_74# HAX1_4/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M9986 HAX1_4/a_9_6# out_global_score[26] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M9987 HAX1_4/a_41_74# HAX1_4/B HAX1_4/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M9988 vdd out_global_score[26] HAX1_4/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M9989 vdd HAX1_4/a_2_74# HAX1_3/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M9990 HAX1_4/a_38_6# HAX1_4/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9991 HAX1_4/YS HAX1_4/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9992 HAX1_4/a_38_6# out_global_score[26] HAX1_4/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9993 HAX1_4/YS HAX1_4/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M9994 HAX1_4/a_2_74# HAX1_4/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M9995 HAX1_4/a_2_74# HAX1_4/B HAX1_4/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M9996 HAX1_4/a_49_54# HAX1_4/B HAX1_4/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M9997 gnd HAX1_4/a_2_74# HAX1_3/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M9998 AND2X2_0/a_2_6# XOR2X1_7/A vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M9999 AND2X2_0/a_9_6# XOR2X1_7/A AND2X2_0/a_2_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=100p ps=50u
M10000 XOR2X1_6/A AND2X2_0/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10001 XOR2X1_6/A AND2X2_0/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10002 vdd FAX1_5/YS AND2X2_0/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10003 gnd FAX1_5/YS AND2X2_0/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10004 AOI21X1_3/A NOR2X1_97/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M10005 NAND3X1_27/a_9_6# NOR2X1_97/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M10006 AOI21X1_3/A NOR2X1_82/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10007 AOI21X1_3/A NOR2X1_82/Y NAND3X1_27/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M10008 vdd NOR2X1_91/Y AOI21X1_3/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10009 NAND3X1_27/a_14_6# NOR2X1_91/Y NAND3X1_27/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M10010 OAI21X1_76/C OAI22X1_3/B vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M10011 NAND3X1_38/a_9_6# OAI22X1_3/B gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M10012 OAI21X1_76/C INVX2_10/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10013 OAI21X1_76/C INVX2_10/Y NAND3X1_38/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M10014 vdd INVX2_83/Y OAI21X1_76/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10015 NAND3X1_38/a_14_6# INVX2_83/Y NAND3X1_38/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M10016 INVX2_87/A INVX2_85/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M10017 NAND3X1_16/a_9_6# INVX2_85/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M10018 INVX2_87/A NOR2X1_73/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10019 INVX2_87/A NOR2X1_73/Y NAND3X1_16/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M10020 vdd INVX2_79/Y INVX2_87/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10021 NAND3X1_16/a_14_6# INVX2_79/Y NAND3X1_16/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M10022 NAND3X1_49/Y INVX2_121/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M10023 NAND3X1_49/a_9_6# INVX2_121/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M10024 NAND3X1_49/Y INVX2_127/A vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10025 NAND3X1_49/Y INVX2_127/A NAND3X1_49/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M10026 vdd NOR2X1_125/Y NAND3X1_49/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10027 NAND3X1_49/a_14_6# NOR2X1_125/Y NAND3X1_49/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M10028 FAX1_17/C INVX2_4/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M10029 FAX1_17/C NOR2X1_17/B NOR2X1_16/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M10030 NOR2X1_16/a_9_54# INVX2_4/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10031 gnd NOR2X1_17/B FAX1_17/C Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10032 FAX1_11/A INVX2_17/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M10033 FAX1_11/A NOR2X1_27/B NOR2X1_27/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M10034 NOR2X1_27/a_9_54# INVX2_17/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10035 gnd NOR2X1_27/B FAX1_11/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10036 NOR2X1_38/Y NOR2X1_40/B gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M10037 NOR2X1_38/Y OR2X1_6/Y NOR2X1_38/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M10038 NOR2X1_38/a_9_54# NOR2X1_40/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10039 gnd OR2X1_6/Y NOR2X1_38/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10040 NOR2X1_49/Y NOR2X1_57/B gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M10041 NOR2X1_49/Y NOR2X1_52/B NOR2X1_49/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M10042 NOR2X1_49/a_9_54# NOR2X1_57/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10043 gnd NOR2X1_52/B NOR2X1_49/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10044 INVX2_205/Y INVX2_205/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10045 INVX2_205/Y INVX2_205/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10046 INVX2_216/Y INVX2_216/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10047 INVX2_216/Y INVX2_216/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10048 OAI21X1_5/A OAI21X1_6/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10049 OAI21X1_5/A OAI21X1_6/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10050 INVX2_238/Y INVX2_238/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10051 INVX2_238/Y INVX2_238/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10052 BUFX2_7/A OAI22X1_5/C gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10053 BUFX2_7/A OAI22X1_5/C vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10054 gnd XNOR2X1_9/Y MUX2X1_12/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M10055 MUX2X1_12/a_17_50# MUX2X1_12/B vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M10056 MUX2X1_12/Y OR2X1_4/Y MUX2X1_12/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M10057 MUX2X1_12/a_30_54# MUX2X1_12/a_2_10# MUX2X1_12/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M10058 MUX2X1_12/a_17_10# MUX2X1_12/B gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10059 vdd OR2X1_4/Y MUX2X1_12/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M10060 MUX2X1_12/a_30_10# OR2X1_4/Y MUX2X1_12/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M10061 gnd OR2X1_4/Y MUX2X1_12/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M10062 vdd XNOR2X1_9/Y MUX2X1_12/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10063 MUX2X1_12/Y MUX2X1_12/a_2_10# MUX2X1_12/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10064 gnd XNOR2X1_4/Y MUX2X1_23/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M10065 MUX2X1_23/a_17_50# NOR2X1_2/A vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M10066 XNOR2X1_3/A OR2X1_2/Y MUX2X1_23/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M10067 MUX2X1_23/a_30_54# MUX2X1_23/a_2_10# XNOR2X1_3/A vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M10068 MUX2X1_23/a_17_10# NOR2X1_2/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10069 vdd OR2X1_2/Y MUX2X1_23/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M10070 MUX2X1_23/a_30_10# OR2X1_2/Y XNOR2X1_3/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M10071 gnd OR2X1_2/Y MUX2X1_23/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M10072 vdd XNOR2X1_4/Y MUX2X1_23/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10073 XNOR2X1_3/A MUX2X1_23/a_2_10# MUX2X1_23/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10074 gnd MUX2X1_34/A MUX2X1_34/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M10075 MUX2X1_34/a_17_50# NOR2X1_0/B vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M10076 NOR2X1_63/B OR2X1_0/Y MUX2X1_34/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M10077 MUX2X1_34/a_30_54# MUX2X1_34/a_2_10# NOR2X1_63/B vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M10078 MUX2X1_34/a_17_10# NOR2X1_0/B gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10079 vdd OR2X1_0/Y MUX2X1_34/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M10080 MUX2X1_34/a_30_10# OR2X1_0/Y NOR2X1_63/B Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M10081 gnd OR2X1_0/Y MUX2X1_34/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M10082 vdd MUX2X1_34/A MUX2X1_34/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10083 NOR2X1_63/B MUX2X1_34/a_2_10# MUX2X1_34/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10084 INVX2_217/A BUFX2_3/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M10085 INVX2_217/A NOR2X1_107/Y NOR2X1_106/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M10086 NOR2X1_106/a_9_54# BUFX2_3/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10087 gnd NOR2X1_107/Y INVX2_217/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10088 NOR2X1_117/Y out_state_main[3] gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M10089 NOR2X1_117/Y INVX2_125/Y NOR2X1_117/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M10090 NOR2X1_117/a_9_54# out_state_main[3] vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10091 gnd INVX2_125/Y NOR2X1_117/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10092 OAI21X1_62/B NOR2X1_79/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M10093 NAND2X1_60/a_9_6# NOR2X1_79/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10094 vdd BUFX2_7/Y OAI21X1_62/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10095 OAI21X1_62/B BUFX2_7/Y NAND2X1_60/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10096 OAI21X1_95/C NOR2X1_55/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M10097 NAND2X1_82/a_9_6# NOR2X1_55/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10098 vdd BUFX2_21/Y OAI21X1_95/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10099 OAI21X1_95/C BUFX2_21/Y NAND2X1_82/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10100 NAND2X1_93/Y NOR2X1_43/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M10101 NAND2X1_93/a_9_6# NOR2X1_43/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10102 vdd BUFX2_21/Y NAND2X1_93/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10103 NAND2X1_93/Y BUFX2_21/Y NAND2X1_93/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10104 OAI21X1_84/C NOR2X1_42/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M10105 NAND2X1_71/a_9_6# NOR2X1_42/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10106 vdd BUFX2_20/Y OAI21X1_84/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10107 OAI21X1_84/C BUFX2_20/Y NAND2X1_71/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10108 INVX2_51/Y INVX2_51/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10109 INVX2_51/Y INVX2_51/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10110 INVX2_73/Y INVX2_73/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10111 INVX2_73/Y INVX2_73/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10112 INVX2_62/Y INVX2_62/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10113 INVX2_62/Y INVX2_62/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10114 INVX2_40/Y INVX2_40/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10115 INVX2_40/Y INVX2_40/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10116 INVX2_95/Y out_temp_cleared[18] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10117 INVX2_95/Y out_temp_cleared[18] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10118 INVX2_84/Y INVX2_84/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10119 INVX2_84/Y INVX2_84/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10120 gnd OAI21X1_6/A OAI21X1_14/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M10121 vdd BUFX2_19/Y INVX2_239/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M10122 INVX2_239/A BUFX2_19/Y OAI21X1_14/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10123 INVX2_239/A NAND3X1_7/Y OAI21X1_14/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M10124 OAI21X1_14/a_9_54# OAI21X1_6/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10125 OAI21X1_14/a_2_6# NAND3X1_7/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10126 gnd INVX2_235/Y OAI21X1_25/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M10127 vdd OAI21X1_25/C OAI21X1_25/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M10128 OAI21X1_25/Y OAI21X1_25/C OAI21X1_25/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10129 OAI21X1_25/Y NOR2X1_66/B OAI21X1_25/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M10130 OAI21X1_25/a_9_54# INVX2_235/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10131 OAI21X1_25/a_2_6# NOR2X1_66/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10132 gnd OR2X1_12/B OAI21X1_36/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M10133 vdd BUFX2_18/Y INVX2_225/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M10134 INVX2_225/A BUFX2_18/Y OAI21X1_36/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10135 INVX2_225/A INVX2_181/Y OAI21X1_36/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M10136 OAI21X1_36/a_9_54# OR2X1_12/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10137 OAI21X1_36/a_2_6# INVX2_181/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10138 gnd INVX2_244/Y OAI21X1_47/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M10139 vdd OAI21X1_47/C OAI21X1_47/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M10140 OAI21X1_47/Y OAI21X1_47/C OAI21X1_47/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10141 OAI21X1_47/Y OAI21X1_9/B OAI21X1_47/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M10142 OAI21X1_47/a_9_54# INVX2_244/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10143 OAI21X1_47/a_2_6# OAI21X1_9/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10144 gnd INVX2_22/Y OAI21X1_69/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M10145 vdd OAI21X1_69/C NOR2X1_84/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M10146 NOR2X1_84/A OAI21X1_69/C OAI21X1_69/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10147 NOR2X1_84/A INVX2_64/Y OAI21X1_69/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M10148 OAI21X1_69/a_9_54# INVX2_22/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10149 OAI21X1_69/a_2_6# INVX2_64/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10150 gnd out_start OAI21X1_58/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M10151 vdd OAI21X1_58/C OAI21X1_58/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M10152 OAI21X1_58/Y OAI21X1_58/C OAI21X1_58/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10153 OAI21X1_58/Y OR2X1_11/A OAI21X1_58/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M10154 OAI21X1_58/a_9_54# out_start vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10155 OAI21X1_58/a_2_6# OR2X1_11/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10156 AND2X2_17/a_2_6# AND2X2_17/A vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M10157 AND2X2_17/a_9_6# AND2X2_17/A AND2X2_17/a_2_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=100p ps=50u
M10158 AND2X2_17/Y AND2X2_17/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10159 AND2X2_17/Y AND2X2_17/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10160 vdd OR2X1_15/Y AND2X2_17/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10161 gnd OR2X1_15/Y AND2X2_17/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10162 gnd XNOR2X1_1/A XNOR2X1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M10163 XNOR2X1_1/Y XNOR2X1_1/A XNOR2X1_1/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M10164 XNOR2X1_1/a_12_41# NOR2X1_0/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10165 XNOR2X1_1/a_18_54# XNOR2X1_1/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M10166 XNOR2X1_1/a_35_6# XNOR2X1_1/a_2_6# XNOR2X1_1/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10167 XNOR2X1_1/a_18_6# XNOR2X1_1/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10168 vdd XNOR2X1_1/A XNOR2X1_1/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M10169 vdd NOR2X1_0/Y XNOR2X1_1/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M10170 XNOR2X1_1/Y XNOR2X1_1/a_2_6# XNOR2X1_1/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M10171 XNOR2X1_1/a_35_54# XNOR2X1_1/A XNOR2X1_1/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10172 XNOR2X1_1/a_12_41# NOR2X1_0/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10173 gnd NOR2X1_0/Y XNOR2X1_1/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10174 DFFNEGX1_80/a_76_6# BUFX2_11/Y DFFNEGX1_80/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M10175 gnd BUFX2_11/Y DFFNEGX1_80/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M10176 DFFNEGX1_80/a_66_6# DFFNEGX1_80/a_2_6# DFFNEGX1_80/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10177 out_temp_cleared[11] DFFNEGX1_80/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10178 DFFNEGX1_80/a_23_6# BUFX2_11/Y DFFNEGX1_80/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M10179 DFFNEGX1_80/a_23_6# DFFNEGX1_80/a_2_6# DFFNEGX1_80/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M10180 gnd DFFNEGX1_80/a_34_4# DFFNEGX1_80/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10181 vdd DFFNEGX1_80/a_34_4# DFFNEGX1_80/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M10182 DFFNEGX1_80/a_61_74# DFFNEGX1_80/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10183 DFFNEGX1_80/a_34_4# DFFNEGX1_80/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10184 DFFNEGX1_80/a_34_4# DFFNEGX1_80/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M10185 vdd out_temp_cleared[11] DFFNEGX1_80/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10186 gnd out_temp_cleared[11] DFFNEGX1_80/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10187 DFFNEGX1_80/a_61_6# DFFNEGX1_80/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10188 DFFNEGX1_80/a_76_84# DFFNEGX1_80/a_2_6# DFFNEGX1_80/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M10189 out_temp_cleared[11] DFFNEGX1_80/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10190 vdd BUFX2_11/Y DFFNEGX1_80/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M10191 DFFNEGX1_80/a_31_6# DFFNEGX1_80/a_2_6# DFFNEGX1_80/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10192 DFFNEGX1_80/a_66_6# BUFX2_11/Y DFFNEGX1_80/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10193 DFFNEGX1_80/a_17_74# OAI22X1_17/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10194 DFFNEGX1_80/a_31_74# BUFX2_11/Y DFFNEGX1_80/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10195 DFFNEGX1_80/a_17_6# OAI22X1_17/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10196 DFFNEGX1_91/a_76_6# BUFX2_11/Y DFFNEGX1_91/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M10197 gnd BUFX2_11/Y DFFNEGX1_91/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M10198 DFFNEGX1_91/a_66_6# DFFNEGX1_91/a_2_6# DFFNEGX1_91/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10199 out_temp_cleared[0] DFFNEGX1_91/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10200 DFFNEGX1_91/a_23_6# BUFX2_11/Y DFFNEGX1_91/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M10201 DFFNEGX1_91/a_23_6# DFFNEGX1_91/a_2_6# DFFNEGX1_91/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M10202 gnd DFFNEGX1_91/a_34_4# DFFNEGX1_91/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10203 vdd DFFNEGX1_91/a_34_4# DFFNEGX1_91/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M10204 DFFNEGX1_91/a_61_74# DFFNEGX1_91/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10205 DFFNEGX1_91/a_34_4# DFFNEGX1_91/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10206 DFFNEGX1_91/a_34_4# DFFNEGX1_91/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M10207 vdd out_temp_cleared[0] DFFNEGX1_91/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10208 gnd out_temp_cleared[0] DFFNEGX1_91/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10209 DFFNEGX1_91/a_61_6# DFFNEGX1_91/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10210 DFFNEGX1_91/a_76_84# DFFNEGX1_91/a_2_6# DFFNEGX1_91/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M10211 out_temp_cleared[0] DFFNEGX1_91/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10212 vdd BUFX2_11/Y DFFNEGX1_91/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M10213 DFFNEGX1_91/a_31_6# DFFNEGX1_91/a_2_6# DFFNEGX1_91/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10214 DFFNEGX1_91/a_66_6# BUFX2_11/Y DFFNEGX1_91/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10215 DFFNEGX1_91/a_17_74# OAI22X1_28/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10216 DFFNEGX1_91/a_31_74# BUFX2_11/Y DFFNEGX1_91/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10217 DFFNEGX1_91/a_17_6# OAI22X1_28/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10218 vdd out_global_score[25] HAX1_5/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M10219 HAX1_5/a_41_74# HAX1_5/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M10220 HAX1_5/a_9_6# out_global_score[25] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10221 HAX1_5/a_41_74# HAX1_5/B HAX1_5/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M10222 vdd out_global_score[25] HAX1_5/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M10223 vdd HAX1_5/a_2_74# HAX1_4/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M10224 HAX1_5/a_38_6# HAX1_5/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10225 HAX1_5/YS HAX1_5/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10226 HAX1_5/a_38_6# out_global_score[25] HAX1_5/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10227 HAX1_5/YS HAX1_5/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M10228 HAX1_5/a_2_74# HAX1_5/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10229 HAX1_5/a_2_74# HAX1_5/B HAX1_5/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10230 HAX1_5/a_49_54# HAX1_5/B HAX1_5/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10231 gnd HAX1_5/a_2_74# HAX1_4/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M10232 AND2X2_1/a_2_6# XOR2X1_8/A vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M10233 AND2X2_1/a_9_6# XOR2X1_8/A AND2X2_1/a_2_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=100p ps=50u
M10234 XOR2X1_7/A AND2X2_1/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10235 XOR2X1_7/A AND2X2_1/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10236 vdd FAX1_6/YS AND2X2_1/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10237 gnd FAX1_6/YS AND2X2_1/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10238 NOR2X1_73/A INVX2_71/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M10239 NAND3X1_17/a_9_6# INVX2_71/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M10240 NOR2X1_73/A NOR2X1_74/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10241 NOR2X1_73/A NOR2X1_74/Y NAND3X1_17/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M10242 vdd INVX2_66/Y NOR2X1_73/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10243 NAND3X1_17/a_14_6# INVX2_66/Y NAND3X1_17/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M10244 NOR2X1_91/B NAND3X1_39/A vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M10245 NAND3X1_39/a_9_6# NAND3X1_39/A gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M10246 NOR2X1_91/B AOI21X1_5/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10247 NOR2X1_91/B AOI21X1_5/Y NAND3X1_39/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M10248 vdd NAND3X1_39/B NOR2X1_91/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10249 NAND3X1_39/a_14_6# NAND3X1_39/B NAND3X1_39/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M10250 NOR2X1_82/B NOR2X1_86/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M10251 NAND3X1_28/a_9_6# NOR2X1_86/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M10252 NOR2X1_82/B NOR2X1_83/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10253 NOR2X1_82/B NOR2X1_83/Y NAND3X1_28/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M10254 vdd NOR2X1_85/Y NOR2X1_82/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10255 NAND3X1_28/a_14_6# NOR2X1_85/Y NAND3X1_28/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M10256 FAX1_15/A INVX2_17/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M10257 FAX1_15/A NOR2X1_17/B NOR2X1_17/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M10258 NOR2X1_17/a_9_54# INVX2_17/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10259 gnd NOR2X1_17/B FAX1_15/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10260 HAX1_32/B INVX2_1/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M10261 HAX1_32/B NOR2X1_32/B NOR2X1_28/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M10262 NOR2X1_28/a_9_54# INVX2_1/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10263 gnd NOR2X1_32/B HAX1_32/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10264 NOR2X1_39/Y NOR2X1_55/A gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M10265 NOR2X1_39/Y NOR2X1_40/B NOR2X1_39/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M10266 NOR2X1_39/a_9_54# NOR2X1_55/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10267 gnd NOR2X1_40/B NOR2X1_39/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10268 INVX2_206/Y INVX2_206/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10269 INVX2_206/Y INVX2_206/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10270 INVX2_239/Y INVX2_239/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10271 INVX2_239/Y INVX2_239/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10272 OAI21X1_7/A OAI21X1_8/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10273 OAI21X1_7/A OAI21X1_8/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10274 INVX2_217/Y INVX2_217/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10275 INVX2_217/Y INVX2_217/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10276 gnd XNOR2X1_8/Y MUX2X1_13/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M10277 MUX2X1_13/a_17_50# NOR2X1_4/A vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M10278 XNOR2X1_7/A OR2X1_4/Y MUX2X1_13/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M10279 MUX2X1_13/a_30_54# MUX2X1_13/a_2_10# XNOR2X1_7/A vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M10280 MUX2X1_13/a_17_10# NOR2X1_4/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10281 vdd OR2X1_4/Y MUX2X1_13/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M10282 MUX2X1_13/a_30_10# OR2X1_4/Y XNOR2X1_7/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M10283 gnd OR2X1_4/Y MUX2X1_13/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M10284 vdd XNOR2X1_8/Y MUX2X1_13/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10285 XNOR2X1_7/A MUX2X1_13/a_2_10# MUX2X1_13/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10286 gnd MUX2X1_24/A MUX2X1_24/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M10287 MUX2X1_24/a_17_50# FAX1_2/YS vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M10288 MUX2X1_24/Y OR2X1_2/Y MUX2X1_24/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M10289 MUX2X1_24/a_30_54# MUX2X1_24/a_2_10# MUX2X1_24/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M10290 MUX2X1_24/a_17_10# FAX1_2/YS gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10291 vdd OR2X1_2/Y MUX2X1_24/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M10292 MUX2X1_24/a_30_10# OR2X1_2/Y MUX2X1_24/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M10293 gnd OR2X1_2/Y MUX2X1_24/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M10294 vdd MUX2X1_24/A MUX2X1_24/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10295 MUX2X1_24/Y MUX2X1_24/a_2_10# MUX2X1_24/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10296 NOR2X1_118/Y BUFX2_3/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M10297 NOR2X1_118/Y NOR2X1_118/B NOR2X1_118/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M10298 NOR2X1_118/a_9_54# BUFX2_3/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10299 gnd NOR2X1_118/B NOR2X1_118/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10300 NOR2X1_107/Y INVX2_129/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M10301 NOR2X1_107/Y BUFX2_3/Y NOR2X1_107/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M10302 NOR2X1_107/a_9_54# INVX2_129/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10303 gnd BUFX2_3/Y NOR2X1_107/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10304 OAI21X1_55/C out_temp_index[1] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M10305 NAND2X1_50/a_9_6# out_temp_index[1] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10306 vdd NOR2X1_67/Y OAI21X1_55/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10307 OAI21X1_55/C NOR2X1_67/Y NAND2X1_50/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10308 NOR2X1_71/B OR2X1_14/A vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M10309 NAND2X1_61/a_9_6# OR2X1_14/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10310 vdd INVX2_85/Y NOR2X1_71/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10311 NOR2X1_71/B INVX2_85/Y NAND2X1_61/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10312 OAI21X1_96/C NOR2X1_54/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M10313 NAND2X1_83/a_9_6# NOR2X1_54/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10314 vdd BUFX2_21/Y OAI21X1_96/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10315 OAI21X1_96/C BUFX2_21/Y NAND2X1_83/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10316 OAI21X1_85/C NOR2X1_41/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M10317 NAND2X1_72/a_9_6# NOR2X1_41/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10318 vdd BUFX2_20/Y OAI21X1_85/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10319 OAI21X1_85/C BUFX2_20/Y NAND2X1_72/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10320 BUFX2_23/A INVX2_217/A vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M10321 NAND2X1_94/a_9_6# INVX2_217/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10322 vdd NOR2X1_104/B BUFX2_23/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10323 BUFX2_23/A NOR2X1_104/B NAND2X1_94/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10324 gnd INVX2_31/Y AOI22X1_70/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M10325 AOI22X1_70/Y out_mines[8] AOI22X1_70/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M10326 AOI22X1_70/a_11_6# INVX2_32/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10327 AOI22X1_70/a_2_54# out_mines[8] vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M10328 AOI22X1_70/a_28_6# out_mines[16] AOI22X1_70/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10329 vdd INVX2_32/Y AOI22X1_70/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10330 AOI22X1_70/Y out_mines[16] AOI22X1_70/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M10331 AOI22X1_70/a_2_54# INVX2_31/Y AOI22X1_70/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10332 INVX2_30/Y out_temp_data_in[4] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10333 INVX2_30/Y out_temp_data_in[4] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10334 INVX2_52/Y INVX2_52/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10335 INVX2_52/Y INVX2_52/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10336 INVX2_63/Y out_temp_decoded[18] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10337 INVX2_63/Y out_temp_decoded[18] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10338 INVX2_41/Y INVX2_41/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10339 INVX2_41/Y INVX2_41/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10340 INVX2_74/Y out_temp_decoded[8] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10341 INVX2_74/Y out_temp_decoded[8] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10342 INVX2_96/Y out_temp_cleared[17] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10343 INVX2_96/Y out_temp_cleared[17] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10344 INVX2_85/Y out_temp_decoded[0] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10345 INVX2_85/Y out_temp_decoded[0] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10346 gnd INVX2_240/Y OAI21X1_15/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M10347 vdd OAI21X1_15/C OAI21X1_15/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M10348 OAI21X1_15/Y OAI21X1_15/C OAI21X1_15/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10349 OAI21X1_15/Y OAI21X1_9/B OAI21X1_15/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M10350 OAI21X1_15/a_9_54# INVX2_240/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10351 OAI21X1_15/a_2_6# OAI21X1_9/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10352 gnd OAI21X1_44/A OAI21X1_26/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M10353 vdd BUFX2_19/Y INVX2_235/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M10354 INVX2_235/A BUFX2_19/Y OAI21X1_26/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10355 INVX2_235/A OAI21X1_30/B OAI21X1_26/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M10356 OAI21X1_26/a_9_54# OAI21X1_44/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10357 OAI21X1_26/a_2_6# OAI21X1_30/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10358 gnd NAND3X1_7/Y OAI21X1_48/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M10359 vdd BUFX2_18/Y INVX2_244/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M10360 INVX2_244/A BUFX2_18/Y OAI21X1_48/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10361 INVX2_244/A OAI21X1_48/B OAI21X1_48/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M10362 OAI21X1_48/a_9_54# NAND3X1_7/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10363 OAI21X1_48/a_2_6# OAI21X1_48/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10364 gnd INVX2_231/Y OAI21X1_37/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M10365 vdd OAI21X1_37/C OAI21X1_37/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M10366 OAI21X1_37/Y OAI21X1_37/C OAI21X1_37/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10367 OAI21X1_37/Y OAI21X1_9/B OAI21X1_37/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M10368 OAI21X1_37/a_9_54# INVX2_231/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10369 OAI21X1_37/a_2_6# OAI21X1_9/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10370 gnd OAI21X1_59/A OAI21X1_59/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M10371 vdd OAI21X1_59/C OAI21X1_59/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M10372 OAI21X1_59/Y OAI21X1_59/C OAI21X1_59/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10373 OAI21X1_59/Y OAI21X1_59/B OAI21X1_59/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M10374 OAI21X1_59/a_9_54# OAI21X1_59/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10375 OAI21X1_59/a_2_6# OAI21X1_59/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10376 AND2X2_18/a_2_6# out_state_main[2] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M10377 AND2X2_18/a_9_6# out_state_main[2] AND2X2_18/a_2_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=100p ps=50u
M10378 AND2X2_18/Y AND2X2_18/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10379 AND2X2_18/Y AND2X2_18/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10380 vdd out_state_main[0] AND2X2_18/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10381 gnd out_state_main[0] AND2X2_18/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10382 gnd NOR2X1_1/A XNOR2X1_2/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M10383 XNOR2X1_2/Y NOR2X1_1/A XNOR2X1_2/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M10384 XNOR2X1_2/a_12_41# FAX1_3/YS gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10385 XNOR2X1_2/a_18_54# XNOR2X1_2/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M10386 XNOR2X1_2/a_35_6# XNOR2X1_2/a_2_6# XNOR2X1_2/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10387 XNOR2X1_2/a_18_6# XNOR2X1_2/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10388 vdd NOR2X1_1/A XNOR2X1_2/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M10389 vdd FAX1_3/YS XNOR2X1_2/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M10390 XNOR2X1_2/Y XNOR2X1_2/a_2_6# XNOR2X1_2/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M10391 XNOR2X1_2/a_35_54# NOR2X1_1/A XNOR2X1_2/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10392 XNOR2X1_2/a_12_41# FAX1_3/YS vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10393 gnd FAX1_3/YS XNOR2X1_2/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10394 DFFNEGX1_70/a_76_6# BUFX2_12/Y DFFNEGX1_70/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M10395 gnd BUFX2_12/Y DFFNEGX1_70/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M10396 DFFNEGX1_70/a_66_6# DFFNEGX1_70/a_2_6# DFFNEGX1_70/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10397 out_temp_cleared[21] DFFNEGX1_70/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10398 DFFNEGX1_70/a_23_6# BUFX2_12/Y DFFNEGX1_70/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M10399 DFFNEGX1_70/a_23_6# DFFNEGX1_70/a_2_6# DFFNEGX1_70/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M10400 gnd DFFNEGX1_70/a_34_4# DFFNEGX1_70/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10401 vdd DFFNEGX1_70/a_34_4# DFFNEGX1_70/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M10402 DFFNEGX1_70/a_61_74# DFFNEGX1_70/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10403 DFFNEGX1_70/a_34_4# DFFNEGX1_70/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10404 DFFNEGX1_70/a_34_4# DFFNEGX1_70/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M10405 vdd out_temp_cleared[21] DFFNEGX1_70/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10406 gnd out_temp_cleared[21] DFFNEGX1_70/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10407 DFFNEGX1_70/a_61_6# DFFNEGX1_70/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10408 DFFNEGX1_70/a_76_84# DFFNEGX1_70/a_2_6# DFFNEGX1_70/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M10409 out_temp_cleared[21] DFFNEGX1_70/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10410 vdd BUFX2_12/Y DFFNEGX1_70/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M10411 DFFNEGX1_70/a_31_6# DFFNEGX1_70/a_2_6# DFFNEGX1_70/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10412 DFFNEGX1_70/a_66_6# BUFX2_12/Y DFFNEGX1_70/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10413 DFFNEGX1_70/a_17_74# OAI22X1_7/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10414 DFFNEGX1_70/a_31_74# BUFX2_12/Y DFFNEGX1_70/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10415 DFFNEGX1_70/a_17_6# OAI22X1_7/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10416 DFFNEGX1_81/a_76_6# BUFX2_11/Y DFFNEGX1_81/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M10417 gnd BUFX2_11/Y DFFNEGX1_81/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M10418 DFFNEGX1_81/a_66_6# DFFNEGX1_81/a_2_6# DFFNEGX1_81/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10419 out_temp_cleared[10] DFFNEGX1_81/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10420 DFFNEGX1_81/a_23_6# BUFX2_11/Y DFFNEGX1_81/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M10421 DFFNEGX1_81/a_23_6# DFFNEGX1_81/a_2_6# DFFNEGX1_81/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M10422 gnd DFFNEGX1_81/a_34_4# DFFNEGX1_81/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10423 vdd DFFNEGX1_81/a_34_4# DFFNEGX1_81/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M10424 DFFNEGX1_81/a_61_74# DFFNEGX1_81/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10425 DFFNEGX1_81/a_34_4# DFFNEGX1_81/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10426 DFFNEGX1_81/a_34_4# DFFNEGX1_81/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M10427 vdd out_temp_cleared[10] DFFNEGX1_81/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10428 gnd out_temp_cleared[10] DFFNEGX1_81/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10429 DFFNEGX1_81/a_61_6# DFFNEGX1_81/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10430 DFFNEGX1_81/a_76_84# DFFNEGX1_81/a_2_6# DFFNEGX1_81/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M10431 out_temp_cleared[10] DFFNEGX1_81/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10432 vdd BUFX2_11/Y DFFNEGX1_81/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M10433 DFFNEGX1_81/a_31_6# DFFNEGX1_81/a_2_6# DFFNEGX1_81/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10434 DFFNEGX1_81/a_66_6# BUFX2_11/Y DFFNEGX1_81/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10435 DFFNEGX1_81/a_17_74# OAI22X1_18/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10436 DFFNEGX1_81/a_31_74# BUFX2_11/Y DFFNEGX1_81/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10437 DFFNEGX1_81/a_17_6# OAI22X1_18/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10438 DFFNEGX1_92/a_76_6# BUFX2_11/Y DFFNEGX1_92/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M10439 gnd BUFX2_11/Y DFFNEGX1_92/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M10440 DFFNEGX1_92/a_66_6# DFFNEGX1_92/a_2_6# DFFNEGX1_92/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10441 out_gameover DFFNEGX1_92/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10442 DFFNEGX1_92/a_23_6# BUFX2_11/Y DFFNEGX1_92/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M10443 DFFNEGX1_92/a_23_6# DFFNEGX1_92/a_2_6# DFFNEGX1_92/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M10444 gnd DFFNEGX1_92/a_34_4# DFFNEGX1_92/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10445 vdd DFFNEGX1_92/a_34_4# DFFNEGX1_92/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M10446 DFFNEGX1_92/a_61_74# DFFNEGX1_92/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10447 DFFNEGX1_92/a_34_4# DFFNEGX1_92/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10448 DFFNEGX1_92/a_34_4# DFFNEGX1_92/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M10449 vdd out_gameover DFFNEGX1_92/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10450 gnd out_gameover DFFNEGX1_92/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10451 DFFNEGX1_92/a_61_6# DFFNEGX1_92/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10452 DFFNEGX1_92/a_76_84# DFFNEGX1_92/a_2_6# DFFNEGX1_92/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M10453 out_gameover DFFNEGX1_92/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10454 vdd BUFX2_11/Y DFFNEGX1_92/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M10455 DFFNEGX1_92/a_31_6# DFFNEGX1_92/a_2_6# DFFNEGX1_92/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10456 DFFNEGX1_92/a_66_6# BUFX2_11/Y DFFNEGX1_92/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10457 DFFNEGX1_92/a_17_74# INVX2_218/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10458 DFFNEGX1_92/a_31_74# BUFX2_11/Y DFFNEGX1_92/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10459 DFFNEGX1_92/a_17_6# INVX2_218/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10460 vdd out_global_score[24] HAX1_6/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M10461 HAX1_6/a_41_74# HAX1_6/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M10462 HAX1_6/a_9_6# out_global_score[24] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10463 HAX1_6/a_41_74# HAX1_6/B HAX1_6/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M10464 vdd out_global_score[24] HAX1_6/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M10465 vdd HAX1_6/a_2_74# HAX1_5/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M10466 HAX1_6/a_38_6# HAX1_6/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10467 HAX1_6/YS HAX1_6/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10468 HAX1_6/a_38_6# out_global_score[24] HAX1_6/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10469 HAX1_6/YS HAX1_6/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M10470 HAX1_6/a_2_74# HAX1_6/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10471 HAX1_6/a_2_74# HAX1_6/B HAX1_6/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10472 HAX1_6/a_49_54# HAX1_6/B HAX1_6/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10473 gnd HAX1_6/a_2_74# HAX1_5/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M10474 AND2X2_2/a_2_6# FAX1_0/YC vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M10475 AND2X2_2/a_9_6# FAX1_0/YC AND2X2_2/a_2_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=100p ps=50u
M10476 XOR2X1_8/A AND2X2_2/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10477 XOR2X1_8/A AND2X2_2/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10478 vdd FAX1_7/YS AND2X2_2/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10479 gnd FAX1_7/YS AND2X2_2/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10480 NOR2X1_83/B INVX2_73/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M10481 NAND3X1_29/a_9_6# INVX2_73/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M10482 NOR2X1_83/B INVX2_58/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10483 NOR2X1_83/B INVX2_58/Y NAND3X1_29/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M10484 vdd INVX2_76/Y NOR2X1_83/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10485 NAND3X1_29/a_14_6# INVX2_76/Y NAND3X1_29/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M10486 OR2X1_14/A AND2X2_15/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M10487 NAND3X1_18/a_9_6# AND2X2_15/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M10488 OR2X1_14/A NOR2X1_75/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10489 OR2X1_14/A NOR2X1_75/Y NAND3X1_18/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M10490 vdd INVX2_84/Y OR2X1_14/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10491 NAND3X1_18/a_14_6# INVX2_84/Y NAND3X1_18/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M10492 FAX1_10/A INVX2_1/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M10493 FAX1_10/A NOR2X1_22/B NOR2X1_18/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M10494 NOR2X1_18/a_9_54# INVX2_1/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10495 gnd NOR2X1_22/B FAX1_10/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10496 HAX1_31/B INVX2_2/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M10497 HAX1_31/B NOR2X1_32/B NOR2X1_29/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M10498 NOR2X1_29/a_9_54# INVX2_2/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10499 gnd NOR2X1_32/B HAX1_31/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10500 INVX2_207/Y INVX2_207/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10501 INVX2_207/Y INVX2_207/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10502 INVX2_229/Y INVX2_229/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10503 INVX2_229/Y INVX2_229/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10504 INVX2_218/Y INVX2_218/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10505 INVX2_218/Y INVX2_218/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10506 gnd HAX1_47/YS MUX2X1_25/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M10507 MUX2X1_25/a_17_50# HAX1_47/A vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M10508 MUX2X1_25/Y OR2X1_1/Y MUX2X1_25/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M10509 MUX2X1_25/a_30_54# MUX2X1_25/a_2_10# MUX2X1_25/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M10510 MUX2X1_25/a_17_10# HAX1_47/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10511 vdd OR2X1_1/Y MUX2X1_25/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M10512 MUX2X1_25/a_30_10# OR2X1_1/Y MUX2X1_25/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M10513 gnd OR2X1_1/Y MUX2X1_25/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M10514 vdd HAX1_47/YS MUX2X1_25/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10515 MUX2X1_25/Y MUX2X1_25/a_2_10# MUX2X1_25/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10516 gnd MUX2X1_14/A MUX2X1_14/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M10517 MUX2X1_14/a_17_50# FAX1_0/YS vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M10518 MUX2X1_14/Y OR2X1_4/Y MUX2X1_14/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M10519 MUX2X1_14/a_30_54# MUX2X1_14/a_2_10# MUX2X1_14/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M10520 MUX2X1_14/a_17_10# FAX1_0/YS gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10521 vdd OR2X1_4/Y MUX2X1_14/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M10522 MUX2X1_14/a_30_10# OR2X1_4/Y MUX2X1_14/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M10523 gnd OR2X1_4/Y MUX2X1_14/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M10524 vdd MUX2X1_14/A MUX2X1_14/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10525 MUX2X1_14/Y MUX2X1_14/a_2_10# MUX2X1_14/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10526 NOR2X1_119/Y BUFX2_3/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M10527 NOR2X1_119/Y NOR2X1_119/B NOR2X1_119/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M10528 NOR2X1_119/a_9_54# BUFX2_3/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10529 gnd NOR2X1_119/B NOR2X1_119/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10530 NOR2X1_108/Y INVX2_21/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M10531 NOR2X1_108/Y NOR2X1_110/B NOR2X1_108/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M10532 NOR2X1_108/a_9_54# INVX2_21/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10533 gnd NOR2X1_110/B NOR2X1_108/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10534 OAI21X1_56/C out_temp_index[0] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M10535 NAND2X1_51/a_9_6# out_temp_index[0] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10536 vdd NOR2X1_67/Y OAI21X1_56/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10537 OAI21X1_56/C NOR2X1_67/Y NAND2X1_51/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10538 OAI21X1_43/C out_mines[4] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M10539 NAND2X1_40/a_9_6# out_mines[4] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10540 vdd INVX2_238/Y OAI21X1_43/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10541 OAI21X1_43/C INVX2_238/Y NAND2X1_40/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10542 OAI21X1_97/C NOR2X1_53/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M10543 NAND2X1_84/a_9_6# NOR2X1_53/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10544 vdd BUFX2_21/Y OAI21X1_97/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10545 OAI21X1_97/C BUFX2_21/Y NAND2X1_84/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10546 OAI21X1_86/C NOR2X1_40/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M10547 NAND2X1_73/a_9_6# NOR2X1_40/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10548 vdd BUFX2_20/Y OAI21X1_86/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10549 OAI21X1_86/C BUFX2_20/Y NAND2X1_73/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10550 NOR2X1_104/B out_decode vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M10551 NAND2X1_95/a_9_6# out_decode gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10552 vdd AND2X2_14/B NOR2X1_104/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10553 NOR2X1_104/B AND2X2_14/B NAND2X1_95/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10554 OAI21X1_65/C out_win vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M10555 NAND2X1_62/a_9_6# out_win gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10556 vdd AOI21X1_2/A OAI21X1_65/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10557 OAI21X1_65/C AOI21X1_2/A NAND2X1_62/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10558 gnd out_mines[3] AOI22X1_60/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M10559 AOI22X1_60/Y NOR2X1_113/Y AOI22X1_60/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M10560 AOI22X1_60/a_11_6# out_mines[4] gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10561 AOI22X1_60/a_2_54# NOR2X1_113/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M10562 AOI22X1_60/a_28_6# NOR2X1_114/Y AOI22X1_60/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10563 vdd out_mines[4] AOI22X1_60/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10564 AOI22X1_60/Y NOR2X1_114/Y AOI22X1_60/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M10565 AOI22X1_60/a_2_54# out_mines[3] AOI22X1_60/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10566 gnd INVX2_31/Y AOI22X1_71/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M10567 AOI22X1_71/Y out_mines[7] AOI22X1_71/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M10568 AOI22X1_71/a_11_6# INVX2_32/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10569 AOI22X1_71/a_2_54# out_mines[7] vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M10570 AOI22X1_71/a_28_6# out_mines[15] AOI22X1_71/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10571 vdd INVX2_32/Y AOI22X1_71/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10572 AOI22X1_71/Y out_mines[15] AOI22X1_71/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M10573 AOI22X1_71/a_2_54# INVX2_31/Y AOI22X1_71/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10574 gnd INVX2_85/Y OAI22X1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M10575 OAI22X1_0/a_2_6# INVX2_83/Y OAI22X1_0/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M10576 OAI22X1_0/Y INVX2_10/Y OAI22X1_0/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10577 OAI22X1_0/Y INVX2_9/Y OAI22X1_0/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M10578 OAI22X1_0/a_28_54# INVX2_10/Y OAI22X1_0/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M10579 OAI22X1_0/a_9_54# INVX2_85/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10580 OAI22X1_0/a_2_6# INVX2_9/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10581 vdd INVX2_83/Y OAI22X1_0/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10582 INVX2_20/Y out_mines[22] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10583 INVX2_20/Y out_mines[22] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10584 INVX2_31/Y INVX2_31/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10585 INVX2_31/Y INVX2_31/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10586 INVX2_42/Y INVX2_42/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10587 INVX2_42/Y INVX2_42/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10588 INVX2_53/Y INVX2_53/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10589 INVX2_53/Y INVX2_53/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10590 INVX2_75/Y out_temp_decoded[7] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10591 INVX2_75/Y out_temp_decoded[7] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10592 INVX2_97/Y out_temp_cleared[16] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10593 INVX2_97/Y out_temp_cleared[16] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10594 INVX2_64/Y out_temp_decoded[17] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10595 INVX2_64/Y out_temp_decoded[17] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10596 INVX2_86/Y INVX2_86/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10597 INVX2_86/Y INVX2_86/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10598 gnd OAI21X1_8/B OAI21X1_16/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M10599 vdd BUFX2_19/Y INVX2_240/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M10600 INVX2_240/A BUFX2_19/Y OAI21X1_16/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10601 INVX2_240/A NAND3X1_7/Y OAI21X1_16/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M10602 OAI21X1_16/a_9_54# OAI21X1_8/B vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10603 OAI21X1_16/a_2_6# NAND3X1_7/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10604 gnd INVX2_222/Y OAI21X1_49/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M10605 vdd OAI21X1_49/C OAI21X1_49/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M10606 OAI21X1_49/Y OAI21X1_49/C OAI21X1_49/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10607 OAI21X1_49/Y OAI21X1_9/B OAI21X1_49/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M10608 OAI21X1_49/a_9_54# INVX2_222/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10609 OAI21X1_49/a_2_6# OAI21X1_9/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10610 gnd OAI21X1_8/A OAI21X1_38/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M10611 vdd BUFX2_18/Y INVX2_231/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M10612 INVX2_231/A BUFX2_18/Y OAI21X1_38/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10613 INVX2_231/A OAI21X1_46/B OAI21X1_38/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M10614 OAI21X1_38/a_9_54# OAI21X1_8/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10615 OAI21X1_38/a_2_6# OAI21X1_46/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10616 gnd INVX2_236/Y OAI21X1_27/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M10617 vdd OAI21X1_27/C OAI21X1_27/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M10618 OAI21X1_27/Y OAI21X1_27/C OAI21X1_27/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10619 OAI21X1_27/Y NOR2X1_66/B OAI21X1_27/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M10620 OAI21X1_27/a_9_54# INVX2_236/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10621 OAI21X1_27/a_2_6# NOR2X1_66/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10622 AND2X2_19/a_2_6# INVX2_124/A vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M10623 AND2X2_19/a_9_6# INVX2_124/A AND2X2_19/a_2_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=100p ps=50u
M10624 AND2X2_19/Y AND2X2_19/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10625 AND2X2_19/Y AND2X2_19/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10626 vdd AND2X2_19/B AND2X2_19/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10627 gnd AND2X2_19/B AND2X2_19/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10628 gnd XNOR2X1_3/A XNOR2X1_3/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M10629 XNOR2X1_3/Y XNOR2X1_3/A XNOR2X1_3/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M10630 XNOR2X1_3/a_12_41# NOR2X1_1/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10631 XNOR2X1_3/a_18_54# XNOR2X1_3/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M10632 XNOR2X1_3/a_35_6# XNOR2X1_3/a_2_6# XNOR2X1_3/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10633 XNOR2X1_3/a_18_6# XNOR2X1_3/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10634 vdd XNOR2X1_3/A XNOR2X1_3/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M10635 vdd NOR2X1_1/Y XNOR2X1_3/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M10636 XNOR2X1_3/Y XNOR2X1_3/a_2_6# XNOR2X1_3/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M10637 XNOR2X1_3/a_35_54# XNOR2X1_3/A XNOR2X1_3/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10638 XNOR2X1_3/a_12_41# NOR2X1_1/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10639 gnd NOR2X1_1/Y XNOR2X1_3/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10640 DFFNEGX1_60/a_76_6# BUFX2_13/Y DFFNEGX1_60/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M10641 gnd BUFX2_13/Y DFFNEGX1_60/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M10642 DFFNEGX1_60/a_66_6# DFFNEGX1_60/a_2_6# DFFNEGX1_60/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10643 out_temp_decoded[6] DFFNEGX1_60/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10644 DFFNEGX1_60/a_23_6# BUFX2_13/Y DFFNEGX1_60/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M10645 DFFNEGX1_60/a_23_6# DFFNEGX1_60/a_2_6# DFFNEGX1_60/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M10646 gnd DFFNEGX1_60/a_34_4# DFFNEGX1_60/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10647 vdd DFFNEGX1_60/a_34_4# DFFNEGX1_60/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M10648 DFFNEGX1_60/a_61_74# DFFNEGX1_60/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10649 DFFNEGX1_60/a_34_4# DFFNEGX1_60/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10650 DFFNEGX1_60/a_34_4# DFFNEGX1_60/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M10651 vdd out_temp_decoded[6] DFFNEGX1_60/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10652 gnd out_temp_decoded[6] DFFNEGX1_60/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10653 DFFNEGX1_60/a_61_6# DFFNEGX1_60/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10654 DFFNEGX1_60/a_76_84# DFFNEGX1_60/a_2_6# DFFNEGX1_60/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M10655 out_temp_decoded[6] DFFNEGX1_60/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10656 vdd BUFX2_13/Y DFFNEGX1_60/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M10657 DFFNEGX1_60/a_31_6# DFFNEGX1_60/a_2_6# DFFNEGX1_60/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10658 DFFNEGX1_60/a_66_6# BUFX2_13/Y DFFNEGX1_60/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10659 DFFNEGX1_60/a_17_74# OAI21X1_88/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10660 DFFNEGX1_60/a_31_74# BUFX2_13/Y DFFNEGX1_60/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10661 DFFNEGX1_60/a_17_6# OAI21X1_88/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10662 DFFNEGX1_93/a_76_6# BUFX2_10/Y DFFNEGX1_93/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M10663 gnd BUFX2_10/Y DFFNEGX1_93/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M10664 DFFNEGX1_93/a_66_6# DFFNEGX1_93/a_2_6# DFFNEGX1_93/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10665 out_win DFFNEGX1_93/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10666 DFFNEGX1_93/a_23_6# BUFX2_10/Y DFFNEGX1_93/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M10667 DFFNEGX1_93/a_23_6# DFFNEGX1_93/a_2_6# DFFNEGX1_93/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M10668 gnd DFFNEGX1_93/a_34_4# DFFNEGX1_93/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10669 vdd DFFNEGX1_93/a_34_4# DFFNEGX1_93/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M10670 DFFNEGX1_93/a_61_74# DFFNEGX1_93/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10671 DFFNEGX1_93/a_34_4# DFFNEGX1_93/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10672 DFFNEGX1_93/a_34_4# DFFNEGX1_93/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M10673 vdd out_win DFFNEGX1_93/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10674 gnd out_win DFFNEGX1_93/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10675 DFFNEGX1_93/a_61_6# DFFNEGX1_93/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10676 DFFNEGX1_93/a_76_84# DFFNEGX1_93/a_2_6# DFFNEGX1_93/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M10677 out_win DFFNEGX1_93/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10678 vdd BUFX2_10/Y DFFNEGX1_93/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M10679 DFFNEGX1_93/a_31_6# DFFNEGX1_93/a_2_6# DFFNEGX1_93/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10680 DFFNEGX1_93/a_66_6# BUFX2_10/Y DFFNEGX1_93/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10681 DFFNEGX1_93/a_17_74# OAI21X1_65/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10682 DFFNEGX1_93/a_31_74# BUFX2_10/Y DFFNEGX1_93/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10683 DFFNEGX1_93/a_17_6# OAI21X1_65/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10684 DFFNEGX1_82/a_76_6# BUFX2_11/Y DFFNEGX1_82/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M10685 gnd BUFX2_11/Y DFFNEGX1_82/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M10686 DFFNEGX1_82/a_66_6# DFFNEGX1_82/a_2_6# DFFNEGX1_82/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10687 out_temp_cleared[9] DFFNEGX1_82/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10688 DFFNEGX1_82/a_23_6# BUFX2_11/Y DFFNEGX1_82/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M10689 DFFNEGX1_82/a_23_6# DFFNEGX1_82/a_2_6# DFFNEGX1_82/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M10690 gnd DFFNEGX1_82/a_34_4# DFFNEGX1_82/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10691 vdd DFFNEGX1_82/a_34_4# DFFNEGX1_82/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M10692 DFFNEGX1_82/a_61_74# DFFNEGX1_82/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10693 DFFNEGX1_82/a_34_4# DFFNEGX1_82/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10694 DFFNEGX1_82/a_34_4# DFFNEGX1_82/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M10695 vdd out_temp_cleared[9] DFFNEGX1_82/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10696 gnd out_temp_cleared[9] DFFNEGX1_82/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10697 DFFNEGX1_82/a_61_6# DFFNEGX1_82/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10698 DFFNEGX1_82/a_76_84# DFFNEGX1_82/a_2_6# DFFNEGX1_82/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M10699 out_temp_cleared[9] DFFNEGX1_82/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10700 vdd BUFX2_11/Y DFFNEGX1_82/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M10701 DFFNEGX1_82/a_31_6# DFFNEGX1_82/a_2_6# DFFNEGX1_82/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10702 DFFNEGX1_82/a_66_6# BUFX2_11/Y DFFNEGX1_82/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10703 DFFNEGX1_82/a_17_74# OAI22X1_19/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10704 DFFNEGX1_82/a_31_74# BUFX2_11/Y DFFNEGX1_82/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10705 DFFNEGX1_82/a_17_6# OAI22X1_19/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10706 DFFNEGX1_71/a_76_6# BUFX2_12/Y DFFNEGX1_71/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M10707 gnd BUFX2_12/Y DFFNEGX1_71/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M10708 DFFNEGX1_71/a_66_6# DFFNEGX1_71/a_2_6# DFFNEGX1_71/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10709 out_temp_cleared[20] DFFNEGX1_71/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10710 DFFNEGX1_71/a_23_6# BUFX2_12/Y DFFNEGX1_71/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M10711 DFFNEGX1_71/a_23_6# DFFNEGX1_71/a_2_6# DFFNEGX1_71/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M10712 gnd DFFNEGX1_71/a_34_4# DFFNEGX1_71/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10713 vdd DFFNEGX1_71/a_34_4# DFFNEGX1_71/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M10714 DFFNEGX1_71/a_61_74# DFFNEGX1_71/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10715 DFFNEGX1_71/a_34_4# DFFNEGX1_71/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10716 DFFNEGX1_71/a_34_4# DFFNEGX1_71/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M10717 vdd out_temp_cleared[20] DFFNEGX1_71/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10718 gnd out_temp_cleared[20] DFFNEGX1_71/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10719 DFFNEGX1_71/a_61_6# DFFNEGX1_71/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10720 DFFNEGX1_71/a_76_84# DFFNEGX1_71/a_2_6# DFFNEGX1_71/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M10721 out_temp_cleared[20] DFFNEGX1_71/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10722 vdd BUFX2_12/Y DFFNEGX1_71/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M10723 DFFNEGX1_71/a_31_6# DFFNEGX1_71/a_2_6# DFFNEGX1_71/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10724 DFFNEGX1_71/a_66_6# BUFX2_12/Y DFFNEGX1_71/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10725 DFFNEGX1_71/a_17_74# OAI22X1_8/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10726 DFFNEGX1_71/a_31_74# BUFX2_12/Y DFFNEGX1_71/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10727 DFFNEGX1_71/a_17_6# OAI22X1_8/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10728 vdd out_global_score[23] HAX1_7/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M10729 HAX1_7/a_41_74# HAX1_7/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M10730 HAX1_7/a_9_6# out_global_score[23] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10731 HAX1_7/a_41_74# HAX1_7/B HAX1_7/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M10732 vdd out_global_score[23] HAX1_7/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M10733 vdd HAX1_7/a_2_74# HAX1_6/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M10734 HAX1_7/a_38_6# HAX1_7/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10735 HAX1_7/YS HAX1_7/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10736 HAX1_7/a_38_6# out_global_score[23] HAX1_7/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10737 HAX1_7/YS HAX1_7/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M10738 HAX1_7/a_2_74# HAX1_7/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10739 HAX1_7/a_2_74# HAX1_7/B HAX1_7/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10740 HAX1_7/a_49_54# HAX1_7/B HAX1_7/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10741 gnd HAX1_7/a_2_74# HAX1_6/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M10742 AND2X2_3/a_2_6# in_incr[0] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M10743 AND2X2_3/a_9_6# in_incr[0] AND2X2_3/a_2_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=100p ps=50u
M10744 FAX1_3/C AND2X2_3/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10745 FAX1_3/C AND2X2_3/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10746 vdd NOR2X1_8/Y AND2X2_3/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10747 gnd NOR2X1_8/Y AND2X2_3/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10748 NOR2X1_75/B INVX2_67/Y vdd vdd pfet w=20 l=2
+  ad=0.22n pd=0.102m as=0 ps=0
M10749 NAND3X1_19/a_9_6# INVX2_67/Y gnd Gnd nfet w=30 l=2
+  ad=90p pd=66u as=0 ps=0
M10750 NOR2X1_75/B NOR2X1_76/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10751 NOR2X1_75/B NOR2X1_76/Y NAND3X1_19/a_14_6# Gnd nfet w=30 l=2
+  ad=0.15n pd=70u as=90p ps=66u
M10752 vdd INVX2_61/Y NOR2X1_75/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10753 NAND3X1_19/a_14_6# INVX2_61/Y NAND3X1_19/a_9_6# Gnd nfet w=30 l=2
+  ad=0 pd=0 as=0 ps=0
M10754 HAX1_33/A INVX2_2/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M10755 HAX1_33/A NOR2X1_22/B NOR2X1_19/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M10756 NOR2X1_19/a_9_54# INVX2_2/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10757 gnd NOR2X1_22/B HAX1_33/A Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10758 INVX2_208/Y INVX2_208/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10759 INVX2_208/Y INVX2_208/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10760 AND2X2_8/A BUFX2_3/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10761 AND2X2_8/A BUFX2_3/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10762 gnd HAX1_43/YS MUX2X1_15/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M10763 MUX2X1_15/a_17_50# HAX1_43/A vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M10764 MUX2X1_15/Y OR2X1_3/Y MUX2X1_15/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M10765 MUX2X1_15/a_30_54# MUX2X1_15/a_2_10# MUX2X1_15/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M10766 MUX2X1_15/a_17_10# HAX1_43/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10767 vdd OR2X1_3/Y MUX2X1_15/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M10768 MUX2X1_15/a_30_10# OR2X1_3/Y MUX2X1_15/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M10769 gnd OR2X1_3/Y MUX2X1_15/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M10770 vdd HAX1_43/YS MUX2X1_15/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10771 MUX2X1_15/Y MUX2X1_15/a_2_10# MUX2X1_15/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10772 gnd HAX1_46/YS MUX2X1_26/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M10773 MUX2X1_26/a_17_50# HAX1_46/A vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M10774 MUX2X1_26/Y OR2X1_1/Y MUX2X1_26/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M10775 MUX2X1_26/a_30_54# MUX2X1_26/a_2_10# MUX2X1_26/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M10776 MUX2X1_26/a_17_10# HAX1_46/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10777 vdd OR2X1_1/Y MUX2X1_26/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M10778 MUX2X1_26/a_30_10# OR2X1_1/Y MUX2X1_26/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M10779 gnd OR2X1_1/Y MUX2X1_26/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M10780 vdd HAX1_46/YS MUX2X1_26/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10781 MUX2X1_26/Y MUX2X1_26/a_2_10# MUX2X1_26/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10782 NOR2X1_109/Y INVX2_24/Y gnd Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=0 ps=0
M10783 NOR2X1_109/Y OAI22X1_38/C NOR2X1_109/a_9_54# vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0.12n ps=86u
M10784 NOR2X1_109/a_9_54# INVX2_24/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10785 gnd OAI22X1_38/C NOR2X1_109/Y Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10786 OAI21X1_44/A NOR2X1_66/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M10787 NAND2X1_41/a_9_6# NOR2X1_66/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10788 vdd NAND3X1_9/A OAI21X1_44/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10789 OAI21X1_44/A NAND3X1_9/A NAND2X1_41/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10790 OAI21X1_29/C out_mines[11] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M10791 NAND2X1_30/a_9_6# out_mines[11] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10792 vdd INVX2_241/Y OAI21X1_29/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10793 OAI21X1_29/C INVX2_241/Y NAND2X1_30/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10794 AND2X2_8/B out_start vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M10795 NAND2X1_52/a_9_6# out_start gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10796 vdd AND2X2_8/A AND2X2_8/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10797 AND2X2_8/B AND2X2_8/A NAND2X1_52/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10798 OAI21X1_98/C NOR2X1_52/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M10799 NAND2X1_85/a_9_6# NOR2X1_52/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10800 vdd BUFX2_21/Y OAI21X1_98/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10801 OAI21X1_98/C BUFX2_21/Y NAND2X1_85/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10802 OAI21X1_87/C NOR2X1_39/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M10803 NAND2X1_74/a_9_6# NOR2X1_39/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10804 vdd BUFX2_20/Y OAI21X1_87/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10805 OAI21X1_87/C BUFX2_20/Y NAND2X1_74/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10806 INVX2_58/A NAND2X1_63/A vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M10807 NAND2X1_63/a_9_6# NAND2X1_63/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10808 vdd NAND2X1_63/B INVX2_58/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10809 INVX2_58/A NAND2X1_63/B NAND2X1_63/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10810 NAND2X1_96/Y in_data[0] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M10811 NAND2X1_96/a_9_6# in_data[0] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10812 vdd NOR2X1_107/Y NAND2X1_96/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10813 NAND2X1_96/Y NOR2X1_107/Y NAND2X1_96/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10814 gnd out_temp_cleared[21] AOI22X1_50/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M10815 NAND3X1_46/B INVX2_23/Y AOI22X1_50/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M10816 AOI22X1_50/a_11_6# NOR2X1_101/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10817 AOI22X1_50/a_2_54# INVX2_23/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M10818 AOI22X1_50/a_28_6# out_mines[21] NAND3X1_46/B Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10819 vdd NOR2X1_101/Y AOI22X1_50/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10820 NAND3X1_46/B out_mines[21] AOI22X1_50/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M10821 AOI22X1_50/a_2_54# out_temp_cleared[21] NAND3X1_46/B vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10822 gnd INVX2_51/A AOI22X1_72/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M10823 AOI22X1_72/Y INVX2_51/Y AOI22X1_72/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M10824 AOI22X1_72/a_11_6# AOI22X1_72/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10825 AOI22X1_72/a_2_54# INVX2_51/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M10826 AOI22X1_72/a_28_6# INVX2_23/Y AOI22X1_72/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10827 vdd AOI22X1_72/A AOI22X1_72/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10828 AOI22X1_72/Y INVX2_23/Y AOI22X1_72/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M10829 AOI22X1_72/a_2_54# INVX2_51/A AOI22X1_72/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10830 gnd out_mines[1] AOI22X1_61/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M10831 AOI22X1_61/Y NOR2X1_111/Y AOI22X1_61/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M10832 AOI22X1_61/a_11_6# out_mines[2] gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10833 AOI22X1_61/a_2_54# NOR2X1_111/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M10834 AOI22X1_61/a_28_6# NOR2X1_112/Y AOI22X1_61/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10835 vdd out_mines[2] AOI22X1_61/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10836 AOI22X1_61/Y NOR2X1_112/Y AOI22X1_61/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M10837 AOI22X1_61/a_2_54# out_mines[1] AOI22X1_61/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10838 gnd INVX2_15/Y OAI22X1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M10839 OAI22X1_1/a_2_6# INVX2_5/Y OAI22X1_1/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M10840 OAI22X1_1/Y OAI22X1_1/D OAI22X1_1/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10841 OAI22X1_1/Y OAI22X1_1/B OAI22X1_1/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M10842 OAI22X1_1/a_28_54# OAI22X1_1/D OAI22X1_1/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M10843 OAI22X1_1/a_9_54# INVX2_15/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10844 OAI22X1_1/a_2_6# OAI22X1_1/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10845 vdd INVX2_5/Y OAI22X1_1/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10846 INVX2_21/Y out_mines[20] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10847 INVX2_21/Y out_mines[20] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10848 INVX2_10/Y out_mines[1] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10849 INVX2_10/Y out_mines[1] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10850 INVX2_54/Y INVX2_54/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10851 INVX2_54/Y INVX2_54/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10852 INVX2_43/Y INVX2_43/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10853 INVX2_43/Y INVX2_43/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10854 INVX2_32/Y INVX2_32/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10855 INVX2_32/Y INVX2_32/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10856 INVX2_65/Y out_temp_decoded[16] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10857 INVX2_65/Y out_temp_decoded[16] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10858 INVX2_76/Y INVX2_76/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10859 INVX2_76/Y INVX2_76/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10860 OR2X1_14/B INVX2_87/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10861 OR2X1_14/B INVX2_87/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10862 INVX2_98/Y out_temp_cleared[15] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10863 INVX2_98/Y out_temp_cleared[15] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10864 gnd INVX2_220/Y OAI21X1_17/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M10865 vdd OAI21X1_17/C OAI21X1_17/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M10866 OAI21X1_17/Y OAI21X1_17/C OAI21X1_17/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10867 OAI21X1_17/Y OAI21X1_9/B OAI21X1_17/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M10868 OAI21X1_17/a_9_54# INVX2_220/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10869 OAI21X1_17/a_2_6# OAI21X1_9/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10870 gnd OAI21X1_44/A OAI21X1_28/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M10871 vdd BUFX2_18/Y INVX2_236/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M10872 INVX2_236/A BUFX2_18/Y OAI21X1_28/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10873 INVX2_236/A OAI21X1_32/B OAI21X1_28/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M10874 OAI21X1_28/a_9_54# OAI21X1_44/A vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10875 OAI21X1_28/a_2_6# OAI21X1_32/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10876 gnd INVX2_232/Y OAI21X1_39/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M10877 vdd OAI21X1_39/C OAI21X1_39/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M10878 OAI21X1_39/Y OAI21X1_39/C OAI21X1_39/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10879 OAI21X1_39/Y OAI21X1_9/B OAI21X1_39/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M10880 OAI21X1_39/a_9_54# INVX2_232/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10881 OAI21X1_39/a_2_6# OAI21X1_9/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10882 gnd NOR2X1_2/A XNOR2X1_4/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M10883 XNOR2X1_4/Y NOR2X1_2/A XNOR2X1_4/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M10884 XNOR2X1_4/a_12_41# FAX1_2/YS gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10885 XNOR2X1_4/a_18_54# XNOR2X1_4/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M10886 XNOR2X1_4/a_35_6# XNOR2X1_4/a_2_6# XNOR2X1_4/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10887 XNOR2X1_4/a_18_6# XNOR2X1_4/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10888 vdd NOR2X1_2/A XNOR2X1_4/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M10889 vdd FAX1_2/YS XNOR2X1_4/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M10890 XNOR2X1_4/Y XNOR2X1_4/a_2_6# XNOR2X1_4/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M10891 XNOR2X1_4/a_35_54# NOR2X1_2/A XNOR2X1_4/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M10892 XNOR2X1_4/a_12_41# FAX1_2/YS vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10893 gnd FAX1_2/YS XNOR2X1_4/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10894 DFFNEGX1_50/a_76_6# BUFX2_14/Y DFFNEGX1_50/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M10895 gnd BUFX2_14/Y DFFNEGX1_50/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M10896 DFFNEGX1_50/a_66_6# DFFNEGX1_50/a_2_6# DFFNEGX1_50/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10897 out_temp_decoded[16] DFFNEGX1_50/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10898 DFFNEGX1_50/a_23_6# BUFX2_14/Y DFFNEGX1_50/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M10899 DFFNEGX1_50/a_23_6# DFFNEGX1_50/a_2_6# DFFNEGX1_50/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M10900 gnd DFFNEGX1_50/a_34_4# DFFNEGX1_50/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10901 vdd DFFNEGX1_50/a_34_4# DFFNEGX1_50/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M10902 DFFNEGX1_50/a_61_74# DFFNEGX1_50/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10903 DFFNEGX1_50/a_34_4# DFFNEGX1_50/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10904 DFFNEGX1_50/a_34_4# DFFNEGX1_50/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M10905 vdd out_temp_decoded[16] DFFNEGX1_50/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10906 gnd out_temp_decoded[16] DFFNEGX1_50/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10907 DFFNEGX1_50/a_61_6# DFFNEGX1_50/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10908 DFFNEGX1_50/a_76_84# DFFNEGX1_50/a_2_6# DFFNEGX1_50/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M10909 out_temp_decoded[16] DFFNEGX1_50/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10910 vdd BUFX2_14/Y DFFNEGX1_50/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M10911 DFFNEGX1_50/a_31_6# DFFNEGX1_50/a_2_6# DFFNEGX1_50/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10912 DFFNEGX1_50/a_66_6# BUFX2_14/Y DFFNEGX1_50/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10913 DFFNEGX1_50/a_17_74# OAI21X1_98/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10914 DFFNEGX1_50/a_31_74# BUFX2_14/Y DFFNEGX1_50/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10915 DFFNEGX1_50/a_17_6# OAI21X1_98/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10916 DFFNEGX1_61/a_76_6# BUFX2_13/Y DFFNEGX1_61/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M10917 gnd BUFX2_13/Y DFFNEGX1_61/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M10918 DFFNEGX1_61/a_66_6# DFFNEGX1_61/a_2_6# DFFNEGX1_61/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10919 out_temp_decoded[5] DFFNEGX1_61/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10920 DFFNEGX1_61/a_23_6# BUFX2_13/Y DFFNEGX1_61/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M10921 DFFNEGX1_61/a_23_6# DFFNEGX1_61/a_2_6# DFFNEGX1_61/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M10922 gnd DFFNEGX1_61/a_34_4# DFFNEGX1_61/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10923 vdd DFFNEGX1_61/a_34_4# DFFNEGX1_61/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M10924 DFFNEGX1_61/a_61_74# DFFNEGX1_61/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10925 DFFNEGX1_61/a_34_4# DFFNEGX1_61/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10926 DFFNEGX1_61/a_34_4# DFFNEGX1_61/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M10927 vdd out_temp_decoded[5] DFFNEGX1_61/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10928 gnd out_temp_decoded[5] DFFNEGX1_61/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10929 DFFNEGX1_61/a_61_6# DFFNEGX1_61/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10930 DFFNEGX1_61/a_76_84# DFFNEGX1_61/a_2_6# DFFNEGX1_61/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M10931 out_temp_decoded[5] DFFNEGX1_61/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10932 vdd BUFX2_13/Y DFFNEGX1_61/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M10933 DFFNEGX1_61/a_31_6# DFFNEGX1_61/a_2_6# DFFNEGX1_61/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10934 DFFNEGX1_61/a_66_6# BUFX2_13/Y DFFNEGX1_61/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10935 DFFNEGX1_61/a_17_74# OAI21X1_87/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10936 DFFNEGX1_61/a_31_74# BUFX2_13/Y DFFNEGX1_61/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10937 DFFNEGX1_61/a_17_6# OAI21X1_87/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10938 DFFNEGX1_94/a_76_6# BUFX2_10/Y DFFNEGX1_94/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M10939 gnd BUFX2_10/Y DFFNEGX1_94/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M10940 DFFNEGX1_94/a_66_6# DFFNEGX1_94/a_2_6# DFFNEGX1_94/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10941 out_global_score[0] DFFNEGX1_94/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10942 DFFNEGX1_94/a_23_6# BUFX2_10/Y DFFNEGX1_94/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M10943 DFFNEGX1_94/a_23_6# DFFNEGX1_94/a_2_6# DFFNEGX1_94/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M10944 gnd DFFNEGX1_94/a_34_4# DFFNEGX1_94/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10945 vdd DFFNEGX1_94/a_34_4# DFFNEGX1_94/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M10946 DFFNEGX1_94/a_61_74# DFFNEGX1_94/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10947 DFFNEGX1_94/a_34_4# DFFNEGX1_94/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10948 DFFNEGX1_94/a_34_4# DFFNEGX1_94/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M10949 vdd out_global_score[0] DFFNEGX1_94/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10950 gnd out_global_score[0] DFFNEGX1_94/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10951 DFFNEGX1_94/a_61_6# DFFNEGX1_94/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10952 DFFNEGX1_94/a_76_84# DFFNEGX1_94/a_2_6# DFFNEGX1_94/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M10953 out_global_score[0] DFFNEGX1_94/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10954 vdd BUFX2_10/Y DFFNEGX1_94/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M10955 DFFNEGX1_94/a_31_6# DFFNEGX1_94/a_2_6# DFFNEGX1_94/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10956 DFFNEGX1_94/a_66_6# BUFX2_10/Y DFFNEGX1_94/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10957 DFFNEGX1_94/a_17_74# INVX2_216/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10958 DFFNEGX1_94/a_31_74# BUFX2_10/Y DFFNEGX1_94/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10959 DFFNEGX1_94/a_17_6# INVX2_216/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10960 DFFNEGX1_83/a_76_6# BUFX2_11/Y DFFNEGX1_83/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M10961 gnd BUFX2_11/Y DFFNEGX1_83/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M10962 DFFNEGX1_83/a_66_6# DFFNEGX1_83/a_2_6# DFFNEGX1_83/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10963 out_temp_cleared[8] DFFNEGX1_83/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10964 DFFNEGX1_83/a_23_6# BUFX2_11/Y DFFNEGX1_83/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M10965 DFFNEGX1_83/a_23_6# DFFNEGX1_83/a_2_6# DFFNEGX1_83/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M10966 gnd DFFNEGX1_83/a_34_4# DFFNEGX1_83/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10967 vdd DFFNEGX1_83/a_34_4# DFFNEGX1_83/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M10968 DFFNEGX1_83/a_61_74# DFFNEGX1_83/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10969 DFFNEGX1_83/a_34_4# DFFNEGX1_83/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10970 DFFNEGX1_83/a_34_4# DFFNEGX1_83/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M10971 vdd out_temp_cleared[8] DFFNEGX1_83/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10972 gnd out_temp_cleared[8] DFFNEGX1_83/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10973 DFFNEGX1_83/a_61_6# DFFNEGX1_83/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10974 DFFNEGX1_83/a_76_84# DFFNEGX1_83/a_2_6# DFFNEGX1_83/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M10975 out_temp_cleared[8] DFFNEGX1_83/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10976 vdd BUFX2_11/Y DFFNEGX1_83/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M10977 DFFNEGX1_83/a_31_6# DFFNEGX1_83/a_2_6# DFFNEGX1_83/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10978 DFFNEGX1_83/a_66_6# BUFX2_11/Y DFFNEGX1_83/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10979 DFFNEGX1_83/a_17_74# OAI22X1_20/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10980 DFFNEGX1_83/a_31_74# BUFX2_11/Y DFFNEGX1_83/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M10981 DFFNEGX1_83/a_17_6# OAI22X1_20/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10982 DFFNEGX1_72/a_76_6# BUFX2_12/Y DFFNEGX1_72/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M10983 gnd BUFX2_12/Y DFFNEGX1_72/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M10984 DFFNEGX1_72/a_66_6# DFFNEGX1_72/a_2_6# DFFNEGX1_72/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10985 out_temp_cleared[19] DFFNEGX1_72/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10986 DFFNEGX1_72/a_23_6# BUFX2_12/Y DFFNEGX1_72/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M10987 DFFNEGX1_72/a_23_6# DFFNEGX1_72/a_2_6# DFFNEGX1_72/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M10988 gnd DFFNEGX1_72/a_34_4# DFFNEGX1_72/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10989 vdd DFFNEGX1_72/a_34_4# DFFNEGX1_72/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M10990 DFFNEGX1_72/a_61_74# DFFNEGX1_72/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M10991 DFFNEGX1_72/a_34_4# DFFNEGX1_72/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M10992 DFFNEGX1_72/a_34_4# DFFNEGX1_72/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M10993 vdd out_temp_cleared[19] DFFNEGX1_72/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M10994 gnd out_temp_cleared[19] DFFNEGX1_72/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10995 DFFNEGX1_72/a_61_6# DFFNEGX1_72/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M10996 DFFNEGX1_72/a_76_84# DFFNEGX1_72/a_2_6# DFFNEGX1_72/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M10997 out_temp_cleared[19] DFFNEGX1_72/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M10998 vdd BUFX2_12/Y DFFNEGX1_72/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M10999 DFFNEGX1_72/a_31_6# DFFNEGX1_72/a_2_6# DFFNEGX1_72/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M11000 DFFNEGX1_72/a_66_6# BUFX2_12/Y DFFNEGX1_72/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11001 DFFNEGX1_72/a_17_74# OAI22X1_9/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11002 DFFNEGX1_72/a_31_74# BUFX2_12/Y DFFNEGX1_72/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11003 DFFNEGX1_72/a_17_6# OAI22X1_9/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M11004 vdd out_global_score[22] HAX1_8/a_2_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.2n ps=100u
M11005 HAX1_8/a_41_74# HAX1_8/a_2_74# vdd vdd pfet w=20 l=2
+  ad=0.22n pd=92u as=0 ps=0
M11006 HAX1_8/a_9_6# out_global_score[22] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M11007 HAX1_8/a_41_74# HAX1_8/B HAX1_8/a_38_6# Gnd nfet w=20 l=2
+  ad=0.12n pd=52u as=0.216n ps=0.102m
M11008 vdd out_global_score[22] HAX1_8/a_49_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M11009 vdd HAX1_8/a_2_74# HAX1_7/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M11010 HAX1_8/a_38_6# HAX1_8/a_2_74# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11011 HAX1_8/YS HAX1_8/a_41_74# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M11012 HAX1_8/a_38_6# out_global_score[22] HAX1_8/a_41_74# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11013 HAX1_8/YS HAX1_8/a_41_74# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M11014 HAX1_8/a_2_74# HAX1_8/B vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11015 HAX1_8/a_2_74# HAX1_8/B HAX1_8/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M11016 HAX1_8/a_49_54# HAX1_8/B HAX1_8/a_41_74# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M11017 gnd HAX1_8/a_2_74# HAX1_7/B Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M11018 AND2X2_4/a_2_6# OR2X1_9/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M11019 AND2X2_4/a_9_6# OR2X1_9/Y AND2X2_4/a_2_6# Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=100p ps=50u
M11020 OR2X1_8/B AND2X2_4/a_2_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M11021 OR2X1_8/B AND2X2_4/a_2_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M11022 vdd out_temp_data_in[2] AND2X2_4/a_2_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11023 gnd out_temp_data_in[2] AND2X2_4/a_9_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11024 INVX2_209/Y INVX2_209/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M11025 INVX2_209/Y INVX2_209/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M11026 gnd HAX1_42/YS MUX2X1_16/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M11027 MUX2X1_16/a_17_50# HAX1_42/A vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M11028 MUX2X1_16/Y OR2X1_3/Y MUX2X1_16/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M11029 MUX2X1_16/a_30_54# MUX2X1_16/a_2_10# MUX2X1_16/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M11030 MUX2X1_16/a_17_10# HAX1_42/A gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M11031 vdd OR2X1_3/Y MUX2X1_16/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M11032 MUX2X1_16/a_30_10# OR2X1_3/Y MUX2X1_16/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M11033 gnd OR2X1_3/Y MUX2X1_16/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M11034 vdd HAX1_42/YS MUX2X1_16/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M11035 MUX2X1_16/Y MUX2X1_16/a_2_10# MUX2X1_16/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11036 gnd XNOR2X1_3/Y MUX2X1_27/a_30_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M11037 MUX2X1_27/a_17_50# MUX2X1_27/B vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M11038 MUX2X1_27/Y OR2X1_1/Y MUX2X1_27/a_17_50# vdd pfet w=40 l=2
+  ad=0.248n pd=100u as=0 ps=0
M11039 MUX2X1_27/a_30_54# MUX2X1_27/a_2_10# MUX2X1_27/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M11040 MUX2X1_27/a_17_10# MUX2X1_27/B gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M11041 vdd OR2X1_1/Y MUX2X1_27/a_2_10# vdd pfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M11042 MUX2X1_27/a_30_10# OR2X1_1/Y MUX2X1_27/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M11043 gnd OR2X1_1/Y MUX2X1_27/a_2_10# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=50p ps=30u
M11044 vdd XNOR2X1_3/Y MUX2X1_27/a_30_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M11045 MUX2X1_27/Y MUX2X1_27/a_2_10# MUX2X1_27/a_17_10# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11046 DFFNEGX1_140/a_76_6# INVX2_259/Y DFFNEGX1_140/a_66_6# Gnd nfet w=10 l=2
+  ad=29.999998p pd=26u as=80p ps=36u
M11047 gnd INVX2_259/Y DFFNEGX1_140/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M11048 DFFNEGX1_140/a_66_6# DFFNEGX1_140/a_2_6# DFFNEGX1_140/a_61_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M11049 out_decode DFFNEGX1_140/a_66_6# gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M11050 DFFNEGX1_140/a_23_6# INVX2_259/Y DFFNEGX1_140/a_17_6# Gnd nfet w=10 l=2
+  ad=59.999996p pd=32u as=40p ps=28u
M11051 DFFNEGX1_140/a_23_6# DFFNEGX1_140/a_2_6# DFFNEGX1_140/a_17_74# vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=80p ps=48u
M11052 gnd DFFNEGX1_140/a_34_4# DFFNEGX1_140/a_31_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M11053 vdd DFFNEGX1_140/a_34_4# DFFNEGX1_140/a_31_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=80p ps=48u
M11054 DFFNEGX1_140/a_61_74# DFFNEGX1_140/a_34_4# vdd vdd pfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M11055 DFFNEGX1_140/a_34_4# DFFNEGX1_140/a_23_6# vdd vdd pfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M11056 DFFNEGX1_140/a_34_4# DFFNEGX1_140/a_23_6# gnd Gnd nfet w=10 l=2
+  ad=50p pd=30u as=0 ps=0
M11057 vdd out_decode DFFNEGX1_140/a_76_84# vdd pfet w=10 l=2
+  ad=0 pd=0 as=29.999998p ps=26u
M11058 gnd out_decode DFFNEGX1_140/a_76_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M11059 DFFNEGX1_140/a_61_6# DFFNEGX1_140/a_34_4# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M11060 DFFNEGX1_140/a_76_84# DFFNEGX1_140/a_2_6# DFFNEGX1_140/a_66_6# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0.15n ps=56u
M11061 out_decode DFFNEGX1_140/a_66_6# vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M11062 vdd INVX2_259/Y DFFNEGX1_140/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M11063 DFFNEGX1_140/a_31_6# DFFNEGX1_140/a_2_6# DFFNEGX1_140/a_23_6# Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M11064 DFFNEGX1_140/a_66_6# INVX2_259/Y DFFNEGX1_140/a_61_74# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11065 DFFNEGX1_140/a_17_74# OAI21X1_158/Y vdd vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11066 DFFNEGX1_140/a_31_74# INVX2_259/Y DFFNEGX1_140/a_23_6# vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11067 DFFNEGX1_140/a_17_6# OAI21X1_158/Y gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M11068 OAI21X1_13/C out_mines[19] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M11069 NAND2X1_20/a_9_6# out_mines[19] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M11070 vdd INVX2_239/Y OAI21X1_13/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11071 OAI21X1_13/C INVX2_239/Y NAND2X1_20/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M11072 OAI21X1_30/B NOR2X1_62/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M11073 NAND2X1_31/a_9_6# NOR2X1_62/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M11074 vdd NOR2X1_65/A OAI21X1_30/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11075 OAI21X1_30/B NOR2X1_65/A NAND2X1_31/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M11076 OAI21X1_45/C out_mines[3] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M11077 NAND2X1_42/a_9_6# out_mines[3] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M11078 vdd INVX2_243/Y OAI21X1_45/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11079 OAI21X1_45/C INVX2_243/Y NAND2X1_42/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M11080 OAI21X1_88/C NOR2X1_38/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M11081 NAND2X1_75/a_9_6# NOR2X1_38/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M11082 vdd BUFX2_20/Y OAI21X1_88/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11083 OAI21X1_88/C BUFX2_20/Y NAND2X1_75/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M11084 OAI21X1_72/B OAI22X1_1/D vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M11085 NAND2X1_64/a_9_6# OAI22X1_1/D gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M11086 vdd INVX2_75/Y OAI21X1_72/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11087 OAI21X1_72/B INVX2_75/Y NAND2X1_64/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M11088 OAI21X1_99/C NOR2X1_51/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M11089 NAND2X1_86/a_9_6# NOR2X1_51/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M11090 vdd BUFX2_21/Y OAI21X1_99/C vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11091 OAI21X1_99/C BUFX2_21/Y NAND2X1_86/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M11092 OAI21X1_57/B OR2X1_13/Y vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M11093 NAND2X1_53/a_9_6# OR2X1_13/Y gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M11094 vdd AND2X2_8/A OAI21X1_57/B vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11095 OAI21X1_57/B AND2X2_8/A NAND2X1_53/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M11096 NAND2X1_97/Y in_data[1] vdd vdd pfet w=20 l=2
+  ad=0.12n pd=52u as=0 ps=0
M11097 NAND2X1_97/a_9_6# in_data[1] gnd Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M11098 vdd NOR2X1_107/Y NAND2X1_97/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11099 NAND2X1_97/Y NOR2X1_107/Y NAND2X1_97/a_9_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M11100 gnd out_temp_cleared[23] AOI22X1_51/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M11101 NAND3X1_46/A out_mines[22] AOI22X1_51/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M11102 AOI22X1_51/a_11_6# out_temp_cleared[22] gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11103 AOI22X1_51/a_2_54# out_mines[22] vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M11104 AOI22X1_51/a_28_6# out_mines[23] NAND3X1_46/A Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11105 vdd out_temp_cleared[22] AOI22X1_51/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M11106 NAND3X1_46/A out_mines[23] AOI22X1_51/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M11107 AOI22X1_51/a_2_54# out_temp_cleared[23] NAND3X1_46/A vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M11108 gnd out_temp_decoded[4] AOI22X1_40/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M11109 OAI21X1_70/C out_mines[3] AOI22X1_40/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M11110 AOI22X1_40/a_11_6# out_temp_decoded[3] gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11111 AOI22X1_40/a_2_54# out_mines[3] vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M11112 AOI22X1_40/a_28_6# out_mines[4] OAI21X1_70/C Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11113 vdd out_temp_decoded[3] AOI22X1_40/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M11114 OAI21X1_70/C out_mines[4] AOI22X1_40/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M11115 AOI22X1_40/a_2_54# out_temp_decoded[4] OAI21X1_70/C vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M11116 gnd INVX2_34/A AOI22X1_73/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M11117 AOI22X1_73/Y INVX2_34/Y AOI22X1_73/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M11118 AOI22X1_73/a_11_6# AOI22X1_73/A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11119 AOI22X1_73/a_2_54# INVX2_34/Y vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M11120 AOI22X1_73/a_28_6# INVX2_23/Y AOI22X1_73/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11121 vdd AOI22X1_73/A AOI22X1_73/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M11122 AOI22X1_73/Y INVX2_23/Y AOI22X1_73/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M11123 AOI22X1_73/a_2_54# INVX2_34/A AOI22X1_73/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M11124 gnd NOR2X1_111/Y AOI22X1_62/a_28_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=59.999996p ps=46u
M11125 AOI22X1_62/Y out_mines[9] AOI22X1_62/a_11_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M11126 AOI22X1_62/a_11_6# NOR2X1_112/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11127 AOI22X1_62/a_2_54# out_mines[9] vdd vdd pfet w=40 l=2
+  ad=0.64n pd=0.272m as=0 ps=0
M11128 AOI22X1_62/a_28_6# out_mines[10] AOI22X1_62/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11129 vdd NOR2X1_112/Y AOI22X1_62/a_2_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M11130 AOI22X1_62/Y out_mines[10] AOI22X1_62/a_2_54# vdd pfet w=40 l=2
+  ad=0.24n pd=92u as=0 ps=0
M11131 AOI22X1_62/a_2_54# NOR2X1_111/Y AOI22X1_62/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M11132 gnd INVX2_8/Y OAI22X1_2/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.32n ps=0.152m
M11133 OAI22X1_2/a_2_6# INVX2_28/Y OAI22X1_2/Y Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.12n ps=52u
M11134 OAI22X1_2/Y OAI22X1_2/D OAI22X1_2/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11135 OAI22X1_2/Y OAI22X1_2/B OAI22X1_2/a_9_54# vdd pfet w=40 l=2
+  ad=0.48n pd=0.104m as=0.12n ps=86u
M11136 OAI22X1_2/a_28_54# OAI22X1_2/D OAI22X1_2/Y vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M11137 OAI22X1_2/a_9_54# INVX2_8/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M11138 OAI22X1_2/a_2_6# OAI22X1_2/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11139 vdd INVX2_28/Y OAI22X1_2/a_28_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M11140 INVX2_11/Y out_mines[15] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M11141 INVX2_11/Y out_mines[15] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M11142 INVX2_22/Y out_mines[17] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M11143 INVX2_22/Y out_mines[17] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M11144 INVX2_33/Y INVX2_33/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M11145 INVX2_33/Y INVX2_33/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M11146 INVX2_44/Y INVX2_44/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M11147 INVX2_44/Y INVX2_44/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M11148 INVX2_77/Y out_temp_decoded[6] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M11149 INVX2_77/Y out_temp_decoded[6] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M11150 INVX2_66/Y out_temp_decoded[15] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M11151 INVX2_66/Y out_temp_decoded[15] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M11152 INVX2_55/Y out_temp_decoded[24] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M11153 INVX2_55/Y out_temp_decoded[24] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M11154 INVX2_88/Y INVX2_88/A gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M11155 INVX2_88/Y INVX2_88/A vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M11156 INVX2_99/Y out_temp_cleared[14] gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M11157 INVX2_99/Y out_temp_cleared[14] vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M11158 gnd INVX2_180/Y OAI21X1_18/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M11159 vdd BUFX2_19/Y INVX2_220/A vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M11160 INVX2_220/A BUFX2_19/Y OAI21X1_18/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M11161 INVX2_220/A NAND3X1_8/Y OAI21X1_18/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M11162 OAI21X1_18/a_9_54# INVX2_180/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M11163 OAI21X1_18/a_2_6# NAND3X1_8/Y gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11164 gnd INVX2_241/Y OAI21X1_29/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=0.102m
M11165 vdd OAI21X1_29/C OAI21X1_29/Y vdd pfet w=20 l=2
+  ad=0 pd=0 as=0.22n ps=92u
M11166 OAI21X1_29/Y OAI21X1_29/C OAI21X1_29/a_2_6# Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M11167 OAI21X1_29/Y OAI21X1_9/B OAI21X1_29/a_9_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M11168 OAI21X1_29/a_9_54# INVX2_241/Y vdd vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M11169 OAI21X1_29/a_2_6# OAI21X1_9/B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11170 gnd XNOR2X1_5/A XNOR2X1_5/a_2_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=100p ps=50u
M11171 XNOR2X1_5/Y XNOR2X1_5/A XNOR2X1_5/a_18_6# Gnd nfet w=20 l=2
+  ad=0.2n pd=60u as=59.999996p ps=46u
M11172 XNOR2X1_5/a_12_41# NOR2X1_2/Y gnd Gnd nfet w=20 l=2
+  ad=100p pd=50u as=0 ps=0
M11173 XNOR2X1_5/a_18_54# XNOR2X1_5/a_12_41# vdd vdd pfet w=40 l=2
+  ad=0.12n pd=86u as=0 ps=0
M11174 XNOR2X1_5/a_35_6# XNOR2X1_5/a_2_6# XNOR2X1_5/Y Gnd nfet w=20 l=2
+  ad=59.999996p pd=46u as=0 ps=0
M11175 XNOR2X1_5/a_18_6# XNOR2X1_5/a_12_41# gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M11176 vdd XNOR2X1_5/A XNOR2X1_5/a_2_6# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.2n ps=90u
M11177 vdd NOR2X1_2/Y XNOR2X1_5/a_35_54# vdd pfet w=40 l=2
+  ad=0 pd=0 as=0.12n ps=86u
M11178 XNOR2X1_5/Y XNOR2X1_5/a_2_6# XNOR2X1_5/a_18_54# vdd pfet w=40 l=2
+  ad=0.4n pd=100u as=0 ps=0
M11179 XNOR2X1_5/a_35_54# XNOR2X1_5/A XNOR2X1_5/Y vdd pfet w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M11180 XNOR2X1_5/a_12_41# NOR2X1_2/Y vdd vdd pfet w=40 l=2
+  ad=0.2n pd=90u as=0 ps=0
M11181 gnd NOR2X1_2/Y XNOR2X1_5/a_35_6# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
C0 vdd out_temp_data_in[3] 8.572948f
C1 vdd INVX2_57/Y 3.08349f
C2 OAI22X1_52/B vdd 3.51999f
C3 vdd INVX2_14/Y 2.67606f
C4 vdd INVX2_119/Y 2.18295f
C5 vdd OAI22X1_52/D 2.32155f
C6 INVX2_257/Y vdd 4.772521f
C7 vdd AND2X2_14/B 2.81034f
C8 vdd OAI21X1_1/B 13.764058f
C9 vdd out_mines[7] 10.365208f
C10 gnd BUFX2_15/Y 2.47932f
C11 OAI21X1_1/A vdd 6.614461f
C12 gnd INVX2_259/Y 2.08161f
C13 INVX2_221/Y vdd 2.01168f
C14 vdd NOR2X1_66/B 6.21009f
C15 vdd OR2X1_0/Y 5.06583f
C16 vdd XNOR2X1_7/A 2.40174f
C17 vdd out_global_score[24] 2.17575f
C18 vdd INVX2_120/A 2.52198f
C19 out_mines[9] vdd 4.622311f
C20 vdd out_state_main[3] 2.96793f
C21 vdd AND2X2_15/Y 2.1996f
C22 gnd BUFX2_25/Y 2.943f
C23 INVX2_65/Y vdd 3.68721f
C24 vdd out_temp_mine_cnt[1] 2.07387f
C25 vdd out_temp_mine_cnt[2] 2.07945f
C26 vdd BUFX2_11/Y 15.124854f
C27 OAI22X1_63/B vdd 3.20931f
C28 vdd out_global_score[1] 2.30418f
C29 AOI21X1_2/A vdd 4.07007f
C30 vdd OAI21X1_9/B 9.294836f
C31 vdd BUFX2_1/Y 2.8971f
C32 vdd out_mines[10] 8.597157f
C33 BUFX2_5/Y vdd 13.448337f
C34 vdd NOR2X1_86/A 2.96451f
C35 OAI21X1_8/A vdd 4.45293f
C36 vdd INVX2_23/Y 2.94894f
C37 INVX2_258/Y vdd 7.66809f
C38 gnd BUFX2_12/Y 2.400211f
C39 vdd out_state_main[2] 3.4695f
C40 BUFX2_10/Y vdd 15.429412f
C41 vdd NOR2X1_107/Y 4.23054f
C42 BUFX2_21/A vdd 2.0736f
C43 INVX2_52/Y vdd 2.66742f
C44 vdd out_state_main[0] 3.26385f
C45 vdd out_place_done 2.87091f
C46 vdd out_display_done 2.66472f
C47 vdd INVX2_82/Y 2.44773f
C48 out_alu vdd 2.87631f
C49 vdd BUFX2_15/Y 16.587536f
C50 vdd BUFX2_23/Y 6.86115f
C51 out_global_score[14] vdd 2.19141f
C52 INVX2_259/Y vdd 16.639463f
C53 vdd INVX2_19/Y 2.09349f
C54 vdd out_start 3.97953f
C55 vdd OAI22X1_63/D 2.4102f
C56 INVX2_2/Y vdd 2.40633f
C57 vdd INVX2_81/Y 2.20338f
C58 vdd OAI22X1_87/D 2.27376f
C59 vdd BUFX2_13/Y 14.846666f
C60 vdd out_temp_data_in[1] 9.251459f
C61 vdd INVX2_10/Y 2.28312f
C62 gnd out_mines[1] 2.580211f
C63 vdd INVX2_32/Y 2.59155f
C64 out_temp_cleared[23] vdd 2.29635f
C65 vdd INVX2_8/Y 3.26952f
C66 vdd NOR2X1_56/B 3.976561f
C67 vdd INVX2_125/Y 2.00871f
C68 vdd out_temp_cleared[14] 2.16207f
C69 BUFX2_25/A vdd 3.56427f
C70 vdd BUFX2_25/Y 3.51351f
C71 out_decode vdd 2.70801f
C72 vdd out_mines[6] 7.53696f
C73 vdd NOR2X1_110/B 2.6118f
C74 vdd INVX2_77/Y 2.69982f
C75 vdd INVX2_255/Y 3.33531f
C76 vdd NOR2X1_27/B 2.14722f
C77 vdd BUFX2_18/Y 10.930049f
C78 out_temp_cleared[12] vdd 2.35368f
C79 vdd out_mines[0] 8.20503f
C80 INVX2_66/Y vdd 2.39688f
C81 vdd out_temp_mine_cnt[0] 2.43729f
C82 vdd INVX2_116/Y 2.04561f
C83 vdd out_global_score[29] 2.11851f
C84 vdd OR2X1_5/Y 5.171311f
C85 NOR2X1_91/Y vdd 2.45772f
C86 OAI22X1_5/C vdd 8.700117f
C87 vdd out_global_score[3] 2.20635f
C88 vdd out_temp_cleared[10] 2.50065f
C89 vdd BUFX2_12/Y 15.600417f
C90 vdd OAI21X1_44/A 2.00646f
C91 NOR2X1_63/B vdd 4.60017f
C92 vdd out_mines[19] 8.01468f
C93 vdd out_state_main[1] 2.72997f
C94 gnd BUFX2_9/Y 3.310111f
C95 OAI22X1_76/B vdd 2.11797f
C96 vdd out_temp_decoded[24] 3.13092f
C97 vdd INVX2_0/A 2.28951f
C98 gnd out_temp_data_in[0] 2.831851f
C99 vdd OAI22X1_75/D 2.11194f
C100 vdd out_mines[13] 7.07445f
C101 vdd INVX2_54/Y 3.44223f
C102 vdd INVX2_79/Y 2.87568f
C103 vdd BUFX2_9/A 2.1519f
C104 vdd out_global_score[25] 2.17071f
C105 vdd out_global_score[16] 2.20743f
C106 vdd out_mines[22] 7.228799f
C107 vdd out_mines[15] 8.380259f
C108 gnd out_mines[17] 2.91447f
C109 INVX2_1/Y vdd 2.13075f
C110 out_mines[1] vdd 7.105411f
C111 vdd out_global_score[30] 2.24631f
C112 gnd BUFX2_3/Y 2.00196f
C113 vdd out_mines[24] 4.209301f
C114 vdd NOR2X1_7/Y 4.66992f
C115 vdd OR2X1_2/Y 5.017681f
C116 OAI21X1_83/C vdd 2.91033f
C117 vdd NOR2X1_67/Y 5.14395f
C118 INVX2_40/A vdd 5.28777f
C119 NOR2X1_84/A vdd 2.97063f
C120 NOR2X1_77/B vdd 3.3183f
C121 gnd OR2X1_11/A 2.45799f
C122 AND2X2_17/A vdd 2.19564f
C123 INVX2_35/Y vdd 2.5272f
C124 vdd NAND3X1_8/Y 2.94336f
C125 INVX2_131/Y vdd 2.40327f
C126 INVX2_251/Y vdd 7.497901f
C127 gnd BUFX2_17/Y 2.23524f
C128 vdd OR2X1_6/A 6.63831f
C129 vdd OAI22X1_87/B 2.3661f
C130 vdd NAND3X1_7/Y 3.89754f
C131 vdd AND2X2_19/B 2.09295f
C132 vdd out_global_score[12] 2.28303f
C133 vdd AOI21X1_3/A 3.61449f
C134 vdd out_mines[12] 8.505089f
C135 vdd AND2X2_8/A 3.76299f
C136 vdd out_mines[5] 7.73613f
C137 vdd OR2X1_3/Y 4.94415f
C138 BUFX2_9/Y vdd 15.075175f
C139 vdd NOR2X1_125/Y 2.79216f
C140 vdd out_temp_data_in[0] 12.810232f
C141 vdd out_mines[18] 7.58322f
C142 NOR2X1_59/B vdd 2.41254f
C143 XOR2X1_29/B vdd 3.35664f
C144 gnd OR2X1_6/Y 2.00457f
C145 vdd NAND3X1_9/A 3.60243f
C146 vdd OAI22X1_88/B 3.464191f
C147 vdd out_mines[11] 11.545738f
C148 vdd BUFX2_19/A 4.222171f
C149 vdd BUFX2_24/Y 3.730861f
C150 vdd NOR2X1_47/B 2.98737f
C151 INVX2_117/Y vdd 3.17538f
C152 vdd out_display 3.47913f
C153 vdd out_mines[17] 8.58087f
C154 vdd NOR2X1_57/B 2.63448f
C155 vdd BUFX2_3/Y 3.85731f
C156 out_temp_cleared[20] vdd 2.53845f
C157 OR2X1_11/B vdd 5.14872f
C158 vdd OR2X1_1/Y 5.80932f
C159 vdd out_gameover 2.61207f
C160 out_global_score[18] vdd 2.11203f
C161 vdd out_mines[23] 9.894237f
C162 vdd INVX2_52/A 3.48318f
C163 vdd out_global_score[15] 2.35719f
C164 INVX2_127/A vdd 3.91851f
C165 vdd INVX2_26/Y 3.40065f
C166 vdd OAI22X1_64/D 2.40408f
C167 vdd BUFX2_21/Y 8.83809f
C168 vdd NOR2X1_78/A 2.29698f
C169 vdd OR2X1_11/A 10.498315f
C170 vdd out_temp_mine_cnt[3] 2.29149f
C171 vdd INVX2_15/Y 3.0042f
C172 out_temp_cleared[19] vdd 2.25f
C173 OAI21X1_90/C vdd 2.69505f
C174 vdd INVX2_130/Y 2.75022f
C175 BUFX2_17/Y vdd 18.440094f
C176 vdd out_alu_done 3.21723f
C177 vdd BUFX2_19/Y 9.102059f
C178 vdd INVX2_67/Y 2.54808f
C179 gnd out_temp_data_in[3] 3.836071f
C180 vdd INVX2_16/Y 3.63753f
C181 gnd vdd 8.424f
C182 out_temp_cleared[13] vdd 2.23911f
C183 OAI22X1_75/B vdd 2.97945f
C184 vdd INVX2_70/Y 2.98188f
C185 vdd out_temp_cleared[21] 2.73123f
C186 vdd HAX1_31/B 2.29671f
C187 out_mines[21] vdd 5.56875f
C188 vdd INVX2_117/A 2.59947f
C189 vdd OAI22X1_64/B 3.31983f
C190 vdd INVX2_30/Y 4.743001f
C191 vdd NOR2X1_77/A 2.03742f
C192 vdd NOR2X1_52/B 2.31255f
C193 out_temp_data_in[4] vdd 9.310227f
C194 vdd OR2X1_4/Y 5.759191f
C195 vdd out_mines[4] 8.800016f
C196 out_mines[8] vdd 7.39989f
C197 INVX2_38/Y vdd 2.90934f
C198 vdd INVX2_31/Y 3.62601f
C199 gnd BUFX2_11/Y 2.546371f
C200 BUFX2_16/Y vdd 20.495787f
C201 HAX1_42/A vdd 2.03796f
C202 vdd OAI22X1_51/B 2.74806f
C203 vdd out_mines[3] 8.458919f
C204 vdd INVX2_119/A 3.93039f
C205 gnd OAI21X1_9/B 2.439811f
C206 vdd BUFX2_22/Y 6.085891f
C207 gnd out_mines[10] 2.687851f
C208 out_mines[20] vdd 7.63497f
C209 vdd XOR2X1_28/A 4.34583f
C210 BUFX2_5/Y gnd 4.744621f
C211 NOR2X1_66/A vdd 2.44701f
C212 INVX2_58/A vdd 2.59236f
C213 vdd INVX2_217/A 3.32964f
C214 vdd INVX2_22/Y 3.32838f
C215 vdd INVX2_85/Y 3.38796f
C216 vdd out_temp_data_in[2] 14.006783f
C217 NOR2X1_22/B vdd 3.482371f
C218 XOR2X1_4/Y vdd 3.480661f
C219 vdd BUFX2_8/Y 2.7864f
C220 vdd BUFX2_20/Y 10.196368f
C221 vdd BUFX2_14/Y 15.145916f
C222 out_mines[14] vdd 6.74928f
C223 vdd NOR2X1_17/B 2.81709f
C224 INVX2_74/Y vdd 2.96748f
C225 vdd out_global_score[10] 2.19339f
C226 vdd XOR2X1_3/Y 3.14721f
C227 vdd NOR2X1_104/B 2.9952f
C228 gnd BUFX2_10/Y 3.819241f
C229 vdd out_mines[2] 14.492783f
C230 OAI21X1_89/C vdd 3.07971f
C231 vdd out_mines[16] 8.785346f
C232 out_temp_mine_cnt[2] 0 29.93778f **FLOATING
C233 out_temp_cleared[8] 0 12.290309f **FLOATING
C234 out_temp_cleared[10] 0 28.74681f **FLOATING
C235 out_temp_decoded[6] 0 15.801449f **FLOATING
C236 out_temp_decoded[9] 0 32.27412f **FLOATING
C237 out_global_score[13] 0 21.72609f **FLOATING
C238 out_global_score[15] 0 21.20481f **FLOATING
C239 out_global_score[29] 0 22.59609f **FLOATING
C240 out_global_score[30] 0 21.468811f **FLOATING
C241 NOR2X1_78/A 0 21.102959f **FLOATING
C242 BUFX2_11/Y 0 0.165133p **FLOATING
C243 out_temp_cleared[17] 0 17.785053f **FLOATING
C244 BUFX2_12/Y 0 0.176761p **FLOATING
C245 out_temp_decoded[12] 0 30.712984f **FLOATING
C246 out_temp_decoded[17] 0 12.595651f **FLOATING
C247 out_mines[15] 0 96.09879f **FLOATING
C248 OR2X1_11/A 0 0.177082p **FLOATING
C249 BUFX2_25/Y 0 79.27437f **FLOATING
C250 OR2X1_15/B 0 17.9817f **FLOATING
C251 BUFX2_24/Y 0 89.24379f **FLOATING
C252 OAI21X1_155/Y 0 10.007521f **FLOATING
C253 OAI21X1_157/A 0 10.1586f **FLOATING
C254 INVX2_77/Y 0 34.500237f **FLOATING
C255 out_temp_cleared[9] 0 13.180049f **FLOATING
C256 AND2X2_17/Y 0 13.73721f **FLOATING
C257 INVX2_121/Y 0 8.258279f **FLOATING
C258 NOR2X1_94/B 0 12.79506f **FLOATING
C259 out_temp_cleared[14] 0 22.136969f **FLOATING
C260 OAI22X1_13/Y 0 11.12574f **FLOATING
C261 INVX2_98/Y 0 10.959781f **FLOATING
C262 out_temp_decoded[13] 0 25.80975f **FLOATING
C263 OAI21X1_78/C 0 12.06021f **FLOATING
C264 INVX2_70/Y 0 29.945099f **FLOATING
C265 INVX2_22/Y 0 32.557697f **FLOATING
C266 INVX2_26/Y 0 41.083134f **FLOATING
C267 NOR2X1_56/B 0 28.087797f **FLOATING
C268 NOR2X1_52/B 0 33.832592f **FLOATING
C269 INVX2_102/Y 0 12.536101f **FLOATING
C270 OAI21X1_92/C 0 10.527f **FLOATING
C271 AOI21X1_5/Y 0 19.609648f **FLOATING
C272 OAI22X1_1/D 0 25.368479f **FLOATING
C273 NAND3X1_35/Y 0 13.812449f **FLOATING
C274 BUFX2_20/Y 0 53.4941f **FLOATING
C275 NAND3X1_41/A 0 12.018849f **FLOATING
C276 NOR2X1_115/Y 0 10.448701f **FLOATING
C277 out_temp_cleared[7] 0 12.00843f **FLOATING
C278 OAI22X1_17/Y 0 10.308779f **FLOATING
C279 NOR2X1_58/A 0 15.77253f **FLOATING
C280 OAI21X1_95/Y 0 11.548019f **FLOATING
C281 INVX2_12/Y 0 8.05614f **FLOATING
C282 NOR2X1_94/Y 0 10.099861f **FLOATING
C283 NOR2X1_116/Y 0 22.831558f **FLOATING
C284 OAI21X1_89/Y 0 14.31198f **FLOATING
C285 NOR2X1_57/Y 0 10.417381f **FLOATING
C286 out_mines[17] 0 0.129715p **FLOATING
C287 OAI21X1_92/Y 0 9.631861f **FLOATING
C288 NOR2X1_36/Y 0 11.433841f **FLOATING
C289 INVX2_54/Y 0 57.161476f **FLOATING
C290 INVX2_97/Y 0 9.80868f **FLOATING
C291 out_temp_cleared[11] 0 18.863308f **FLOATING
C292 OAI21X1_160/Y 0 10.630321f **FLOATING
C293 NOR2X1_87/B 0 12.303479f **FLOATING
C294 out_mines[10] 0 0.12941p **FLOATING
C295 NOR2X1_46/Y 0 10.455f **FLOATING
C296 OAI21X1_159/Y 0 12.042662f **FLOATING
C297 INVX2_7/Y 0 12.807f **FLOATING
C298 NOR2X1_45/Y 0 11.2953f **FLOATING
C299 OAI21X1_88/C 0 12.35646f **FLOATING
C300 NOR2X1_44/Y 0 8.899321f **FLOATING
C301 OAI21X1_104/Y 0 11.412059f **FLOATING
C302 NOR2X1_85/B 0 9.90846f **FLOATING
C303 INVX2_16/Y 0 45.65755f **FLOATING
C304 NAND2X1_91/Y 0 12.01968f **FLOATING
C305 out_mines[11] 0 0.112077p **FLOATING
C306 OAI21X1_106/Y 0 13.2999f **FLOATING
C307 OAI22X1_1/Y 0 11.31066f **FLOATING
C308 out_temp_decoded[24] 0 33.53814f **FLOATING
C309 INVX2_57/Y 0 25.37553f **FLOATING
C310 OAI22X1_20/Y 0 10.308781f **FLOATING
C311 BUFX2_23/A 0 24.266521f **FLOATING
C312 OAI21X1_87/C 0 9.351542f **FLOATING
C313 INVX2_61/Y 0 11.81928f **FLOATING
C314 INVX2_91/Y 0 11.295599f **FLOATING
C315 out_temp_decoded[5] 0 24.90014f **FLOATING
C316 OAI21X1_103/Y 0 11.16996f **FLOATING
C317 INVX2_76/Y 0 15.38988f **FLOATING
C318 OAI21X1_101/Y 0 11.939011f **FLOATING
C319 out_temp_decoded[21] 0 16.442013f **FLOATING
C320 out_mines[22] 0 80.22717f **FLOATING
C321 INVX2_85/Y 0 45.630135f **FLOATING
C322 INVX2_130/Y 0 46.39129f **FLOATING
C323 AOI21X1_5/C 0 9.693181f **FLOATING
C324 OAI22X1_9/Y 0 12.574679f **FLOATING
C325 INVX2_82/Y 0 23.727898f **FLOATING
C326 INVX2_80/Y 0 15.24826f **FLOATING
C327 INVX2_21/Y 0 27.592957f **FLOATING
C328 AND2X2_14/B 0 19.05999f **FLOATING
C329 OAI21X1_84/C 0 12.331261f **FLOATING
C330 INVX2_59/Y 0 29.620792f **FLOATING
C331 OAI21X1_59/A 0 13.63761f **FLOATING
C332 OAI21X1_68/C 0 11.537701f **FLOATING
C333 INVX2_184/A 0 17.06685f **FLOATING
C334 NOR2X1_90/Y 0 13.312379f **FLOATING
C335 out_mines[18] 0 0.106582p **FLOATING
C336 AOI21X1_22/Y 0 10.544491f **FLOATING
C337 NOR2X1_40/Y 0 10.32396f **FLOATING
C338 INVX2_133/Y 0 8.35146f **FLOATING
C339 BUFX2_1/Y 0 25.937529f **FLOATING
C340 out_mines[19] 0 98.34232f **FLOATING
C341 out_display_done 0 23.03547f **FLOATING
C342 NOR2X1_101/Y 0 14.448361f **FLOATING
C343 INVX2_124/Y 0 8.93118f **FLOATING
C344 INVX2_23/Y 0 83.89878f **FLOATING
C345 NAND3X1_46/B 0 10.468439f **FLOATING
C346 out_temp_data_in[3] 0 0.146224p **FLOATING
C347 OAI22X1_87/B 0 36.9134f **FLOATING
C348 BUFX2_3/Y 0 71.82505f **FLOATING
C349 OAI22X1_2/Y 0 10.163819f **FLOATING
C350 OAI22X1_84/Y 0 9.407041f **FLOATING
C351 OAI22X1_86/Y 0 11.47194f **FLOATING
C352 out_mines[23] 0 0.106086p **FLOATING
C353 out_temp_data_in[1] 0 0.13572p **FLOATING
C354 out_state_main[1] 0 32.35193f **FLOATING
C355 AND2X2_6/Y 0 17.585793f **FLOATING
C356 OAI22X1_83/Y 0 9.844021f **FLOATING
C357 OAI22X1_88/D 0 28.511255f **FLOATING
C358 OAI22X1_87/D 0 33.429634f **FLOATING
C359 OAI22X1_3/D 0 19.6473f **FLOATING
C360 OAI21X1_1/B 0 0.127745p **FLOATING
C361 OAI21X1_153/Y 0 9.80076f **FLOATING
C362 INVX2_9/Y 0 15.031772f **FLOATING
C363 INVX2_84/Y 0 13.349939f **FLOATING
C364 OAI22X1_79/Y 0 13.03488f **FLOATING
C365 AOI21X1_17/A 0 14.655779f **FLOATING
C366 INVX2_8/Y 0 18.094873f **FLOATING
C367 INVX2_28/Y 0 13.564679f **FLOATING
C368 OAI22X1_2/D 0 16.298101f **FLOATING
C369 AOI22X1_78/Y 0 9.233459f **FLOATING
C370 out_temp_cleared[0] 0 12.00843f **FLOATING
C371 OAI22X1_25/Y 0 10.308779f **FLOATING
C372 OAI21X1_80/B 0 9.824401f **FLOATING
C373 INVX2_108/Y 0 15.888721f **FLOATING
C374 INVX2_123/Y 0 27.217796f **FLOATING
C375 INVX2_126/Y 0 8.261461f **FLOATING
C376 out_gameover 0 27.426567f **FLOATING
C377 NOR2X1_107/Y 0 36.768436f **FLOATING
C378 OAI22X1_39/Y 0 9.216239f **FLOATING
C379 OAI22X1_35/Y 0 10.388282f **FLOATING
C380 OAI22X1_82/Y 0 10.0686f **FLOATING
C381 INVX2_36/A 0 21.519688f **FLOATING
C382 OR2X1_10/B 0 19.986992f **FLOATING
C383 AOI21X1_23/C 0 10.49664f **FLOATING
C384 OAI21X1_110/Y 0 12.42834f **FLOATING
C385 OAI21X1_111/Y 0 12.428341f **FLOATING
C386 OAI22X1_24/Y 0 14.437561f **FLOATING
C387 INVX2_87/A 0 12.682769f **FLOATING
C388 AOI21X1_18/Y 0 11.687789f **FLOATING
C389 OAI22X1_62/Y 0 8.933039f **FLOATING
C390 AOI21X1_17/Y 0 11.64765f **FLOATING
C391 INVX2_42/Y 0 14.667121f **FLOATING
C392 OAI21X1_138/Y 0 11.14386f **FLOATING
C393 AOI21X1_26/A 0 9.97116f **FLOATING
C394 OAI22X1_34/C 0 11.5116f **FLOATING
C395 OAI22X1_61/Y 0 9.14856f **FLOATING
C396 OAI21X1_137/Y 0 11.07771f **FLOATING
C397 AOI22X1_0/Y 0 11.0649f **FLOATING
C398 NOR2X1_114/Y 0 27.02155f **FLOATING
C399 AOI22X1_70/Y 0 9.234301f **FLOATING
C400 OR2X1_7/Y 0 14.21052f **FLOATING
C401 OAI21X1_60/Y 0 11.11179f **FLOATING
C402 XOR2X1_18/Y 0 13.58874f **FLOATING
C403 out_place_done 0 18.392609f **FLOATING
C404 XNOR2X1_25/A 0 13.36071f **FLOATING
C405 OAI22X1_64/D 0 43.06368f **FLOATING
C406 AOI21X1_8/B 0 19.001698f **FLOATING
C407 OAI22X1_59/Y 0 10.917601f **FLOATING
C408 INVX2_34/A 0 16.978352f **FLOATING
C409 AOI21X1_13/B 0 14.213281f **FLOATING
C410 INVX2_48/A 0 25.600258f **FLOATING
C411 OAI22X1_60/Y 0 10.968959f **FLOATING
C412 INVX2_185/A 0 10.776541f **FLOATING
C413 INVX2_0/A 0 19.809149f **FLOATING
C414 AOI21X1_9/A 0 16.2876f **FLOATING
C415 INVX2_255/Y 0 0.125624p **FLOATING
C416 OR2X1_13/Y 0 16.0077f **FLOATING
C417 OR2X1_13/A 0 10.81875f **FLOATING
C418 XNOR2X1_27/A 0 12.776371f **FLOATING
C419 INVX2_46/A 0 8.99013f **FLOATING
C420 AOI21X1_13/Y 0 9.72213f **FLOATING
C421 HAX1_0/B 0 13.12728f **FLOATING
C422 AOI22X1_62/Y 0 13.114621f **FLOATING
C423 INVX2_49/A 0 21.43566f **FLOATING
C424 INVX2_51/A 0 23.99007f **FLOATING
C425 XOR2X1_25/Y 0 15.247231f **FLOATING
C426 INVX2_50/Y 0 18.22584f **FLOATING
C427 AOI22X1_64/Y 0 9.385019f **FLOATING
C428 OR2X1_11/Y 0 14.409842f **FLOATING
C429 XNOR2X1_28/A 0 12.733109f **FLOATING
C430 XOR2X1_26/Y 0 14.567881f **FLOATING
C431 XOR2X1_22/Y 0 15.496561f **FLOATING
C432 OAI21X1_0/C 0 14.99223f **FLOATING
C433 OR2X1_9/Y 0 14.15127f **FLOATING
C434 OR2X1_8/Y 0 9.39612f **FLOATING
C435 XNOR2X1_21/Y 0 16.37181f **FLOATING
C436 XNOR2X1_28/B 0 9.178679f **FLOATING
C437 XOR2X1_3/Y 0 31.377092f **FLOATING
C438 XOR2X1_11/Y 0 20.59986f **FLOATING
C439 OAI22X1_68/Y 0 11.078699f **FLOATING
C440 INVX2_190/A 0 8.5323f **FLOATING
C441 OAI21X1_21/Y 0 12.415561f **FLOATING
C442 OAI22X1_67/Y 0 9.930779f **FLOATING
C443 out_temp_mine_cnt[3] 0 28.632122f **FLOATING
C444 OAI21X1_3/C 0 17.332441f **FLOATING
C445 OAI22X1_47/Y 0 16.637878f **FLOATING
C446 HAX1_4/B 0 13.220099f **FLOATING
C447 HAX1_3/YS 0 10.997251f **FLOATING
C448 out_temp_mine_cnt[4] 0 20.50488f **FLOATING
C449 OAI22X1_71/Y 0 11.147639f **FLOATING
C450 HAX1_3/B 0 11.586299f **FLOATING
C451 XOR2X1_1/Y 0 9.001141f **FLOATING
C452 AND2X2_9/Y 0 10.754701f **FLOATING
C453 out_global_score[26] 0 21.545908f **FLOATING
C454 BUFX2_8/Y 0 40.152676f **FLOATING
C455 OAI21X1_23/Y 0 11.74776f **FLOATING
C456 OAI21X1_3/Y 0 11.72886f **FLOATING
C457 AOI22X1_72/Y 0 14.99682f **FLOATING
C458 AOI21X1_16/A 0 9.490199f **FLOATING
C459 OAI22X1_69/Y 0 12.31092f **FLOATING
C460 OAI21X1_44/A 0 41.168922f **FLOATING
C461 OAI21X1_33/Y 0 13.064102f **FLOATING
C462 OAI21X1_47/Y 0 10.99626f **FLOATING
C463 INVX2_229/A 0 10.02318f **FLOATING
C464 OAI22X1_70/Y 0 12.992341f **FLOATING
C465 INVX2_231/Y 0 14.712899f **FLOATING
C466 INVX2_231/A 0 10.17846f **FLOATING
C467 OAI21X1_35/Y 0 10.553221f **FLOATING
C468 OAI22X1_42/Y 0 11.597881f **FLOATING
C469 BUFX2_18/Y 0 53.660206f **FLOATING
C470 NAND3X1_8/Y 0 34.70743f **FLOATING
C471 BUFX2_19/A 0 42.81912f **FLOATING
C472 HAX1_6/B 0 12.29184f **FLOATING
C473 INVX2_193/Y 0 11.327579f **FLOATING
C474 AND2X2_13/Y 0 11.47875f **FLOATING
C475 INVX2_240/Y 0 11.620621f **FLOATING
C476 OAI21X1_7/C 0 9.129241f **FLOATING
C477 out_global_score[24] 0 19.010609f **FLOATING
C478 out_global_score[23] 0 14.925629f **FLOATING
C479 INVX2_29/Y 0 8.49102f **FLOATING
C480 OAI21X1_51/Y 0 10.22112f **FLOATING
C481 INVX2_181/Y 0 11.697959f **FLOATING
C482 OAI21X1_4/Y 0 14.724299f **FLOATING
C483 OAI22X1_75/Y 0 9.76344f **FLOATING
C484 INVX2_243/A 0 8.59506f **FLOATING
C485 OR2X1_12/A 0 34.695858f **FLOATING
C486 OAI22X1_73/Y 0 10.11708f **FLOATING
C487 OAI21X1_7/Y 0 13.0707f **FLOATING
C488 OAI22X1_52/Y 0 9.32718f **FLOATING
C489 OAI21X1_146/Y 0 10.38066f **FLOATING
C490 OR2X1_12/B 0 26.53467f **FLOATING
C491 OAI22X1_76/Y 0 9.95598f **FLOATING
C492 HAX1_37/YS 0 14.624732f **FLOATING
C493 INVX2_226/A 0 11.871121f **FLOATING
C494 OAI21X1_19/Y 0 13.875602f **FLOATING
C495 out_global_score[21] 0 18.654211f **FLOATING
C496 OAI21X1_9/Y 0 13.75686f **FLOATING
C497 NOR2X1_66/Y 0 19.478281f **FLOATING
C498 FAX1_11/C 0 17.01567f **FLOATING
C499 INVX2_196/A 0 9.15792f **FLOATING
C500 OAI21X1_17/Y 0 13.41462f **FLOATING
C501 out_global_score[3] 0 19.25829f **FLOATING
C502 NOR2X1_67/Y 0 47.027435f **FLOATING
C503 OAI21X1_11/Y 0 12.46314f **FLOATING
C504 FAX1_13/B 0 17.41263f **FLOATING
C505 INVX2_196/Y 0 8.787181f **FLOATING
C506 INVX2_213/Y 0 10.923481f **FLOATING
C507 out_global_score[4] 0 18.28863f **FLOATING
C508 OAI21X1_53/Y 0 13.31982f **FLOATING
C509 FAX1_13/C 0 13.759529f **FLOATING
C510 FAX1_11/B 0 15.625471f **FLOATING
C511 out_global_score[20] 0 19.374329f **FLOATING
C512 out_temp_index[2] 0 15.96975f **FLOATING
C513 FAX1_11/A 0 17.49699f **FLOATING
C514 out_temp_index[4] 0 16.660769f **FLOATING
C515 OAI21X1_5/Y 0 13.44384f **FLOATING
C516 FAX1_12/B 0 16.374903f **FLOATING
C517 INVX2_197/A 0 8.43066f **FLOATING
C518 out_temp_index[3] 0 16.528948f **FLOATING
C519 HAX1_31/A 0 12.528239f **FLOATING
C520 FAX1_5/B 0 17.696913f **FLOATING
C521 out_global_score[19] 0 18.908491f **FLOATING
C522 HAX1_28/B 0 12.6729f **FLOATING
C523 XNOR2X1_1/A 0 21.820591f **FLOATING
C524 MUX2X1_32/B 0 9.09192f **FLOATING
C525 out_global_score[2] 0 14.925631f **FLOATING
C526 out_global_score[6] 0 15.923189f **FLOATING
C527 FAX1_4/C 0 14.529271f **FLOATING
C528 FAX1_14/B 0 16.23321f **FLOATING
C529 HAX1_24/YS 0 10.290271f **FLOATING
C530 XNOR2X1_1/Y 0 9.17841f **FLOATING
C531 NOR2X1_8/Y 0 12.90882f **FLOATING
C532 FAX1_10/B 0 17.150372f **FLOATING
C533 FAX1_5/C 0 14.10627f **FLOATING
C534 INVX2_214/Y 0 11.199121f **FLOATING
C535 NOR2X1_0/Y 0 12.731702f **FLOATING
C536 NOR2X1_0/A 0 18.36129f **FLOATING
C537 HAX1_30/A 0 14.21646f **FLOATING
C538 FAX1_8/A 0 17.07561f **FLOATING
C539 FAX1_7/B 0 16.69182f **FLOATING
C540 OR2X1_1/Y 0 38.928356f **FLOATING
C541 FAX1_8/C 0 15.10707f **FLOATING
C542 FAX1_16/C 0 15.98928f **FLOATING
C543 FAX1_7/A 0 15.40053f **FLOATING
C544 XOR2X1_5/A 0 14.249642f **FLOATING
C545 INVX2_198/A 0 9.898381f **FLOATING
C546 FAX1_3/YS 0 18.277647f **FLOATING
C547 FAX1_7/C 0 13.13309f **FLOATING
C548 XOR2X1_8/A 0 13.15248f **FLOATING
C549 FAX1_2/A 0 19.28292f **FLOATING
C550 HAX1_49/YS 0 10.87473f **FLOATING
C551 out_global_score[16] 0 19.38837f **FLOATING
C552 out_global_score[12] 0 19.959211f **FLOATING
C553 HAX1_19/YS 0 10.60365f **FLOATING
C554 HAX1_49/A 0 16.646881f **FLOATING
C555 XNOR2X1_3/Y 0 10.544669f **FLOATING
C556 FAX1_1/C 0 14.301269f **FLOATING
C557 XOR2X1_9/Y 0 19.028881f **FLOATING
C558 OR2X1_5/Y 0 36.77742f **FLOATING
C559 NOR2X1_7/Y 0 33.256924f **FLOATING
C560 NOR2X1_6/Y 0 15.374041f **FLOATING
C561 INVX2_208/A 0 8.13648f **FLOATING
C562 XNOR2X1_5/A 0 20.37639f **FLOATING
C563 NOR2X1_4/Y 0 14.332621f **FLOATING
C564 MUX2X1_7/Y 0 10.222141f **FLOATING
C565 NOR2X1_5/Y 0 13.016101f **FLOATING
C566 HAX1_16/B 0 14.803139f **FLOATING
C567 HAX1_47/B 0 15.01608f **FLOATING
C568 HAX1_15/B 0 13.69104f **FLOATING
C569 HAX1_43/B 0 12.058951f **FLOATING
C570 MUX2X1_15/Y 0 13.7775f **FLOATING
C571 MUX2X1_0/B 0 16.133432f **FLOATING
C572 INVX2_202/Y 0 9.691381f **FLOATING
C573 out_global_score[10] 0 19.37541f **FLOATING
C574 out_global_score[9] 0 15.378511f **FLOATING
C575 OR2X1_1/B 0 8.6436f **FLOATING
C576 HAX1_42/B 0 13.02174f **FLOATING
C577 MUX2X1_0/A 0 10.122509f **FLOATING
C578 MUX2X1_20/Y 0 8.98788f **FLOATING
C579 MUX2X1_10/Y 0 8.99418f **FLOATING
C580 HAX1_45/B 0 12.012541f **FLOATING
C581 HAX1_45/A 0 15.909598f **FLOATING
C582 OR2X1_3/Y 0 38.47968f **FLOATING
C583 HAX1_41/B 0 12.01254f **FLOATING
C584 HAX1_39/B 0 12.01704f **FLOATING
C585 MUX2X1_16/Y 0 13.38978f **FLOATING
C586 out_display 0 26.636568f **FLOATING
C587 INVX2_121/A 0 15.04806f **FLOATING
C588 OAI21X1_156/Y 0 11.563862f **FLOATING
C589 NAND3X1_49/Y 0 9.88605f **FLOATING
C590 INVX2_120/A 0 27.268408f **FLOATING
C591 INVX2_117/A 0 24.610292f **FLOATING
C592 INVX2_128/Y 0 10.88208f **FLOATING
C593 INVX2_128/A 0 8.64501f **FLOATING
C594 NOR2X1_125/Y 0 29.079119f **FLOATING
C595 NOR2X1_124/Y 0 23.341913f **FLOATING
C596 INVX2_119/Y 0 15.640198f **FLOATING
C597 NAND3X1_52/Y 0 10.699651f **FLOATING
C598 INVX2_119/A 0 35.698727f **FLOATING
C599 INVX2_125/Y 0 24.43611f **FLOATING
C600 out_state_main[2] 0 39.98532f **FLOATING
C601 AND2X2_18/Y 0 9.13881f **FLOATING
C602 NOR2X1_122/Y 0 8.142241f **FLOATING
C603 INVX2_126/A 0 9.52818f **FLOATING
C604 out_state_main[3] 0 39.90015f **FLOATING
C605 out_state_main[0] 0 30.153156f **FLOATING
C606 NOR2X1_117/Y 0 8.436241f **FLOATING
C607 INVX2_123/A 0 11.278709f **FLOATING
C608 NOR2X1_120/Y 0 12.135181f **FLOATING
C609 INVX2_116/Y 0 18.44869f **FLOATING
C610 AOI21X1_26/C 0 9.99042f **FLOATING
C611 INVX2_118/Y 0 12.861361f **FLOATING
C612 INVX2_133/A 0 9.79305f **FLOATING
C613 OR2X1_15/A 0 17.74113f **FLOATING
C614 OR2X1_15/Y 0 11.629771f **FLOATING
C615 INVX2_122/A 0 13.224091f **FLOATING
C616 in_data_in 0 12.45708f **FLOATING
C617 AND2X2_19/B 0 16.958218f **FLOATING
C618 out_load 0 22.16591f **FLOATING
C619 AND2X2_19/Y 0 9.25725f **FLOATING
C620 AOI21X1_24/Y 0 15.23352f **FLOATING
C621 AOI21X1_25/Y 0 11.15469f **FLOATING
C622 OR2X1_16/Y 0 14.181481f **FLOATING
C623 XOR2X1_2/Y 0 8.8935f **FLOATING
C624 out_global_score[31] 0 17.498398f **FLOATING
C625 HAX1_0/YS 0 12.64647f **FLOATING
C626 INVX2_187/Y 0 11.303821f **FLOATING
C627 AND2X2_14/Y 0 8.366791f **FLOATING
C628 INVX2_186/A 0 8.11314f **FLOATING
C629 INVX2_191/A 0 10.845061f **FLOATING
C630 out_global_score[25] 0 19.825771f **FLOATING
C631 INVX2_187/A 0 9.64086f **FLOATING
C632 HAX1_1/B 0 12.083099f **FLOATING
C633 out_start 0 56.282654f **FLOATING
C634 INVX2_132/Y 0 11.862961f **FLOATING
C635 OAI21X1_59/Y 0 11.70111f **FLOATING
C636 INVX2_184/Y 0 15.56616f **FLOATING
C637 out_alu_done 0 28.94754f **FLOATING
C638 OAI22X1_21/Y 0 10.576621f **FLOATING
C639 out_temp_decoded[7] 0 18.685411f **FLOATING
C640 OAI21X1_71/C 0 11.346449f **FLOATING
C641 INVX2_15/Y 0 29.158005f **FLOATING
C642 OAI22X1_1/B 0 18.421381f **FLOATING
C643 NOR2X1_85/Y 0 15.08328f **FLOATING
C644 OAI21X1_58/Y 0 15.27528f **FLOATING
C645 INVX2_111/Y 0 12.175802f **FLOATING
C646 OAI21X1_57/Y 0 11.27628f **FLOATING
C647 OAI22X1_28/Y 0 10.576619f **FLOATING
C648 OAI22X1_27/Y 0 10.77798f **FLOATING
C649 INVX2_218/Y 0 9.44658f **FLOATING
C650 OAI21X1_66/C 0 9.4605f **FLOATING
C651 out_temp_decoded[8] 0 14.78124f **FLOATING
C652 OAI22X1_19/Y 0 11.18082f **FLOATING
C653 OAI22X1_3/Y 0 9.178319f **FLOATING
C654 NOR2X1_82/B 0 20.96001f **FLOATING
C655 NOR2X1_83/B 0 8.674289f **FLOATING
C656 NOR2X1_87/A 0 8.99709f **FLOATING
C657 INVX2_71/Y 0 25.018682f **FLOATING
C658 INVX2_103/Y 0 9.069539f **FLOATING
C659 INVX2_104/Y 0 21.14664f **FLOATING
C660 INVX2_73/Y 0 6.67872f **FLOATING
C661 NOR2X1_90/A 0 8.69106f **FLOATING
C662 NOR2X1_69/Y 0 9.79398f **FLOATING
C663 HAX1_2/YS 0 10.763371f **FLOATING
C664 INVX2_190/Y 0 10.401779f **FLOATING
C665 INVX2_188/A 0 8.2485f **FLOATING
C666 INVX2_188/Y 0 11.92524f **FLOATING
C667 HAX1_2/B 0 15.615301f **FLOATING
C668 INVX2_192/A 0 13.326211f **FLOATING
C669 INVX2_195/A 0 13.471979f **FLOATING
C670 HAX1_5/B 0 19.870382f **FLOATING
C671 INVX2_197/Y 0 8.604779f **FLOATING
C672 INVX2_200/Y 0 11.21502f **FLOATING
C673 HAX1_9/B 0 12.59868f **FLOATING
C674 out_global_score[22] 0 15.092158f **FLOATING
C675 INVX2_193/A 0 10.625701f **FLOATING
C676 INVX2_194/A 0 8.01198f **FLOATING
C677 XNOR2X1_24/Y 0 9.36609f **FLOATING
C678 INVX2_0/Y 0 8.7408f **FLOATING
C679 AND2X2_8/A 0 26.99898f **FLOATING
C680 AND2X2_8/B 0 12.835709f **FLOATING
C681 OAI22X1_3/B 0 15.89616f **FLOATING
C682 INVX2_10/Y 0 32.976383f **FLOATING
C683 OAI21X1_84/Y 0 11.208481f **FLOATING
C684 NOR2X1_83/A 0 13.685069f **FLOATING
C685 INVX2_217/A 0 44.174362f **FLOATING
C686 BUFX2_9/A 0 31.196962f **FLOATING
C687 out_win 0 18.09807f **FLOATING
C688 OAI21X1_65/Y 0 14.6436f **FLOATING
C689 INVX2_83/Y 0 24.019318f **FLOATING
C690 INVX2_84/A 0 12.580651f **FLOATING
C691 OAI22X1_0/Y 0 16.567741f **FLOATING
C692 NOR2X1_87/Y 0 13.83664f **FLOATING
C693 BUFX2_7/A 0 8.403271f **FLOATING
C694 NOR2X1_82/Y 0 7.946701f **FLOATING
C695 NOR2X1_82/A 0 10.414891f **FLOATING
C696 NOR2X1_88/Y 0 10.44264f **FLOATING
C697 INVX2_73/A 0 16.11396f **FLOATING
C698 OAI21X1_67/C 0 7.269899f **FLOATING
C699 BUFX2_13/Y 0 0.169197p **FLOATING
C700 OAI21X1_94/C 0 13.051619f **FLOATING
C701 BUFX2_22/Y 0 81.04724f **FLOATING
C702 NOR2X1_58/Y 0 9.33456f **FLOATING
C703 OAI21X1_85/C 0 13.16004f **FLOATING
C704 OAI21X1_75/C 0 12.986851f **FLOATING
C705 AOI21X1_3/A 0 44.600204f **FLOATING
C706 OAI21X1_85/Y 0 11.144521f **FLOATING
C707 OAI21X1_80/C 0 10.08849f **FLOATING
C708 BUFX2_5/A 0 6.56301f **FLOATING
C709 out_n_nearby[0] 0 14.325271f **FLOATING
C710 HAX1_35/B 0 16.81674f **FLOATING
C711 XNOR2X1_22/Y 0 10.629809f **FLOATING
C712 HAX1_36/B 0 11.5872f **FLOATING
C713 out_temp_mine_cnt[1] 0 27.42366f **FLOATING
C714 out_temp_mine_cnt[0] 0 25.670462f **FLOATING
C715 OAI21X1_62/Y 0 10.373401f **FLOATING
C716 OAI21X1_62/B 0 14.732221f **FLOATING
C717 OAI22X1_2/B 0 17.602621f **FLOATING
C718 AOI21X1_6/C 0 10.131181f **FLOATING
C719 INVX2_6/Y 0 20.664122f **FLOATING
C720 OAI21X1_70/C 0 10.454161f **FLOATING
C721 out_temp_decoded[3] 0 15.563551f **FLOATING
C722 INVX2_81/Y 0 31.37677f **FLOATING
C723 NOR2X1_38/Y 0 8.336221f **FLOATING
C724 NOR2X1_73/A 0 27.733288f **FLOATING
C725 NOR2X1_78/B 0 9.66609f **FLOATING
C726 OAI22X1_16/Y 0 10.60566f **FLOATING
C727 NOR2X1_55/Y 0 7.49442f **FLOATING
C728 OAI21X1_87/Y 0 11.144522f **FLOATING
C729 OAI21X1_86/C 0 11.54844f **FLOATING
C730 OAI21X1_86/Y 0 11.144521f **FLOATING
C731 NOR2X1_74/Y 0 12.21078f **FLOATING
C732 NOR2X1_40/B 0 26.35265f **FLOATING
C733 out_mines[4] 0 0.1147p **FLOATING
C734 out_temp_cleared[5] 0 16.26141f **FLOATING
C735 INVX2_86/A 0 18.88695f **FLOATING
C736 in_clka 0 15.67584f **FLOATING
C737 NOR2X1_72/A 0 7.138051f **FLOATING
C738 XNOR2X1_26/A 0 10.94439f **FLOATING
C739 OAI21X1_37/Y 0 11.29992f **FLOATING
C740 AND2X2_12/Y 0 10.748251f **FLOATING
C741 HAX1_10/B 0 13.44222f **FLOATING
C742 INVX2_215/A 0 7.963619f **FLOATING
C743 HAX1_29/YS 0 11.70525f **FLOATING
C744 INVX2_213/A 0 8.11314f **FLOATING
C745 HAX1_13/B 0 14.603101f **FLOATING
C746 out_global_score[1] 0 20.96421f **FLOATING
C747 HAX1_27/YS 0 12.57357f **FLOATING
C748 INVX2_212/A 0 8.2485f **FLOATING
C749 HAX1_26/YS 0 11.595571f **FLOATING
C750 BUFX2_8/A 0 7.72872f **FLOATING
C751 OAI21X1_47/C 0 8.630341f **FLOATING
C752 INVX2_79/Y 0 27.230436f **FLOATING
C753 AND2X2_15/Y 0 21.525446f **FLOATING
C754 NOR2X1_77/Y 0 9.228871f **FLOATING
C755 NOR2X1_77/A 0 18.677769f **FLOATING
C756 out_temp_decoded[4] 0 25.85217f **FLOATING
C757 OR2X1_14/A 0 19.301313f **FLOATING
C758 NOR2X1_75/Y 0 8.208841f **FLOATING
C759 XOR2X1_20/Y 0 22.013008f **FLOATING
C760 XOR2X1_23/Y 0 12.69852f **FLOATING
C761 INVX2_88/A 0 10.30908f **FLOATING
C762 OR2X1_14/Y 0 20.92968f **FLOATING
C763 OR2X1_14/B 0 15.28494f **FLOATING
C764 XNOR2X1_25/B 0 9.520199f **FLOATING
C765 XOR2X1_24/Y 0 9.3543f **FLOATING
C766 XOR2X1_23/B 0 11.99934f **FLOATING
C767 XOR2X1_24/A 0 17.58858f **FLOATING
C768 NOR2X1_104/B 0 14.73871f **FLOATING
C769 NOR2X1_96/Y 0 13.1091f **FLOATING
C770 NAND2X1_89/Y 0 9.10434f **FLOATING
C771 INVX2_30/Y 0 29.993118f **FLOATING
C772 BUFX2_15/Y 0 0.178619p **FLOATING
C773 OAI22X1_8/Y 0 13.528379f **FLOATING
C774 NOR2X1_99/Y 0 15.225301f **FLOATING
C775 NOR2X1_86/A 0 26.53953f **FLOATING
C776 NOR2X1_75/B 0 24.836027f **FLOATING
C777 INVX2_67/Y 0 27.189238f **FLOATING
C778 out_mines[12] 0 0.1232p **FLOATING
C779 NOR2X1_93/Y 0 10.9344f **FLOATING
C780 OAI21X1_96/C 0 12.439139f **FLOATING
C781 NAND2X1_88/Y 0 9.68214f **FLOATING
C782 NOR2X1_76/Y 0 7.96254f **FLOATING
C783 INVX2_62/A 0 13.718147f **FLOATING
C784 out_temp_data_in[0] 0 0.149337p **FLOATING
C785 NOR2X1_97/B 0 8.674289f **FLOATING
C786 INVX2_14/Y 0 46.002567f **FLOATING
C787 INVX2_94/Y 0 10.07031f **FLOATING
C788 NAND3X1_44/B 0 9.011339f **FLOATING
C789 INVX2_217/Y 0 42.359486f **FLOATING
C790 INVX2_31/Y 0 47.440647f **FLOATING
C791 INVX2_13/Y 0 17.524439f **FLOATING
C792 out_mines[13] 0 0.11289p **FLOATING
C793 NAND3X1_39/B 0 10.610161f **FLOATING
C794 NOR2X1_91/B 0 9.700891f **FLOATING
C795 OAI21X1_97/C 0 13.51944f **FLOATING
C796 BUFX2_21/Y 0 58.74002f **FLOATING
C797 NOR2X1_50/Y 0 7.56102f **FLOATING
C798 OAI21X1_100/Y 0 16.2435f **FLOATING
C799 out_mines[16] 0 86.42235f **FLOATING
C800 OAI21X1_98/Y 0 10.65756f **FLOATING
C801 OAI21X1_98/C 0 9.68574f **FLOATING
C802 NOR2X1_53/Y 0 7.56102f **FLOATING
C803 NOR2X1_57/B 0 44.99598f **FLOATING
C804 NOR2X1_55/A 0 40.42625f **FLOATING
C805 NOR2X1_52/Y 0 7.56102f **FLOATING
C806 NOR2X1_47/B 0 26.472397f **FLOATING
C807 XNOR2X1_27/B 0 9.97902f **FLOATING
C808 OAI21X1_39/Y 0 11.144522f **FLOATING
C809 INVX2_226/Y 0 10.36056f **FLOATING
C810 OAI21X1_39/C 0 8.146441f **FLOATING
C811 INVX2_232/Y 0 9.477601f **FLOATING
C812 INVX2_232/A 0 9.772019f **FLOATING
C813 INVX2_45/Y 0 8.073541f **FLOATING
C814 XNOR2X1_26/B 0 9.831199f **FLOATING
C815 OAI21X1_108/Y 0 13.2681f **FLOATING
C816 INVX2_45/A 0 34.23672f **FLOATING
C817 INVX2_44/A 0 27.710114f **FLOATING
C818 NOR2X1_108/Y 0 8.7906f **FLOATING
C819 INVX2_32/A 0 27.421886f **FLOATING
C820 OAI22X1_37/D 0 9.61098f **FLOATING
C821 OAI21X1_114/Y 0 10.34646f **FLOATING
C822 AND2X2_16/Y 0 20.265808f **FLOATING
C823 XOR2X1_25/B 0 40.802185f **FLOATING
C824 OAI21X1_41/C 0 9.100141f **FLOATING
C825 OAI21X1_48/B 0 22.992722f **FLOATING
C826 HAX1_27/B 0 12.639899f **FLOATING
C827 HAX1_26/B 0 12.490501f **FLOATING
C828 HAX1_28/YS 0 10.16799f **FLOATING
C829 HAX1_13/YS 0 9.87783f **FLOATING
C830 HAX1_14/B 0 14.225579f **FLOATING
C831 INVX2_114/Y 0 9.281881f **FLOATING
C832 INVX2_216/A 0 9.14826f **FLOATING
C833 INVX2_214/A 0 8.261459f **FLOATING
C834 HAX1_24/B 0 13.686299f **FLOATING
C835 HAX1_25/B 0 14.1897f **FLOATING
C836 OAI21X1_49/C 0 8.08944f **FLOATING
C837 INVX2_237/Y 0 10.19298f **FLOATING
C838 OAI21X1_41/Y 0 14.410558f **FLOATING
C839 INVX2_222/Y 0 8.94756f **FLOATING
C840 NOR2X1_64/Y 0 13.273801f **FLOATING
C841 NOR2X1_65/Y 0 8.208841f **FLOATING
C842 OAI21X1_31/Y 0 10.490218f **FLOATING
C843 OAI21X1_9/B 0 0.148881p **FLOATING
C844 OAI21X1_29/Y 0 11.82246f **FLOATING
C845 INVX2_47/Y 0 7.497841f **FLOATING
C846 OAI22X1_40/D 0 10.084379f **FLOATING
C847 OAI21X1_116/Y 0 12.29982f **FLOATING
C848 AOI22X1_60/Y 0 9.50952f **FLOATING
C849 INVX2_242/Y 0 14.401502f **FLOATING
C850 INVX2_235/Y 0 10.400579f **FLOATING
C851 OAI21X1_25/Y 0 12.371161f **FLOATING
C852 NOR2X1_66/B 0 0.11511p **FLOATING
C853 INVX2_235/A 0 9.09366f **FLOATING
C854 NOR2X1_64/A 0 11.273069f **FLOATING
C855 INVX2_211/A 0 7.610041f **FLOATING
C856 HAX1_25/YS 0 10.322251f **FLOATING
C857 HAX1_16/YS 0 9.72225f **FLOATING
C858 INVX2_203/Y 0 10.36098f **FLOATING
C859 INVX2_210/A 0 8.2485f **FLOATING
C860 INVX2_202/A 0 10.947899f **FLOATING
C861 INVX2_206/Y 0 11.303821f **FLOATING
C862 INVX2_205/Y 0 12.10038f **FLOATING
C863 INVX2_205/A 0 8.11314f **FLOATING
C864 HAX1_22/B 0 15.898261f **FLOATING
C865 HAX1_23/YS 0 9.845429f **FLOATING
C866 INVX2_209/A 0 7.89246f **FLOATING
C867 HAX1_19/B 0 15.87642f **FLOATING
C868 HAX1_21/YS 0 11.173591f **FLOATING
C869 HAX1_21/B 0 12.086699f **FLOATING
C870 INVX2_206/A 0 8.11314f **FLOATING
C871 HAX1_22/YS 0 10.322251f **FLOATING
C872 OAI21X1_56/C 0 8.31858f **FLOATING
C873 HAX1_48/B 0 11.73816f **FLOATING
C874 OR2X1_0/B 0 9.88308f **FLOATING
C875 HAX1_48/A 0 14.45508f **FLOATING
C876 NAND3X1_9/A 0 27.99871f **FLOATING
C877 OAI21X1_56/Y 0 10.85157f **FLOATING
C878 NAND3X1_7/Y 0 48.14422f **FLOATING
C879 OAI21X1_30/B 0 16.18188f **FLOATING
C880 NOR2X1_62/Y 0 17.314259f **FLOATING
C881 OR2X1_12/Y 0 8.85576f **FLOATING
C882 OAI21X1_32/B 0 21.167099f **FLOATING
C883 INVX2_230/A 0 8.973359f **FLOATING
C884 INVX2_236/Y 0 14.197619f **FLOATING
C885 OAI22X1_36/C 0 10.08918f **FLOATING
C886 AOI21X1_9/C 0 9.47925f **FLOATING
C887 out_temp_data_in[2] 0 0.150713p **FLOATING
C888 OAI22X1_10/Y 0 10.04838f **FLOATING
C889 INVX2_95/Y 0 14.91882f **FLOATING
C890 INVX2_24/Y 0 12.69576f **FLOATING
C891 AOI22X1_55/Y 0 8.731501f **FLOATING
C892 INVX2_42/A 0 8.577089f **FLOATING
C893 INVX2_32/Y 0 53.619453f **FLOATING
C894 AOI21X1_8/C 0 15.779877f **FLOATING
C895 INVX2_41/A 0 21.70554f **FLOATING
C896 BUFX2_14/Y 0 0.168468p **FLOATING
C897 INVX2_64/Y 0 20.362976f **FLOATING
C898 BUFX2_23/Y 0 89.22652f **FLOATING
C899 AOI22X1_71/Y 0 10.21704f **FLOATING
C900 AOI22X1_63/Y 0 8.901481f **FLOATING
C901 BUFX2_19/Y 0 57.403248f **FLOATING
C902 INVX2_180/Y 0 10.964642f **FLOATING
C903 OAI21X1_54/Y 0 12.13344f **FLOATING
C904 OAI21X1_8/B 0 19.56918f **FLOATING
C905 OAI21X1_27/Y 0 13.912801f **FLOATING
C906 OAI21X1_8/Y 0 9.398459f **FLOATING
C907 INVX2_220/A 0 13.73982f **FLOATING
C908 INVX2_234/A 0 12.051419f **FLOATING
C909 OAI21X1_6/Y 0 22.47954f **FLOATING
C910 INVX2_239/A 0 11.244961f **FLOATING
C911 OAI21X1_15/C 0 8.146441f **FLOATING
C912 AOI22X1_61/Y 0 11.631241f **FLOATING
C913 AOI22X1_69/B 0 19.608599f **FLOATING
C914 AOI22X1_59/Y 0 9.617221f **FLOATING
C915 AND2X2_16/B 0 8.878711f **FLOATING
C916 NOR2X1_112/Y 0 27.897177f **FLOATING
C917 INVX2_89/Y 0 14.4516f **FLOATING
C918 INVX2_54/A 0 11.362771f **FLOATING
C919 INVX2_11/Y 0 10.31658f **FLOATING
C920 OAI21X1_79/C 0 11.03145f **FLOATING
C921 NAND2X1_90/Y 0 15.49242f **FLOATING
C922 AOI21X1_7/Y 0 12.00429f **FLOATING
C923 NOR2X1_97/A 0 13.74607f **FLOATING
C924 out_mines[24] 0 60.634747f **FLOATING
C925 AOI22X1_68/Y 0 8.1408f **FLOATING
C926 NOR2X1_110/B 0 37.42078f **FLOATING
C927 OR2X1_6/A 0 80.41687f **FLOATING
C928 INVX2_20/Y 0 9.01524f **FLOATING
C929 AOI22X1_67/Y 0 10.261501f **FLOATING
C930 out_mines[6] 0 0.126525p **FLOATING
C931 out_mines[7] 0 0.126729p **FLOATING
C932 NAND2X1_63/A 0 11.138579f **FLOATING
C933 INVX2_18/Y 0 22.767437f **FLOATING
C934 AOI21X1_18/A 0 19.4949f **FLOATING
C935 INVX2_56/Y 0 12.56856f **FLOATING
C936 OAI22X1_5/Y 0 11.503139f **FLOATING
C937 INVX2_90/Y 0 7.67754f **FLOATING
C938 out_mines[5] 0 79.21423f **FLOATING
C939 OAI22X1_80/Y 0 9.09378f **FLOATING
C940 out_mines[0] 0 97.429436f **FLOATING
C941 AOI21X1_12/Y 0 12.93189f **FLOATING
C942 OAI22X1_63/Y 0 9.400501f **FLOATING
C943 OAI22X1_43/Y 0 8.43162f **FLOATING
C944 INVX2_224/Y 0 10.05258f **FLOATING
C945 INVX2_220/Y 0 15.448802f **FLOATING
C946 AOI22X1_72/A 0 10.833721f **FLOATING
C947 OAI22X1_45/Y 0 9.44892f **FLOATING
C948 INVX2_52/A 0 38.424114f **FLOATING
C949 OAI22X1_55/Y 0 11.24202f **FLOATING
C950 OAI22X1_64/Y 0 14.131619f **FLOATING
C951 NAND3X1_46/A 0 13.7931f **FLOATING
C952 OAI21X1_77/C 0 8.964451f **FLOATING
C953 INVX2_92/Y 0 8.9082f **FLOATING
C954 INVX2_53/Y 0 8.85789f **FLOATING
C955 OAI22X1_49/Y 0 9.30834f **FLOATING
C956 INVX2_53/A 0 14.027582f **FLOATING
C957 OAI22X1_51/B 0 45.1084f **FLOATING
C958 OAI22X1_48/Y 0 10.873501f **FLOATING
C959 OR2X1_0/Y 0 33.377396f **FLOATING
C960 in_incr[0] 0 4.99065f **FLOATING
C961 OR2X1_0/A 0 16.0935f **FLOATING
C962 INVX2_207/A 0 8.224979f **FLOATING
C963 HAX1_46/YS 0 8.304689f **FLOATING
C964 MUX2X1_27/Y 0 11.828699f **FLOATING
C965 MUX2X1_27/B 0 6.84966f **FLOATING
C966 HAX1_46/A 0 14.804729f **FLOATING
C967 NOR2X1_1/Y 0 14.58312f **FLOATING
C968 MUX2X1_24/Y 0 10.742339f **FLOATING
C969 XNOR2X1_2/Y 0 9.43125f **FLOATING
C970 NOR2X1_1/A 0 21.399902f **FLOATING
C971 FAX1_2/C 0 19.594889f **FLOATING
C972 FAX1_3/C 0 15.114539f **FLOATING
C973 HAX1_34/B 0 13.268641f **FLOATING
C974 NOR2X1_9/A 0 30.777721f **FLOATING
C975 FAX1_10/C 0 17.16912f **FLOATING
C976 FAX1_18/C 0 17.917528f **FLOATING
C977 NOR2X1_17/B 0 24.959547f **FLOATING
C978 FAX1_16/B 0 20.665018f **FLOATING
C979 FAX1_17/B 0 17.71875f **FLOATING
C980 OAI21X1_5/C 0 8.407441f **FLOATING
C981 OAI21X1_9/A 0 10.20798f **FLOATING
C982 HAX1_32/B 0 9.72912f **FLOATING
C983 OAI21X1_5/A 0 10.615141f **FLOATING
C984 OAI22X1_52/D 0 36.319736f **FLOATING
C985 OAI22X1_88/B 0 31.809212f **FLOATING
C986 INVX2_19/Y 0 41.212547f **FLOATING
C987 out_temp_cleared[21] 0 19.637129f **FLOATING
C988 out_mines[3] 0 0.101478p **FLOATING
C989 INVX2_37/Y 0 9.281519f **FLOATING
C990 OAI22X1_64/B 0 42.465984f **FLOATING
C991 out_mines[2] 0 0.170767p **FLOATING
C992 OAI22X1_63/D 0 32.095284f **FLOATING
C993 OAI22X1_81/Y 0 8.284681f **FLOATING
C994 OAI22X1_53/Y 0 9.974641f **FLOATING
C995 OAI22X1_85/Y 0 8.320619f **FLOATING
C996 OAI22X1_87/Y 0 12.203879f **FLOATING
C997 OAI22X1_88/Y 0 14.57268f **FLOATING
C998 OAI21X1_154/Y 0 9.07758f **FLOATING
C999 OAI22X1_77/Y 0 10.562281f **FLOATING
C1000 OAI22X1_78/Y 0 12.17526f **FLOATING
C1001 AOI21X1_17/B 0 9.466621f **FLOATING
C1002 OAI22X1_58/Y 0 11.178301f **FLOATING
C1003 OAI22X1_57/Y 0 9.15912f **FLOATING
C1004 INVX2_37/A 0 19.3776f **FLOATING
C1005 OAI22X1_76/D 0 31.111256f **FLOATING
C1006 OAI22X1_75/D 0 32.10847f **FLOATING
C1007 AOI21X1_18/B 0 10.458961f **FLOATING
C1008 AOI21X1_14/A 0 9.613801f **FLOATING
C1009 INVX2_36/Y 0 11.009881f **FLOATING
C1010 AOI22X1_75/Y 0 9.75222f **FLOATING
C1011 OAI21X1_148/Y 0 8.38662f **FLOATING
C1012 XOR2X1_28/A 0 27.392408f **FLOATING
C1013 INVX2_34/Y 0 16.894861f **FLOATING
C1014 AOI22X1_73/Y 0 10.111739f **FLOATING
C1015 OR2X1_10/Y 0 10.059091f **FLOATING
C1016 AOI21X1_13/A 0 15.796619f **FLOATING
C1017 AOI21X1_15/A 0 8.84676f **FLOATING
C1018 OAI22X1_72/Y 0 9.721921f **FLOATING
C1019 OR2X1_8/B 0 15.742561f **FLOATING
C1020 AOI21X1_15/Y 0 9.83355f **FLOATING
C1021 OAI21X1_140/Y 0 8.705819f **FLOATING
C1022 AOI21X1_15/B 0 15.58324f **FLOATING
C1023 OAI22X1_65/Y 0 9.556979f **FLOATING
C1024 OAI22X1_66/Y 0 9.579719f **FLOATING
C1025 AOI21X1_16/B 0 9.807421f **FLOATING
C1026 AOI22X1_74/Y 0 11.12862f **FLOATING
C1027 OAI21X1_145/Y 0 7.87782f **FLOATING
C1028 OAI22X1_74/Y 0 21.46935f **FLOATING
C1029 FAX1_14/C 0 18.896519f **FLOATING
C1030 FAX1_15/C 0 15.150631f **FLOATING
C1031 FAX1_15/B 0 15.446913f **FLOATING
C1032 FAX1_15/A 0 17.052391f **FLOATING
C1033 MUX2X1_22/B 0 6.498059f **FLOATING
C1034 HAX1_44/YS 0 8.01429f **FLOATING
C1035 HAX1_47/A 0 16.378378f **FLOATING
C1036 HAX1_45/YS 0 8.10309f **FLOATING
C1037 OR2X1_2/Y 0 35.903835f **FLOATING
C1038 NOR2X1_2/A 0 20.4699f **FLOATING
C1039 FAX1_1/A 0 20.932802f **FLOATING
C1040 FAX1_9/C 0 15.587669f **FLOATING
C1041 FAX1_9/B 0 15.85902f **FLOATING
C1042 FAX1_9/A 0 17.728199f **FLOATING
C1043 FAX1_13/A 0 17.99703f **FLOATING
C1044 INVX2_3/Y 0 34.182274f **FLOATING
C1045 HAX1_31/B 0 17.81208f **FLOATING
C1046 FAX1_12/C 0 14.959739f **FLOATING
C1047 FAX1_12/A 0 17.49441f **FLOATING
C1048 NOR2X1_27/B 0 31.420958f **FLOATING
C1049 NOR2X1_32/B 0 31.622597f **FLOATING
C1050 INVX2_4/Y 0 33.29524f **FLOATING
C1051 FAX1_4/B 0 16.824091f **FLOATING
C1052 FAX1_0/A 0 23.969398f **FLOATING
C1053 FAX1_16/A 0 14.827169f **FLOATING
C1054 FAX1_2/YS 0 21.949106f **FLOATING
C1055 MUX2X1_19/Y 0 9.66618f **FLOATING
C1056 HAX1_44/A 0 20.201937f **FLOATING
C1057 MUX2X1_17/B 0 6.84966f **FLOATING
C1058 FAX1_1/YS 0 20.897366f **FLOATING
C1059 XNOR2X1_6/Y 0 9.26847f **FLOATING
C1060 NOR2X1_3/Y 0 19.119001f **FLOATING
C1061 XNOR2X1_7/A 0 23.04702f **FLOATING
C1062 FAX1_0/C 0 12.739349f **FLOATING
C1063 FAX1_0/YS 0 24.157558f **FLOATING
C1064 FAX1_7/YS 0 18.668459f **FLOATING
C1065 FAX1_6/C 0 13.73325f **FLOATING
C1066 FAX1_6/B 0 16.352102f **FLOATING
C1067 FAX1_6/A 0 14.102133f **FLOATING
C1068 INVX2_17/Y 0 34.23489f **FLOATING
C1069 FAX1_5/A 0 20.326738f **FLOATING
C1070 FAX1_4/A 0 19.702621f **FLOATING
C1071 MUX2X1_12/B 0 7.11246f **FLOATING
C1072 HAX1_40/YS 0 8.01429f **FLOATING
C1073 OR2X1_4/Y 0 32.41662f **FLOATING
C1074 MUX2X1_8/Y 0 17.978369f **FLOATING
C1075 FAX1_0/YC 0 17.601389f **FLOATING
C1076 FAX1_5/YS 0 16.036558f **FLOATING
C1077 XOR2X1_7/A 0 14.12958f **FLOATING
C1078 XOR2X1_6/A 0 12.985261f **FLOATING
C1079 MUX2X1_7/B 0 6.498059f **FLOATING
C1080 MUX2X1_5/Y 0 15.590641f **FLOATING
C1081 XOR2X1_8/Y 0 22.616922f **FLOATING
C1082 FAX1_4/YS 0 14.88312f **FLOATING
C1083 HAX1_41/YS 0 8.10309f **FLOATING
C1084 HAX1_43/A 0 16.685938f **FLOATING
C1085 MUX2X1_2/Y 0 9.2415f **FLOATING
C1086 XOR2X1_6/Y 0 14.668321f **FLOATING
C1087 OR2X1_5/B 0 8.8116f **FLOATING
C1088 OR2X1_5/A 0 6.996f **FLOATING
C1089 HAX1_41/A 0 16.378378f **FLOATING
C1090 FAX1_4/YC 0 15.189781f **FLOATING
C1091 XOR2X1_0/A 0 17.5761f **FLOATING
C1092 NOR2X1_7/A 0 12.2829f **FLOATING
C1093 vdd 0 18.918516p **FLOATING
C1094 FAX1_6/YS 0 16.345291f **FLOATING
C1095 XNOR2X1_5/Y 0 11.54667f **FLOATING
C1096 XNOR2X1_5/a_2_6# 0 6.77121f **FLOATING
C1097 XNOR2X1_5/a_12_41# 0 7.905991f **FLOATING
C1098 OAI21X1_29/a_2_6# 0 2.78652f **FLOATING
C1099 OAI21X1_18/a_2_6# 0 2.78652f **FLOATING
C1100 INVX2_88/Y 0 9.44856f **FLOATING
C1101 INVX2_44/Y 0 11.615879f **FLOATING
C1102 INVX2_33/Y 0 5.96766f **FLOATING
C1103 out_temp_cleared[12] 0 29.68209f **FLOATING
C1104 INVX2_259/Y 0 0.174577p **FLOATING
C1105 OAI22X1_2/a_2_6# 0 4.25172f **FLOATING
C1106 OAI22X1_50/Y 0 9.866341f **FLOATING
C1107 AOI22X1_62/a_2_54# 0 6.66f **FLOATING
C1108 AOI22X1_73/a_2_54# 0 6.66f **FLOATING
C1109 AOI22X1_40/a_2_54# 0 6.66f **FLOATING
C1110 AOI22X1_51/a_2_54# 0 6.66f **FLOATING
C1111 NAND2X1_97/Y 0 6.87006f **FLOATING
C1112 OAI21X1_57/B 0 7.08252f **FLOATING
C1113 OAI21X1_45/C 0 6.87006f **FLOATING
C1114 OAI21X1_13/C 0 6.87006f **FLOATING
C1115 OR2X1_6/Y 0 39.649754f **FLOATING
C1116 DFFNEGX1_140/a_66_6# 0 6.40992f **FLOATING
C1117 DFFNEGX1_140/a_23_6# 0 6.85692f **FLOATING
C1118 DFFNEGX1_140/a_34_4# 0 4.93023f **FLOATING
C1119 DFFNEGX1_140/a_2_6# 0 9.33504f **FLOATING
C1120 OAI21X1_158/Y 0 12.98496f **FLOATING
C1121 MUX2X1_27/a_2_10# 0 6.0456f **FLOATING
C1122 MUX2X1_16/a_2_10# 0 6.0456f **FLOATING
C1123 AND2X2_4/a_2_6# 0 6.03567f **FLOATING
C1124 HAX1_8/a_38_6# 0 2.442f **FLOATING
C1125 HAX1_8/a_41_74# 0 5.99325f **FLOATING
C1126 HAX1_8/a_2_74# 0 7.65318f **FLOATING
C1127 DFFNEGX1_72/a_66_6# 0 6.40992f **FLOATING
C1128 out_temp_cleared[19] 0 18.78807f **FLOATING
C1129 DFFNEGX1_72/a_23_6# 0 6.85692f **FLOATING
C1130 DFFNEGX1_72/a_34_4# 0 4.93023f **FLOATING
C1131 DFFNEGX1_72/a_2_6# 0 9.33504f **FLOATING
C1132 DFFNEGX1_83/a_66_6# 0 6.40992f **FLOATING
C1133 DFFNEGX1_83/a_23_6# 0 6.85692f **FLOATING
C1134 DFFNEGX1_83/a_34_4# 0 4.93023f **FLOATING
C1135 DFFNEGX1_83/a_2_6# 0 9.33504f **FLOATING
C1136 DFFNEGX1_94/a_66_6# 0 6.40992f **FLOATING
C1137 DFFNEGX1_94/a_23_6# 0 6.85692f **FLOATING
C1138 DFFNEGX1_94/a_34_4# 0 4.93023f **FLOATING
C1139 DFFNEGX1_94/a_2_6# 0 9.33504f **FLOATING
C1140 INVX2_216/Y 0 10.173361f **FLOATING
C1141 DFFNEGX1_61/a_66_6# 0 6.40992f **FLOATING
C1142 DFFNEGX1_61/a_23_6# 0 6.85692f **FLOATING
C1143 DFFNEGX1_61/a_34_4# 0 4.93023f **FLOATING
C1144 DFFNEGX1_61/a_2_6# 0 9.33504f **FLOATING
C1145 DFFNEGX1_50/a_66_6# 0 6.40992f **FLOATING
C1146 DFFNEGX1_50/a_23_6# 0 6.85692f **FLOATING
C1147 DFFNEGX1_50/a_34_4# 0 4.93023f **FLOATING
C1148 DFFNEGX1_50/a_2_6# 0 9.33504f **FLOATING
C1149 XNOR2X1_4/Y 0 9.22011f **FLOATING
C1150 XNOR2X1_4/a_2_6# 0 6.77121f **FLOATING
C1151 XNOR2X1_4/a_12_41# 0 7.905991f **FLOATING
C1152 INVX2_238/A 0 14.823421f **FLOATING
C1153 INVX2_241/A 0 8.48274f **FLOATING
C1154 OAI21X1_39/a_2_6# 0 2.78652f **FLOATING
C1155 OAI21X1_28/a_2_6# 0 2.78652f **FLOATING
C1156 OAI21X1_17/a_2_6# 0 2.78652f **FLOATING
C1157 OAI21X1_17/C 0 6.86169f **FLOATING
C1158 out_temp_decoded[16] 0 14.53077f **FLOATING
C1159 INVX2_43/Y 0 10.14474f **FLOATING
C1160 out_temp_cleared[2] 0 19.290129f **FLOATING
C1161 OAI22X1_1/a_2_6# 0 4.25172f **FLOATING
C1162 AOI22X1_61/a_2_54# 0 6.66f **FLOATING
C1163 AOI22X1_72/a_2_54# 0 6.66f **FLOATING
C1164 INVX2_51/Y 0 12.18555f **FLOATING
C1165 AOI22X1_50/a_2_54# 0 6.66f **FLOATING
C1166 OAI21X1_29/C 0 6.87006f **FLOATING
C1167 MUX2X1_26/Y 0 6.36198f **FLOATING
C1168 MUX2X1_26/a_2_10# 0 6.0456f **FLOATING
C1169 MUX2X1_15/a_2_10# 0 6.0456f **FLOATING
C1170 HAX1_33/A 0 14.034389f **FLOATING
C1171 AND2X2_3/a_2_6# 0 6.03567f **FLOATING
C1172 HAX1_7/a_38_6# 0 2.442f **FLOATING
C1173 HAX1_7/a_41_74# 0 5.99325f **FLOATING
C1174 HAX1_7/a_2_74# 0 7.65318f **FLOATING
C1175 DFFNEGX1_71/a_66_6# 0 6.40992f **FLOATING
C1176 DFFNEGX1_71/a_23_6# 0 6.85692f **FLOATING
C1177 DFFNEGX1_71/a_34_4# 0 4.93023f **FLOATING
C1178 DFFNEGX1_71/a_2_6# 0 9.33504f **FLOATING
C1179 DFFNEGX1_82/a_66_6# 0 6.40992f **FLOATING
C1180 DFFNEGX1_82/a_23_6# 0 6.85692f **FLOATING
C1181 DFFNEGX1_82/a_34_4# 0 4.93023f **FLOATING
C1182 DFFNEGX1_82/a_2_6# 0 9.33504f **FLOATING
C1183 DFFNEGX1_93/a_66_6# 0 6.40992f **FLOATING
C1184 DFFNEGX1_93/a_23_6# 0 6.85692f **FLOATING
C1185 DFFNEGX1_93/a_34_4# 0 4.93023f **FLOATING
C1186 DFFNEGX1_93/a_2_6# 0 9.33504f **FLOATING
C1187 DFFNEGX1_60/a_66_6# 0 6.40992f **FLOATING
C1188 DFFNEGX1_60/a_23_6# 0 6.85692f **FLOATING
C1189 DFFNEGX1_60/a_34_4# 0 4.93023f **FLOATING
C1190 DFFNEGX1_60/a_2_6# 0 9.33504f **FLOATING
C1191 XNOR2X1_3/a_2_6# 0 6.77121f **FLOATING
C1192 XNOR2X1_3/a_12_41# 0 7.905991f **FLOATING
C1193 AND2X2_19/a_2_6# 0 6.03567f **FLOATING
C1194 OAI21X1_27/a_2_6# 0 2.78652f **FLOATING
C1195 OAI21X1_38/a_2_6# 0 2.78652f **FLOATING
C1196 OAI21X1_49/a_2_6# 0 2.78652f **FLOATING
C1197 OAI21X1_49/Y 0 10.32552f **FLOATING
C1198 OAI21X1_16/a_2_6# 0 2.78652f **FLOATING
C1199 INVX2_86/Y 0 14.119862f **FLOATING
C1200 INVX2_31/A 0 19.663923f **FLOATING
C1201 HAX1_7/YS 0 10.12317f **FLOATING
C1202 XOR2X1_1/A 0 13.27659f **FLOATING
C1203 HAX1_7/B 0 13.508699f **FLOATING
C1204 OAI22X1_0/a_2_6# 0 4.25172f **FLOATING
C1205 OAI22X1_54/Y 0 9.832621f **FLOATING
C1206 AOI22X1_71/a_2_54# 0 6.66f **FLOATING
C1207 AOI22X1_60/a_2_54# 0 6.66f **FLOATING
C1208 OAI21X1_65/C 0 6.87006f **FLOATING
C1209 out_temp_index[0] 0 17.025751f **FLOATING
C1210 NOR2X1_119/B 0 10.753769f **FLOATING
C1211 MUX2X1_14/Y 0 9.97854f **FLOATING
C1212 MUX2X1_14/A 0 6.05058f **FLOATING
C1213 MUX2X1_14/a_2_10# 0 6.0456f **FLOATING
C1214 MUX2X1_25/a_2_10# 0 6.0456f **FLOATING
C1215 FAX1_10/A 0 14.75937f **FLOATING
C1216 INVX2_58/Y 0 7.020599f **FLOATING
C1217 AND2X2_2/a_2_6# 0 6.03567f **FLOATING
C1218 INVX2_27/Y 0 8.093459f **FLOATING
C1219 HAX1_6/a_38_6# 0 2.442f **FLOATING
C1220 HAX1_6/YS 0 6.99546f **FLOATING
C1221 HAX1_6/a_41_74# 0 5.99325f **FLOATING
C1222 HAX1_6/a_2_74# 0 7.65318f **FLOATING
C1223 DFFNEGX1_92/a_66_6# 0 6.40992f **FLOATING
C1224 DFFNEGX1_92/a_23_6# 0 6.85692f **FLOATING
C1225 DFFNEGX1_92/a_34_4# 0 4.93023f **FLOATING
C1226 DFFNEGX1_92/a_2_6# 0 9.33504f **FLOATING
C1227 DFFNEGX1_81/a_66_6# 0 6.40992f **FLOATING
C1228 DFFNEGX1_81/a_23_6# 0 6.85692f **FLOATING
C1229 DFFNEGX1_81/a_34_4# 0 4.93023f **FLOATING
C1230 DFFNEGX1_81/a_2_6# 0 9.33504f **FLOATING
C1231 OAI22X1_18/Y 0 10.427939f **FLOATING
C1232 DFFNEGX1_70/a_66_6# 0 6.40992f **FLOATING
C1233 DFFNEGX1_70/a_23_6# 0 6.85692f **FLOATING
C1234 DFFNEGX1_70/a_34_4# 0 4.93023f **FLOATING
C1235 DFFNEGX1_70/a_2_6# 0 9.33504f **FLOATING
C1236 OAI22X1_7/Y 0 11.25366f **FLOATING
C1237 INVX2_68/Y 0 18.277023f **FLOATING
C1238 XNOR2X1_2/a_2_6# 0 6.77121f **FLOATING
C1239 XNOR2X1_2/a_12_41# 0 7.905991f **FLOATING
C1240 OAI21X1_43/C 0 7.94154f **FLOATING
C1241 AND2X2_18/a_2_6# 0 6.03567f **FLOATING
C1242 OAI21X1_59/a_2_6# 0 2.78652f **FLOATING
C1243 OAI21X1_59/C 0 6.86169f **FLOATING
C1244 OAI21X1_37/a_2_6# 0 2.78652f **FLOATING
C1245 OAI21X1_37/C 0 6.86169f **FLOATING
C1246 OAI21X1_48/a_2_6# 0 2.78652f **FLOATING
C1247 INVX2_244/A 0 6.92922f **FLOATING
C1248 OAI21X1_26/a_2_6# 0 2.78652f **FLOATING
C1249 OAI21X1_15/a_2_6# 0 2.78652f **FLOATING
C1250 OAI21X1_129/Y 0 8.025811f **FLOATING
C1251 AOI22X1_70/a_2_54# 0 6.66f **FLOATING
C1252 OAI21X1_55/C 0 8.08944f **FLOATING
C1253 INVX2_189/A 0 8.11314f **FLOATING
C1254 NOR2X1_118/B 0 12.02118f **FLOATING
C1255 MUX2X1_24/A 0 6.13938f **FLOATING
C1256 MUX2X1_24/a_2_10# 0 6.0456f **FLOATING
C1257 MUX2X1_13/a_2_10# 0 6.0456f **FLOATING
C1258 INVX2_239/Y 0 10.97868f **FLOATING
C1259 NOR2X1_39/Y 0 6.2739f **FLOATING
C1260 NOR2X1_83/Y 0 8.409901f **FLOATING
C1261 NOR2X1_86/Y 0 10.837259f **FLOATING
C1262 out_mines[1] 0 0.116304p **FLOATING
C1263 NOR2X1_119/Y 0 11.606281f **FLOATING
C1264 AND2X2_1/a_2_6# 0 6.03567f **FLOATING
C1265 HAX1_5/a_38_6# 0 2.442f **FLOATING
C1266 HAX1_5/YS 0 6.92886f **FLOATING
C1267 HAX1_5/a_41_74# 0 5.99325f **FLOATING
C1268 HAX1_5/a_2_74# 0 7.65318f **FLOATING
C1269 DFFNEGX1_91/a_66_6# 0 6.40992f **FLOATING
C1270 DFFNEGX1_91/a_23_6# 0 6.85692f **FLOATING
C1271 DFFNEGX1_91/a_34_4# 0 4.93023f **FLOATING
C1272 DFFNEGX1_91/a_2_6# 0 9.33504f **FLOATING
C1273 DFFNEGX1_80/a_66_6# 0 6.40992f **FLOATING
C1274 DFFNEGX1_80/a_23_6# 0 6.85692f **FLOATING
C1275 DFFNEGX1_80/a_34_4# 0 4.93023f **FLOATING
C1276 DFFNEGX1_80/a_2_6# 0 9.33504f **FLOATING
C1277 INVX2_78/Y 0 27.014141f **FLOATING
C1278 XNOR2X1_1/a_2_6# 0 6.77121f **FLOATING
C1279 XNOR2X1_1/a_12_41# 0 7.905991f **FLOATING
C1280 AND2X2_17/a_2_6# 0 6.03567f **FLOATING
C1281 AND2X2_17/A 0 17.98425f **FLOATING
C1282 OAI21X1_58/a_2_6# 0 2.78652f **FLOATING
C1283 OAI21X1_69/a_2_6# 0 2.78652f **FLOATING
C1284 OAI21X1_47/a_2_6# 0 2.78652f **FLOATING
C1285 OAI21X1_36/a_2_6# 0 2.78652f **FLOATING
C1286 INVX2_225/A 0 6.0849f **FLOATING
C1287 OAI21X1_25/a_2_6# 0 2.78652f **FLOATING
C1288 OAI21X1_14/a_2_6# 0 2.78652f **FLOATING
C1289 INVX2_62/Y 0 5.62842f **FLOATING
C1290 HAX1_8/YS 0 9.83463f **FLOATING
C1291 HAX1_8/B 0 12.3081f **FLOATING
C1292 MUX2X1_34/A 0 6.13938f **FLOATING
C1293 MUX2X1_34/a_2_10# 0 6.0456f **FLOATING
C1294 XNOR2X1_3/A 0 22.189049f **FLOATING
C1295 MUX2X1_23/a_2_10# 0 6.0456f **FLOATING
C1296 MUX2X1_12/Y 0 6.36198f **FLOATING
C1297 MUX2X1_12/a_2_10# 0 6.0456f **FLOATING
C1298 INVX2_238/Y 0 10.02582f **FLOATING
C1299 NOR2X1_49/Y 0 6.2739f **FLOATING
C1300 FAX1_17/C 0 16.55049f **FLOATING
C1301 AND2X2_0/a_2_6# 0 6.03567f **FLOATING
C1302 HAX1_4/a_38_6# 0 2.442f **FLOATING
C1303 HAX1_4/YS 0 6.99546f **FLOATING
C1304 HAX1_4/a_41_74# 0 5.99325f **FLOATING
C1305 HAX1_4/a_2_74# 0 7.65318f **FLOATING
C1306 DFFNEGX1_90/a_66_6# 0 6.40992f **FLOATING
C1307 DFFNEGX1_90/a_23_6# 0 6.85692f **FLOATING
C1308 DFFNEGX1_90/a_34_4# 0 4.93023f **FLOATING
C1309 DFFNEGX1_90/a_2_6# 0 9.33504f **FLOATING
C1310 INVX2_93/Y 0 8.811f **FLOATING
C1311 INVX1_0/Y 0 5.6358f **FLOATING
C1312 XNOR2X1_0/Y 0 9.10131f **FLOATING
C1313 XNOR2X1_0/a_2_6# 0 6.77121f **FLOATING
C1314 XNOR2X1_0/a_12_41# 0 7.905991f **FLOATING
C1315 INVX2_237/A 0 9.07926f **FLOATING
C1316 AND2X2_16/a_2_6# 0 6.03567f **FLOATING
C1317 OAI21X1_79/a_2_6# 0 2.78652f **FLOATING
C1318 NOR2X1_94/A 0 6.771f **FLOATING
C1319 OAI21X1_57/a_2_6# 0 2.78652f **FLOATING
C1320 OAI21X1_68/a_2_6# 0 2.78652f **FLOATING
C1321 OAI21X1_46/a_2_6# 0 2.78652f **FLOATING
C1322 OAI21X1_24/a_2_6# 0 2.78652f **FLOATING
C1323 OAI21X1_35/a_2_6# 0 2.78652f **FLOATING
C1324 OAI21X1_13/a_2_6# 0 2.78652f **FLOATING
C1325 out_temp_decoded[1] 0 12.277711f **FLOATING
C1326 out_temp_decoded[19] 0 21.382141f **FLOATING
C1327 OAI21X1_83/C 0 13.565429f **FLOATING
C1328 MUX2X1_33/a_2_10# 0 6.0456f **FLOATING
C1329 MUX2X1_22/Y 0 7.2063f **FLOATING
C1330 MUX2X1_22/a_2_10# 0 6.0456f **FLOATING
C1331 MUX2X1_11/Y 0 8.18202f **FLOATING
C1332 MUX2X1_11/a_2_10# 0 6.0456f **FLOATING
C1333 INVX2_215/Y 0 10.993021f **FLOATING
C1334 INVX2_204/Y 0 12.089221f **FLOATING
C1335 INVX2_204/A 0 8.11314f **FLOATING
C1336 NOR2X1_48/Y 0 9.13794f **FLOATING
C1337 NOR2X1_59/Y 0 6.2739f **FLOATING
C1338 NOR2X1_59/B 0 25.510616f **FLOATING
C1339 NOR2X1_37/Y 0 11.33742f **FLOATING
C1340 FAX1_18/B 0 17.56059f **FLOATING
C1341 INVX2_131/Y 0 16.850458f **FLOATING
C1342 HAX1_3/a_38_6# 0 2.442f **FLOATING
C1343 HAX1_3/a_41_74# 0 5.99325f **FLOATING
C1344 HAX1_3/a_2_74# 0 7.65318f **FLOATING
C1345 AND2X2_15/a_2_6# 0 6.03567f **FLOATING
C1346 OR2X1_16/a_2_54# 0 6.27999f **FLOATING
C1347 OAI21X1_89/a_2_6# 0 2.78652f **FLOATING
C1348 OAI21X1_78/a_2_6# 0 2.78652f **FLOATING
C1349 OAI21X1_67/a_2_6# 0 2.78652f **FLOATING
C1350 OAI21X1_56/a_2_6# 0 2.78652f **FLOATING
C1351 OAI21X1_23/a_2_6# 0 2.78652f **FLOATING
C1352 OAI21X1_45/a_2_6# 0 2.78652f **FLOATING
C1353 OAI21X1_34/a_2_6# 0 2.78652f **FLOATING
C1354 OAI21X1_12/a_2_6# 0 2.78652f **FLOATING
C1355 out_global_score[27] 0 18.269371f **FLOATING
C1356 MUX2X1_32/a_2_10# 0 6.0456f **FLOATING
C1357 MUX2X1_21/Y 0 8.18202f **FLOATING
C1358 MUX2X1_21/a_2_10# 0 6.0456f **FLOATING
C1359 MUX2X1_10/a_2_10# 0 6.0456f **FLOATING
C1360 INVX2_203/A 0 9.661799f **FLOATING
C1361 NAND3X1_36/Y 0 6.97965f **FLOATING
C1362 NAND3X1_50/Y 0 9.911551f **FLOATING
C1363 HAX1_2/a_38_6# 0 2.442f **FLOATING
C1364 HAX1_2/a_41_74# 0 5.99325f **FLOATING
C1365 HAX1_2/a_2_74# 0 7.65318f **FLOATING
C1366 AND2X2_14/a_2_6# 0 6.03567f **FLOATING
C1367 OR2X1_15/a_2_54# 0 6.27999f **FLOATING
C1368 OAI21X1_99/a_2_6# 0 2.78652f **FLOATING
C1369 OAI21X1_99/C 0 10.55064f **FLOATING
C1370 OAI21X1_88/a_2_6# 0 2.78652f **FLOATING
C1371 OAI21X1_77/a_2_6# 0 2.78652f **FLOATING
C1372 OAI21X1_66/a_2_6# 0 2.78652f **FLOATING
C1373 OAI21X1_55/a_2_6# 0 2.78652f **FLOATING
C1374 OAI21X1_55/Y 0 12.530281f **FLOATING
C1375 OAI21X1_33/a_2_6# 0 2.78652f **FLOATING
C1376 OAI21X1_22/a_2_6# 0 2.78652f **FLOATING
C1377 OAI21X1_44/a_2_6# 0 2.78652f **FLOATING
C1378 OAI21X1_11/a_2_6# 0 2.78652f **FLOATING
C1379 OAI21X1_11/C 0 6.86169f **FLOATING
C1380 HAX1_0/YC 0 11.435069f **FLOATING
C1381 AOI21X1_2/A 0 37.655674f **FLOATING
C1382 HAX1_48/YS 0 11.26437f **FLOATING
C1383 MUX2X1_31/a_2_10# 0 6.0456f **FLOATING
C1384 MUX2X1_20/a_2_10# 0 6.0456f **FLOATING
C1385 INVX2_257/Y 0 0.106892p **FLOATING
C1386 XOR2X1_14/Y 0 9.064739f **FLOATING
C1387 NOR2X1_35/Y 0 10.484581f **FLOATING
C1388 HAX1_32/A 0 12.496619f **FLOATING
C1389 INVX2_2/Y 0 30.08525f **FLOATING
C1390 BUFX2_25/A 0 37.04236f **FLOATING
C1391 BUFX2_21/A 0 21.442198f **FLOATING
C1392 HAX1_1/a_38_6# 0 2.442f **FLOATING
C1393 HAX1_1/a_41_74# 0 5.99325f **FLOATING
C1394 HAX1_1/a_2_74# 0 7.65318f **FLOATING
C1395 AND2X2_13/a_2_6# 0 6.03567f **FLOATING
C1396 OR2X1_14/a_2_54# 0 6.27999f **FLOATING
C1397 OAI21X1_98/a_2_6# 0 2.78652f **FLOATING
C1398 OAI21X1_65/a_2_6# 0 2.78652f **FLOATING
C1399 OAI21X1_76/a_2_6# 0 2.78652f **FLOATING
C1400 OAI21X1_76/C 0 12.496051f **FLOATING
C1401 OAI21X1_87/a_2_6# 0 2.78652f **FLOATING
C1402 OAI21X1_21/a_2_6# 0 2.78652f **FLOATING
C1403 INVX2_229/Y 0 16.069983f **FLOATING
C1404 OAI21X1_43/a_2_6# 0 2.78652f **FLOATING
C1405 OAI21X1_43/Y 0 12.073442f **FLOATING
C1406 OAI21X1_32/a_2_6# 0 2.78652f **FLOATING
C1407 INVX2_242/A 0 6.0849f **FLOATING
C1408 OAI21X1_54/a_2_6# 0 2.78652f **FLOATING
C1409 OAI21X1_10/a_2_6# 0 2.78652f **FLOATING
C1410 OR2X1_2/B 0 8.8116f **FLOATING
C1411 BUFX2_7/Y 0 15.099481f **FLOATING
C1412 NOR2X1_124/B 0 6.08568f **FLOATING
C1413 MUX2X1_30/a_2_10# 0 6.0456f **FLOATING
C1414 OR2X1_11/B 0 0.122423p **FLOATING
C1415 INVX2_245/Y 0 12.208021f **FLOATING
C1416 INVX2_201/Y 0 11.646931f **FLOATING
C1417 INVX2_201/A 0 8.03022f **FLOATING
C1418 NOR2X1_78/Y 0 15.20712f **FLOATING
C1419 NOR2X1_56/Y 0 6.2739f **FLOATING
C1420 HAX1_33/B 0 13.62348f **FLOATING
C1421 FAX1_17/A 0 21.12963f **FLOATING
C1422 NAND3X1_34/C 0 13.30176f **FLOATING
C1423 OAI21X1_77/B 0 9.784981f **FLOATING
C1424 HAX1_0/a_38_6# 0 2.442f **FLOATING
C1425 HAX1_0/a_41_74# 0 5.99325f **FLOATING
C1426 HAX1_0/a_2_74# 0 7.65318f **FLOATING
C1427 NOR2X1_68/Y 0 10.19124f **FLOATING
C1428 AND2X2_12/a_2_6# 0 6.03567f **FLOATING
C1429 OR2X1_13/a_2_54# 0 6.27999f **FLOATING
C1430 OR2X1_13/B 0 17.375288f **FLOATING
C1431 OAI21X1_97/a_2_6# 0 2.78652f **FLOATING
C1432 OAI21X1_64/a_2_6# 0 2.78652f **FLOATING
C1433 INVX2_256/A 0 17.23056f **FLOATING
C1434 OAI21X1_75/a_2_6# 0 2.78652f **FLOATING
C1435 NOR2X1_89/B 0 7.529939f **FLOATING
C1436 OAI21X1_86/a_2_6# 0 2.78652f **FLOATING
C1437 OAI21X1_31/a_2_6# 0 2.78652f **FLOATING
C1438 OAI21X1_31/C 0 6.86169f **FLOATING
C1439 OAI21X1_42/a_2_6# 0 2.78652f **FLOATING
C1440 OAI21X1_46/B 0 22.598103f **FLOATING
C1441 OAI21X1_53/a_2_6# 0 2.78652f **FLOATING
C1442 OAI21X1_53/C 0 10.92264f **FLOATING
C1443 OAI21X1_20/a_2_6# 0 2.78652f **FLOATING
C1444 OR2X1_4/B 0 8.8116f **FLOATING
C1445 OR2X1_16/B 0 11.39076f **FLOATING
C1446 out_temp_cleared[24] 0 16.00557f **FLOATING
C1447 INVX2_244/Y 0 10.245f **FLOATING
C1448 INVX2_200/A 0 8.11314f **FLOATING
C1449 NOR2X1_33/Y 0 9.98682f **FLOATING
C1450 NOR2X1_22/B 0 38.1562f **FLOATING
C1451 FAX1_18/A 0 18.15975f **FLOATING
C1452 NOR2X1_89/Y 0 9.094381f **FLOATING
C1453 AOI21X1_6/Y 0 20.320797f **FLOATING
C1454 NAND3X1_44/A 0 9.394199f **FLOATING
C1455 OAI21X1_8/A 0 53.754803f **FLOATING
C1456 out_temp_cleared[20] 0 27.070229f **FLOATING
C1457 AND2X2_11/a_2_6# 0 6.03567f **FLOATING
C1458 OR2X1_12/a_2_54# 0 6.27999f **FLOATING
C1459 OAI21X1_85/a_2_6# 0 2.78652f **FLOATING
C1460 OAI21X1_96/a_2_6# 0 2.78652f **FLOATING
C1461 OAI21X1_74/a_2_6# 0 2.78652f **FLOATING
C1462 OAI21X1_63/a_2_6# 0 2.78652f **FLOATING
C1463 OAI21X1_63/Y 0 6.5451f **FLOATING
C1464 OAI21X1_41/a_2_6# 0 2.78652f **FLOATING
C1465 OAI21X1_30/a_2_6# 0 2.78652f **FLOATING
C1466 OAI21X1_52/a_2_6# 0 2.78652f **FLOATING
C1467 OAI22X1_19/a_2_6# 0 4.25172f **FLOATING
C1468 OR2X1_9/a_2_54# 0 6.27999f **FLOATING
C1469 out_temp_data_in[4] 0 91.656006f **FLOATING
C1470 NOR2X1_98/Y 0 6.8172f **FLOATING
C1471 NOR2X1_43/B 0 6.08568f **FLOATING
C1472 NOR2X1_54/Y 0 6.2739f **FLOATING
C1473 HAX1_34/A 0 9.284161f **FLOATING
C1474 NOR2X1_77/B 0 13.432339f **FLOATING
C1475 NAND3X1_41/B 0 8.3577f **FLOATING
C1476 AOI21X1_20/Y 0 12.31401f **FLOATING
C1477 AND2X2_10/a_2_6# 0 6.03567f **FLOATING
C1478 OR2X1_11/a_2_54# 0 6.27999f **FLOATING
C1479 OAI21X1_84/a_2_6# 0 2.78652f **FLOATING
C1480 OAI21X1_95/a_2_6# 0 2.78652f **FLOATING
C1481 OAI21X1_95/C 0 6.86169f **FLOATING
C1482 OAI21X1_73/a_2_6# 0 2.78652f **FLOATING
C1483 OAI21X1_62/a_2_6# 0 2.78652f **FLOATING
C1484 OAI21X1_40/a_2_6# 0 2.78652f **FLOATING
C1485 OAI21X1_51/a_2_6# 0 2.78652f **FLOATING
C1486 OAI22X1_29/a_2_6# 0 4.25172f **FLOATING
C1487 OAI22X1_18/a_2_6# 0 4.25172f **FLOATING
C1488 INVX2_230/Y 0 13.028521f **FLOATING
C1489 OR2X1_8/a_2_54# 0 6.27999f **FLOATING
C1490 NOR2X1_110/Y 0 6.311941f **FLOATING
C1491 NOR2X1_97/Y 0 10.38471f **FLOATING
C1492 INVX2_240/A 0 11.18778f **FLOATING
C1493 OAI21X1_91/C 0 10.70784f **FLOATING
C1494 OAI21X1_6/A 0 19.46268f **FLOATING
C1495 out_mines[21] 0 69.52224f **FLOATING
C1496 OR2X1_10/a_2_54# 0 6.27999f **FLOATING
C1497 OAI21X1_83/a_2_6# 0 2.78652f **FLOATING
C1498 OAI21X1_83/Y 0 13.13226f **FLOATING
C1499 OAI21X1_94/a_2_6# 0 2.78652f **FLOATING
C1500 OAI21X1_61/a_2_6# 0 2.78652f **FLOATING
C1501 OAI21X1_61/Y 0 9.85554f **FLOATING
C1502 XNOR2X1_20/Y 0 7.55235f **FLOATING
C1503 OAI21X1_72/a_2_6# 0 2.78652f **FLOATING
C1504 OAI21X1_72/C 0 11.01525f **FLOATING
C1505 OAI21X1_50/a_2_6# 0 2.78652f **FLOATING
C1506 INVX2_222/A 0 11.797681f **FLOATING
C1507 OAI22X1_28/a_2_6# 0 4.25172f **FLOATING
C1508 OAI22X1_39/a_2_6# 0 4.25172f **FLOATING
C1509 OAI22X1_17/a_2_6# 0 4.25172f **FLOATING
C1510 OR2X1_7/a_2_54# 0 6.27999f **FLOATING
C1511 BUFX2_19/a_2_6# 0 5.63946f **FLOATING
C1512 NOR2X1_7/B 0 15.043921f **FLOATING
C1513 NOR2X1_41/Y 0 8.64978f **FLOATING
C1514 INVX2_224/A 0 15.098761f **FLOATING
C1515 OAI21X1_81/C 0 11.485651f **FLOATING
C1516 out_temp_decoded[2] 0 14.84049f **FLOATING
C1517 INVX2_127/A 0 45.089657f **FLOATING
C1518 OAI21X1_82/a_2_6# 0 2.78652f **FLOATING
C1519 OAI21X1_93/a_2_6# 0 2.78652f **FLOATING
C1520 OAI21X1_60/a_2_6# 0 2.78652f **FLOATING
C1521 OAI21X1_60/C 0 7.93494f **FLOATING
C1522 OAI21X1_71/a_2_6# 0 2.78652f **FLOATING
C1523 OAI22X1_27/a_2_6# 0 4.25172f **FLOATING
C1524 OAI22X1_38/a_2_6# 0 4.25172f **FLOATING
C1525 OAI22X1_38/C 0 17.019361f **FLOATING
C1526 OAI22X1_16/a_2_6# 0 4.25172f **FLOATING
C1527 OAI22X1_49/a_2_6# 0 4.25172f **FLOATING
C1528 OR2X1_6/a_2_54# 0 6.27999f **FLOATING
C1529 AOI21X1_19/a_2_54# 0 4.3068f **FLOATING
C1530 HAX1_30/B 0 14.47212f **FLOATING
C1531 BUFX2_18/a_2_6# 0 5.63946f **FLOATING
C1532 XNOR2X1_19/a_2_6# 0 6.77121f **FLOATING
C1533 XNOR2X1_19/a_12_41# 0 7.905991f **FLOATING
C1534 AOI21X1_4/Y 0 13.812331f **FLOATING
C1535 NAND2X1_6/B 0 14.605862f **FLOATING
C1536 FAX1_9/a_46_6# 0 2.442f **FLOATING
C1537 FAX1_9/a_2_6# 0 2.5308f **FLOATING
C1538 FAX1_9/a_46_54# 0 4.1292f **FLOATING
C1539 FAX1_9/a_2_54# 0 4.3068f **FLOATING
C1540 FAX1_9/a_70_6# 0 6.54516f **FLOATING
C1541 FAX1_9/a_25_6# 0 9.36792f **FLOATING
C1542 NOR2X1_95/Y 0 12.013378f **FLOATING
C1543 out_temp_cleared[13] 0 25.98684f **FLOATING
C1544 NOR2X1_73/Y 0 14.16606f **FLOATING
C1545 AND2X2_16/A 0 9.07974f **FLOATING
C1546 out_temp_decoded[20] 0 24.89595f **FLOATING
C1547 INVX2_5/Y 0 6.71694f **FLOATING
C1548 OAI21X1_92/a_2_6# 0 2.78652f **FLOATING
C1549 OAI21X1_70/a_2_6# 0 2.78652f **FLOATING
C1550 INVX2_80/A 0 6.0849f **FLOATING
C1551 OAI21X1_81/a_2_6# 0 2.78652f **FLOATING
C1552 AOI21X1_7/C 0 10.43922f **FLOATING
C1553 OAI22X1_59/a_2_6# 0 4.25172f **FLOATING
C1554 OAI22X1_37/a_2_6# 0 4.25172f **FLOATING
C1555 OAI22X1_26/a_2_6# 0 4.25172f **FLOATING
C1556 OAI22X1_48/a_2_6# 0 4.25172f **FLOATING
C1557 OAI22X1_15/a_2_6# 0 4.25172f **FLOATING
C1558 OR2X1_5/a_2_54# 0 6.27999f **FLOATING
C1559 AOI21X1_18/a_2_54# 0 4.3068f **FLOATING
C1560 BUFX2_17/a_2_6# 0 5.63946f **FLOATING
C1561 OR2X1_3/B 0 8.670599f **FLOATING
C1562 XNOR2X1_18/a_2_6# 0 6.77121f **FLOATING
C1563 XNOR2X1_18/a_12_41# 0 7.905991f **FLOATING
C1564 XNOR2X1_29/a_2_6# 0 6.77121f **FLOATING
C1565 XNOR2X1_29/a_12_41# 0 7.905991f **FLOATING
C1566 NOR2X1_79/B 0 11.101291f **FLOATING
C1567 HAX1_38/B 0 13.04418f **FLOATING
C1568 FAX1_8/a_46_6# 0 2.442f **FLOATING
C1569 FAX1_8/a_2_6# 0 2.5308f **FLOATING
C1570 FAX1_8/a_46_54# 0 4.1292f **FLOATING
C1571 FAX1_8/a_2_54# 0 4.3068f **FLOATING
C1572 FAX1_8/a_70_6# 0 6.54516f **FLOATING
C1573 FAX1_8/a_25_6# 0 9.36792f **FLOATING
C1574 FAX1_8/B 0 13.157999f **FLOATING
C1575 BUFX2_16/Y 0 0.19702p **FLOATING
C1576 NOR2X1_72/Y 0 6.311941f **FLOATING
C1577 out_decode 0 23.59515f **FLOATING
C1578 OAI21X1_23/C 0 8.146441f **FLOATING
C1579 OAI21X1_90/C 0 20.199959f **FLOATING
C1580 INVX2_233/A 0 11.649938f **FLOATING
C1581 FAX1_18/a_46_6# 0 2.442f **FLOATING
C1582 FAX1_18/a_2_6# 0 2.5308f **FLOATING
C1583 FAX1_18/a_46_54# 0 4.1292f **FLOATING
C1584 FAX1_18/a_2_54# 0 4.3068f **FLOATING
C1585 FAX1_18/a_70_6# 0 6.54516f **FLOATING
C1586 FAX1_18/a_25_6# 0 9.36792f **FLOATING
C1587 OAI21X1_91/a_2_6# 0 2.78652f **FLOATING
C1588 OAI21X1_80/a_2_6# 0 2.78652f **FLOATING
C1589 OAI22X1_69/a_2_6# 0 4.25172f **FLOATING
C1590 OAI22X1_36/a_2_6# 0 4.25172f **FLOATING
C1591 OAI22X1_58/a_2_6# 0 4.25172f **FLOATING
C1592 OAI22X1_47/a_2_6# 0 4.25172f **FLOATING
C1593 OAI22X1_25/a_2_6# 0 4.25172f **FLOATING
C1594 OAI22X1_14/a_2_6# 0 4.25172f **FLOATING
C1595 OR2X1_4/a_2_54# 0 6.27999f **FLOATING
C1596 AOI21X1_17/a_2_54# 0 4.3068f **FLOATING
C1597 BUFX2_16/a_2_6# 0 5.63946f **FLOATING
C1598 XNOR2X1_28/a_2_6# 0 6.77121f **FLOATING
C1599 XNOR2X1_28/a_12_41# 0 7.905991f **FLOATING
C1600 INVX2_39/A 0 24.355228f **FLOATING
C1601 XNOR2X1_17/a_2_6# 0 6.77121f **FLOATING
C1602 XNOR2X1_17/a_12_41# 0 7.905991f **FLOATING
C1603 NOR2X1_79/A 0 13.206931f **FLOATING
C1604 AOI21X1_9/a_2_54# 0 4.3068f **FLOATING
C1605 HAX1_40/B 0 12.93174f **FLOATING
C1606 FAX1_7/a_46_6# 0 2.442f **FLOATING
C1607 FAX1_7/a_2_6# 0 2.5308f **FLOATING
C1608 FAX1_7/a_46_54# 0 4.1292f **FLOATING
C1609 FAX1_7/a_2_54# 0 4.3068f **FLOATING
C1610 FAX1_7/a_70_6# 0 6.54516f **FLOATING
C1611 FAX1_7/a_25_6# 0 9.36792f **FLOATING
C1612 BUFX2_9/a_2_6# 0 5.63946f **FLOATING
C1613 NOR2X1_71/Y 0 9.2895f **FLOATING
C1614 NOR2X1_71/B 0 6.08568f **FLOATING
C1615 NOR2X1_61/Y 0 14.768552f **FLOATING
C1616 FAX1_17/a_46_6# 0 2.442f **FLOATING
C1617 FAX1_17/a_2_6# 0 2.5308f **FLOATING
C1618 FAX1_17/a_46_54# 0 4.1292f **FLOATING
C1619 FAX1_17/a_2_54# 0 4.3068f **FLOATING
C1620 FAX1_17/a_70_6# 0 6.54516f **FLOATING
C1621 FAX1_17/a_25_6# 0 9.36792f **FLOATING
C1622 out_temp_cleared[18] 0 22.339352f **FLOATING
C1623 OAI22X1_5/C 0 0.105496p **FLOATING
C1624 OAI21X1_90/a_2_6# 0 2.78652f **FLOATING
C1625 DFFNEGX1_9/a_66_6# 0 6.40992f **FLOATING
C1626 DFFNEGX1_9/a_23_6# 0 6.85692f **FLOATING
C1627 DFFNEGX1_9/a_34_4# 0 4.93023f **FLOATING
C1628 DFFNEGX1_9/a_2_6# 0 9.33504f **FLOATING
C1629 INVX2_60/Y 0 21.3291f **FLOATING
C1630 OAI22X1_68/a_2_6# 0 4.25172f **FLOATING
C1631 OAI22X1_79/a_2_6# 0 4.25172f **FLOATING
C1632 OAI22X1_57/a_2_6# 0 4.25172f **FLOATING
C1633 OAI22X1_35/a_2_6# 0 4.25172f **FLOATING
C1634 OAI22X1_46/a_2_6# 0 4.25172f **FLOATING
C1635 OAI22X1_24/a_2_6# 0 4.25172f **FLOATING
C1636 OAI22X1_13/a_2_6# 0 4.25172f **FLOATING
C1637 INVX2_225/Y 0 12.67092f **FLOATING
C1638 OR2X1_3/a_2_54# 0 6.27999f **FLOATING
C1639 HAX1_19/a_38_6# 0 2.442f **FLOATING
C1640 HAX1_18/B 0 12.009359f **FLOATING
C1641 HAX1_19/a_41_74# 0 5.99325f **FLOATING
C1642 HAX1_19/a_2_74# 0 7.65318f **FLOATING
C1643 AOI21X1_16/a_2_54# 0 4.3068f **FLOATING
C1644 XOR2X1_7/Y 0 21.324808f **FLOATING
C1645 BUFX2_15/a_2_6# 0 5.63946f **FLOATING
C1646 XNOR2X1_27/a_2_6# 0 6.77121f **FLOATING
C1647 XNOR2X1_27/a_12_41# 0 7.905991f **FLOATING
C1648 XNOR2X1_16/a_2_6# 0 6.77121f **FLOATING
C1649 XNOR2X1_16/a_12_41# 0 7.905991f **FLOATING
C1650 AOI21X1_8/a_2_54# 0 4.3068f **FLOATING
C1651 INVX2_251/Y 0 0.103067p **FLOATING
C1652 FAX1_6/a_46_6# 0 2.442f **FLOATING
C1653 FAX1_6/a_2_6# 0 2.5308f **FLOATING
C1654 FAX1_6/a_46_54# 0 4.1292f **FLOATING
C1655 FAX1_6/a_2_54# 0 4.3068f **FLOATING
C1656 FAX1_6/a_70_6# 0 6.54516f **FLOATING
C1657 FAX1_6/a_25_6# 0 9.36792f **FLOATING
C1658 AOI22X1_65/Y 0 8.14098f **FLOATING
C1659 BUFX2_2/Y 0 15.007832f **FLOATING
C1660 BUFX2_8/a_2_6# 0 5.63946f **FLOATING
C1661 NOR2X1_70/Y 0 10.12821f **FLOATING
C1662 NOR2X1_81/Y 0 10.040161f **FLOATING
C1663 BUFX2_6/Y 0 17.117552f **FLOATING
C1664 FAX1_16/a_46_6# 0 2.442f **FLOATING
C1665 FAX1_16/a_2_6# 0 2.5308f **FLOATING
C1666 FAX1_16/a_46_54# 0 4.1292f **FLOATING
C1667 FAX1_16/a_2_54# 0 4.3068f **FLOATING
C1668 FAX1_16/a_70_6# 0 6.54516f **FLOATING
C1669 FAX1_16/a_25_6# 0 9.36792f **FLOATING
C1670 DFFNEGX1_8/a_66_6# 0 6.40992f **FLOATING
C1671 DFFNEGX1_8/a_23_6# 0 6.85692f **FLOATING
C1672 DFFNEGX1_8/a_34_4# 0 4.93023f **FLOATING
C1673 DFFNEGX1_8/a_2_6# 0 9.33504f **FLOATING
C1674 OAI22X1_78/a_2_6# 0 4.25172f **FLOATING
C1675 OAI22X1_67/a_2_6# 0 4.25172f **FLOATING
C1676 OAI22X1_56/a_2_6# 0 4.25172f **FLOATING
C1677 OAI22X1_45/a_2_6# 0 4.25172f **FLOATING
C1678 OAI22X1_34/a_2_6# 0 4.25172f **FLOATING
C1679 OAI22X1_23/a_2_6# 0 4.25172f **FLOATING
C1680 OAI22X1_12/a_2_6# 0 4.25172f **FLOATING
C1681 OAI21X1_7/A 0 12.80892f **FLOATING
C1682 INVX2_221/Y 0 16.088577f **FLOATING
C1683 OR2X1_2/a_2_54# 0 6.27999f **FLOATING
C1684 HAX1_29/a_38_6# 0 2.442f **FLOATING
C1685 HAX1_29/a_41_74# 0 5.99325f **FLOATING
C1686 HAX1_29/a_2_74# 0 7.65318f **FLOATING
C1687 out_global_score[0] 0 20.9754f **FLOATING
C1688 HAX1_18/a_38_6# 0 2.442f **FLOATING
C1689 HAX1_18/YS 0 7.70586f **FLOATING
C1690 HAX1_17/B 0 13.94946f **FLOATING
C1691 HAX1_18/a_41_74# 0 5.99325f **FLOATING
C1692 HAX1_18/a_2_74# 0 7.65318f **FLOATING
C1693 AOI21X1_15/a_2_54# 0 4.3068f **FLOATING
C1694 AOI21X1_26/a_2_54# 0 4.3068f **FLOATING
C1695 NAND3X1_57/Y 0 9.10041f **FLOATING
C1696 BUFX2_14/a_2_6# 0 5.63946f **FLOATING
C1697 BUFX2_25/a_2_6# 0 5.63946f **FLOATING
C1698 XNOR2X1_26/a_2_6# 0 6.77121f **FLOATING
C1699 XNOR2X1_26/a_12_41# 0 7.905991f **FLOATING
C1700 XNOR2X1_15/a_2_6# 0 6.77121f **FLOATING
C1701 XNOR2X1_15/a_12_41# 0 7.905991f **FLOATING
C1702 AOI21X1_7/a_2_54# 0 4.3068f **FLOATING
C1703 AOI21X1_7/A 0 10.7952f **FLOATING
C1704 HAX1_44/B 0 15.494401f **FLOATING
C1705 FAX1_5/a_46_6# 0 2.442f **FLOATING
C1706 FAX1_5/a_2_6# 0 2.5308f **FLOATING
C1707 FAX1_5/a_46_54# 0 4.1292f **FLOATING
C1708 FAX1_5/a_2_54# 0 4.3068f **FLOATING
C1709 FAX1_5/a_70_6# 0 6.54516f **FLOATING
C1710 FAX1_5/a_25_6# 0 9.36792f **FLOATING
C1711 BUFX2_7/a_2_6# 0 5.63946f **FLOATING
C1712 OAI21X1_109/a_2_6# 0 2.78652f **FLOATING
C1713 NOR2X1_80/Y 0 10.89264f **FLOATING
C1714 INVX2_58/A 0 46.64106f **FLOATING
C1715 FAX1_15/a_46_6# 0 2.442f **FLOATING
C1716 FAX1_15/a_2_6# 0 2.5308f **FLOATING
C1717 FAX1_15/a_46_54# 0 4.1292f **FLOATING
C1718 FAX1_15/a_2_54# 0 4.3068f **FLOATING
C1719 FAX1_15/a_70_6# 0 6.54516f **FLOATING
C1720 FAX1_15/a_25_6# 0 9.36792f **FLOATING
C1721 DFFNEGX1_7/a_66_6# 0 6.40992f **FLOATING
C1722 DFFNEGX1_7/a_23_6# 0 6.85692f **FLOATING
C1723 DFFNEGX1_7/a_34_4# 0 4.93023f **FLOATING
C1724 DFFNEGX1_7/a_2_6# 0 9.33504f **FLOATING
C1725 OAI22X1_77/a_2_6# 0 4.25172f **FLOATING
C1726 OAI22X1_88/a_2_6# 0 4.25172f **FLOATING
C1727 out_mines[20] 0 93.0717f **FLOATING
C1728 OAI22X1_44/a_2_6# 0 4.25172f **FLOATING
C1729 OAI22X1_55/a_2_6# 0 4.25172f **FLOATING
C1730 OAI22X1_66/a_2_6# 0 4.25172f **FLOATING
C1731 OAI22X1_33/a_2_6# 0 4.25172f **FLOATING
C1732 OAI22X1_11/a_2_6# 0 4.25172f **FLOATING
C1733 INVX2_96/Y 0 8.0085f **FLOATING
C1734 OAI22X1_22/a_2_6# 0 4.25172f **FLOATING
C1735 OAI21X1_9/a_2_6# 0 2.78652f **FLOATING
C1736 OR2X1_1/a_2_54# 0 6.27999f **FLOATING
C1737 HAX1_28/a_38_6# 0 2.442f **FLOATING
C1738 HAX1_28/a_41_74# 0 5.99325f **FLOATING
C1739 HAX1_28/a_2_74# 0 7.65318f **FLOATING
C1740 HAX1_17/a_38_6# 0 2.442f **FLOATING
C1741 HAX1_17/a_41_74# 0 5.99325f **FLOATING
C1742 HAX1_17/a_2_74# 0 7.65318f **FLOATING
C1743 HAX1_39/a_38_6# 0 2.442f **FLOATING
C1744 MUX2X1_5/A 0 8.10309f **FLOATING
C1745 HAX1_39/a_41_74# 0 5.99325f **FLOATING
C1746 HAX1_39/a_2_74# 0 7.65318f **FLOATING
C1747 AOI21X1_14/a_2_54# 0 4.3068f **FLOATING
C1748 AOI21X1_25/a_2_54# 0 4.3068f **FLOATING
C1749 AOI21X1_26/Y 0 13.274969f **FLOATING
C1750 BUFX2_24/a_2_6# 0 5.63946f **FLOATING
C1751 BUFX2_13/a_2_6# 0 5.63946f **FLOATING
C1752 AOI22X1_1/A 0 7.09215f **FLOATING
C1753 XNOR2X1_25/a_2_6# 0 6.77121f **FLOATING
C1754 XNOR2X1_25/a_12_41# 0 7.905991f **FLOATING
C1755 XNOR2X1_14/a_2_6# 0 6.77121f **FLOATING
C1756 XNOR2X1_14/a_12_41# 0 7.905991f **FLOATING
C1757 AOI21X1_6/a_2_54# 0 4.3068f **FLOATING
C1758 HAX1_46/B 0 14.95275f **FLOATING
C1759 AOI22X1_73/A 0 12.400081f **FLOATING
C1760 FAX1_4/a_46_6# 0 2.442f **FLOATING
C1761 FAX1_4/a_2_6# 0 2.5308f **FLOATING
C1762 FAX1_4/a_46_54# 0 4.1292f **FLOATING
C1763 FAX1_4/a_2_54# 0 4.3068f **FLOATING
C1764 FAX1_4/a_70_6# 0 6.54516f **FLOATING
C1765 FAX1_4/a_25_6# 0 9.36792f **FLOATING
C1766 BUFX2_6/a_2_6# 0 5.63946f **FLOATING
C1767 OAI21X1_119/a_2_6# 0 2.78652f **FLOATING
C1768 OAI21X1_108/a_2_6# 0 2.78652f **FLOATING
C1769 FAX1_14/a_46_6# 0 2.442f **FLOATING
C1770 FAX1_14/a_2_6# 0 2.5308f **FLOATING
C1771 FAX1_14/a_46_54# 0 4.1292f **FLOATING
C1772 FAX1_14/a_2_54# 0 4.3068f **FLOATING
C1773 FAX1_14/a_70_6# 0 6.54516f **FLOATING
C1774 FAX1_14/a_25_6# 0 9.36792f **FLOATING
C1775 out_temp_decoded[14] 0 13.01307f **FLOATING
C1776 INVX2_129/Y 0 11.273641f **FLOATING
C1777 out_temp_cleared[6] 0 12.311551f **FLOATING
C1778 DFFNEGX1_6/a_66_6# 0 6.40992f **FLOATING
C1779 DFFNEGX1_6/a_23_6# 0 6.85692f **FLOATING
C1780 DFFNEGX1_6/a_34_4# 0 4.93023f **FLOATING
C1781 DFFNEGX1_6/a_2_6# 0 9.33504f **FLOATING
C1782 INVX2_63/Y 0 31.05316f **FLOATING
C1783 OAI22X1_87/a_2_6# 0 4.25172f **FLOATING
C1784 OAI22X1_54/a_2_6# 0 4.25172f **FLOATING
C1785 OAI22X1_65/a_2_6# 0 4.25172f **FLOATING
C1786 OAI22X1_76/a_2_6# 0 4.25172f **FLOATING
C1787 OAI22X1_43/a_2_6# 0 4.25172f **FLOATING
C1788 OAI22X1_32/a_2_6# 0 4.25172f **FLOATING
C1789 OAI22X1_10/a_2_6# 0 4.25172f **FLOATING
C1790 OAI22X1_21/a_2_6# 0 4.25172f **FLOATING
C1791 OAI21X1_8/a_2_6# 0 2.78652f **FLOATING
C1792 OR2X1_0/a_2_54# 0 6.27999f **FLOATING
C1793 HAX1_49/a_38_6# 0 2.442f **FLOATING
C1794 HAX1_49/a_41_74# 0 5.99325f **FLOATING
C1795 HAX1_49/a_2_74# 0 7.65318f **FLOATING
C1796 HAX1_27/a_38_6# 0 2.442f **FLOATING
C1797 HAX1_27/a_41_74# 0 5.99325f **FLOATING
C1798 HAX1_27/a_2_74# 0 7.65318f **FLOATING
C1799 HAX1_16/a_38_6# 0 2.442f **FLOATING
C1800 HAX1_16/a_41_74# 0 5.99325f **FLOATING
C1801 HAX1_16/a_2_74# 0 7.65318f **FLOATING
C1802 HAX1_38/a_38_6# 0 2.442f **FLOATING
C1803 MUX2X1_6/A 0 8.10309f **FLOATING
C1804 HAX1_38/a_41_74# 0 5.99325f **FLOATING
C1805 HAX1_38/a_2_74# 0 7.65318f **FLOATING
C1806 AOI21X1_13/a_2_54# 0 4.3068f **FLOATING
C1807 AOI21X1_24/a_2_54# 0 4.3068f **FLOATING
C1808 NOR2X1_3/A 0 17.425138f **FLOATING
C1809 BUFX2_12/a_2_6# 0 5.63946f **FLOATING
C1810 BUFX2_23/a_2_6# 0 5.63946f **FLOATING
C1811 XNOR2X1_24/a_2_6# 0 6.77121f **FLOATING
C1812 XNOR2X1_24/a_12_41# 0 7.905991f **FLOATING
C1813 MUX2X1_2/A 0 10.764989f **FLOATING
C1814 XNOR2X1_13/a_2_6# 0 6.77121f **FLOATING
C1815 XNOR2X1_13/a_12_41# 0 7.905991f **FLOATING
C1816 AOI21X1_5/a_2_54# 0 4.3068f **FLOATING
C1817 NOR2X1_92/Y 0 6.77838f **FLOATING
C1818 AOI22X1_75/A 0 11.277359f **FLOATING
C1819 FAX1_3/a_46_6# 0 2.442f **FLOATING
C1820 FAX1_3/a_2_6# 0 2.5308f **FLOATING
C1821 FAX1_3/a_46_54# 0 4.1292f **FLOATING
C1822 FAX1_3/a_2_54# 0 4.3068f **FLOATING
C1823 FAX1_3/a_70_6# 0 6.54516f **FLOATING
C1824 FAX1_3/a_25_6# 0 9.36792f **FLOATING
C1825 in_incr[1] 0 6.02205f **FLOATING
C1826 BUFX2_5/a_2_6# 0 5.63946f **FLOATING
C1827 OAI21X1_118/a_2_6# 0 2.78652f **FLOATING
C1828 OAI21X1_118/Y 0 12.197461f **FLOATING
C1829 OAI21X1_107/a_2_6# 0 2.78652f **FLOATING
C1830 NAND2X1_96/Y 0 6.86169f **FLOATING
C1831 OAI21X1_129/a_2_6# 0 2.78652f **FLOATING
C1832 OAI21X1_93/C 0 11.02494f **FLOATING
C1833 FAX1_13/a_46_6# 0 2.442f **FLOATING
C1834 FAX1_13/a_2_6# 0 2.5308f **FLOATING
C1835 FAX1_13/a_46_54# 0 4.1292f **FLOATING
C1836 FAX1_13/a_2_54# 0 4.3068f **FLOATING
C1837 FAX1_13/a_70_6# 0 6.54516f **FLOATING
C1838 FAX1_13/a_25_6# 0 9.36792f **FLOATING
C1839 AOI21X1_16/Y 0 12.29553f **FLOATING
C1840 INVX2_76/A 0 8.41374f **FLOATING
C1841 NOR2X1_91/Y 0 29.622074f **FLOATING
C1842 DFFNEGX1_5/a_66_6# 0 6.40992f **FLOATING
C1843 DFFNEGX1_5/a_23_6# 0 6.85692f **FLOATING
C1844 DFFNEGX1_5/a_34_4# 0 4.93023f **FLOATING
C1845 DFFNEGX1_5/a_2_6# 0 9.33504f **FLOATING
C1846 OAI22X1_86/a_2_6# 0 4.25172f **FLOATING
C1847 OAI22X1_64/a_2_6# 0 4.25172f **FLOATING
C1848 OAI22X1_53/a_2_6# 0 4.25172f **FLOATING
C1849 OAI22X1_75/a_2_6# 0 4.25172f **FLOATING
C1850 OAI22X1_31/a_2_6# 0 4.25172f **FLOATING
C1851 OAI22X1_20/a_2_6# 0 4.25172f **FLOATING
C1852 OAI22X1_42/a_2_6# 0 4.25172f **FLOATING
C1853 OAI21X1_7/a_2_6# 0 2.78652f **FLOATING
C1854 HAX1_37/a_38_6# 0 2.442f **FLOATING
C1855 HAX1_37/a_41_74# 0 5.99325f **FLOATING
C1856 HAX1_37/a_2_74# 0 7.65318f **FLOATING
C1857 HAX1_26/a_38_6# 0 2.442f **FLOATING
C1858 HAX1_26/a_41_74# 0 5.99325f **FLOATING
C1859 HAX1_26/a_2_74# 0 7.65318f **FLOATING
C1860 HAX1_48/a_38_6# 0 2.442f **FLOATING
C1861 HAX1_49/B 0 12.947281f **FLOATING
C1862 HAX1_48/a_41_74# 0 5.99325f **FLOATING
C1863 HAX1_48/a_2_74# 0 7.65318f **FLOATING
C1864 HAX1_15/a_38_6# 0 2.442f **FLOATING
C1865 HAX1_15/a_41_74# 0 5.99325f **FLOATING
C1866 HAX1_15/a_2_74# 0 7.65318f **FLOATING
C1867 AOI21X1_23/a_2_54# 0 4.3068f **FLOATING
C1868 AOI21X1_12/a_2_54# 0 4.3068f **FLOATING
C1869 NOR2X1_2/Y 0 12.198901f **FLOATING
C1870 BUFX2_22/a_2_6# 0 5.63946f **FLOATING
C1871 BUFX2_11/a_2_6# 0 5.63946f **FLOATING
C1872 XNOR2X1_23/Y 0 8.247869f **FLOATING
C1873 XNOR2X1_23/a_2_6# 0 6.77121f **FLOATING
C1874 XNOR2X1_23/a_12_41# 0 7.905991f **FLOATING
C1875 MUX2X1_3/A 0 11.607269f **FLOATING
C1876 XNOR2X1_12/a_2_6# 0 6.77121f **FLOATING
C1877 XNOR2X1_12/a_12_41# 0 7.905991f **FLOATING
C1878 AOI21X1_4/a_2_54# 0 4.3068f **FLOATING
C1879 INVX2_107/Y 0 18.84034f **FLOATING
C1880 INVX2_101/Y 0 7.67754f **FLOATING
C1881 OAI22X1_76/B 0 34.611176f **FLOATING
C1882 BUFX2_17/Y 0 0.176059p **FLOATING
C1883 FAX1_2/a_46_6# 0 2.442f **FLOATING
C1884 FAX1_2/a_2_6# 0 2.5308f **FLOATING
C1885 FAX1_2/a_46_54# 0 4.1292f **FLOATING
C1886 FAX1_2/a_2_54# 0 4.3068f **FLOATING
C1887 FAX1_2/a_70_6# 0 6.54516f **FLOATING
C1888 FAX1_2/a_25_6# 0 9.36792f **FLOATING
C1889 in_incr[2] 0 6.02205f **FLOATING
C1890 BUFX2_4/a_2_6# 0 5.63946f **FLOATING
C1891 OAI21X1_139/a_2_6# 0 2.78652f **FLOATING
C1892 OAI21X1_117/a_2_6# 0 2.78652f **FLOATING
C1893 INVX2_50/A 0 13.522079f **FLOATING
C1894 OAI21X1_106/a_2_6# 0 2.78652f **FLOATING
C1895 NAND2X1_93/Y 0 6.86169f **FLOATING
C1896 OAI21X1_128/a_2_6# 0 2.78652f **FLOATING
C1897 FAX1_12/a_46_6# 0 2.442f **FLOATING
C1898 FAX1_12/a_2_6# 0 2.5308f **FLOATING
C1899 FAX1_12/a_46_54# 0 4.1292f **FLOATING
C1900 FAX1_12/a_2_54# 0 4.3068f **FLOATING
C1901 FAX1_12/a_70_6# 0 6.54516f **FLOATING
C1902 FAX1_12/a_25_6# 0 9.36792f **FLOATING
C1903 OAI22X1_56/Y 0 8.24718f **FLOATING
C1904 HAX1_38/A 0 21.094738f **FLOATING
C1905 OAI21X1_69/C 0 8.869499f **FLOATING
C1906 XOR2X1_9/a_2_6# 0 8.278139f **FLOATING
C1907 XOR2X1_9/a_13_43# 0 7.836241f **FLOATING
C1908 DFFNEGX1_4/a_66_6# 0 6.40992f **FLOATING
C1909 DFFNEGX1_4/a_23_6# 0 6.85692f **FLOATING
C1910 DFFNEGX1_4/a_34_4# 0 4.93023f **FLOATING
C1911 DFFNEGX1_4/a_2_6# 0 9.33504f **FLOATING
C1912 OAI22X1_63/a_2_6# 0 4.25172f **FLOATING
C1913 OAI22X1_85/a_2_6# 0 4.25172f **FLOATING
C1914 OAI22X1_74/a_2_6# 0 4.25172f **FLOATING
C1915 OAI22X1_30/a_2_6# 0 4.25172f **FLOATING
C1916 OAI22X1_41/a_2_6# 0 4.25172f **FLOATING
C1917 OAI22X1_52/a_2_6# 0 4.25172f **FLOATING
C1918 OAI21X1_6/a_2_6# 0 2.78652f **FLOATING
C1919 HAX1_36/a_38_6# 0 2.442f **FLOATING
C1920 HAX1_36/YS 0 7.40268f **FLOATING
C1921 HAX1_36/a_41_74# 0 5.99325f **FLOATING
C1922 HAX1_36/a_2_74# 0 7.65318f **FLOATING
C1923 HAX1_25/a_38_6# 0 2.442f **FLOATING
C1924 HAX1_25/a_41_74# 0 5.99325f **FLOATING
C1925 HAX1_25/a_2_74# 0 7.65318f **FLOATING
C1926 HAX1_47/a_38_6# 0 2.442f **FLOATING
C1927 HAX1_47/YS 0 8.10309f **FLOATING
C1928 HAX1_47/a_41_74# 0 5.99325f **FLOATING
C1929 HAX1_47/a_2_74# 0 7.65318f **FLOATING
C1930 AOI21X1_11/Y 0 7.18191f **FLOATING
C1931 AOI21X1_11/a_2_54# 0 4.3068f **FLOATING
C1932 AOI21X1_22/a_2_54# 0 4.3068f **FLOATING
C1933 HAX1_14/a_38_6# 0 2.442f **FLOATING
C1934 HAX1_14/YS 0 6.99546f **FLOATING
C1935 HAX1_14/a_41_74# 0 5.99325f **FLOATING
C1936 HAX1_14/a_2_74# 0 7.65318f **FLOATING
C1937 BUFX2_21/a_2_6# 0 5.63946f **FLOATING
C1938 BUFX2_10/a_2_6# 0 5.63946f **FLOATING
C1939 XNOR2X1_22/a_2_6# 0 6.77121f **FLOATING
C1940 XNOR2X1_22/a_12_41# 0 7.905991f **FLOATING
C1941 MUX2X1_7/A 0 10.543229f **FLOATING
C1942 XNOR2X1_11/a_2_6# 0 6.77121f **FLOATING
C1943 XNOR2X1_11/a_12_41# 0 7.905991f **FLOATING
C1944 AOI21X1_3/Y 0 8.65788f **FLOATING
C1945 AOI21X1_3/a_2_54# 0 4.3068f **FLOATING
C1946 FAX1_1/a_46_6# 0 2.442f **FLOATING
C1947 FAX1_1/a_2_6# 0 2.5308f **FLOATING
C1948 FAX1_1/a_46_54# 0 4.1292f **FLOATING
C1949 FAX1_1/a_2_54# 0 4.3068f **FLOATING
C1950 FAX1_1/a_70_6# 0 6.54516f **FLOATING
C1951 FAX1_1/a_25_6# 0 9.36792f **FLOATING
C1952 in_incr[3] 0 6.02205f **FLOATING
C1953 BUFX2_3/a_2_6# 0 5.63946f **FLOATING
C1954 OAI21X1_149/a_2_6# 0 2.78652f **FLOATING
C1955 OAI21X1_138/a_2_6# 0 2.78652f **FLOATING
C1956 OAI21X1_116/a_2_6# 0 2.78652f **FLOATING
C1957 OAI22X1_40/Y 0 9.911041f **FLOATING
C1958 NOR2X1_109/Y 0 9.616139f **FLOATING
C1959 OAI21X1_105/a_2_6# 0 2.78652f **FLOATING
C1960 NAND2X1_92/Y 0 10.81764f **FLOATING
C1961 OAI21X1_127/a_2_6# 0 2.78652f **FLOATING
C1962 AOI21X1_12/B 0 7.33464f **FLOATING
C1963 INVX2_52/Y 0 18.277441f **FLOATING
C1964 XOR2X1_19/Y 0 12.84477f **FLOATING
C1965 XOR2X1_19/a_2_6# 0 8.278139f **FLOATING
C1966 XOR2X1_19/a_13_43# 0 7.836241f **FLOATING
C1967 INVX2_40/Y 0 23.014063f **FLOATING
C1968 NOR2X1_51/Y 0 10.612081f **FLOATING
C1969 FAX1_11/a_46_6# 0 2.442f **FLOATING
C1970 FAX1_11/a_2_6# 0 2.5308f **FLOATING
C1971 FAX1_11/a_46_54# 0 4.1292f **FLOATING
C1972 FAX1_11/a_2_54# 0 4.3068f **FLOATING
C1973 FAX1_11/a_70_6# 0 6.54516f **FLOATING
C1974 FAX1_11/a_25_6# 0 9.36792f **FLOATING
C1975 HAX1_39/A 0 18.769289f **FLOATING
C1976 OR2X1_16/A 0 9.381721f **FLOATING
C1977 AND2X2_11/Y 0 12.49959f **FLOATING
C1978 NAND2X1_63/B 0 13.20522f **FLOATING
C1979 MUX2X1_9/Y 0 9.89586f **FLOATING
C1980 MUX2X1_9/A 0 6.13938f **FLOATING
C1981 MUX2X1_9/a_2_10# 0 6.0456f **FLOATING
C1982 XOR2X1_8/a_2_6# 0 8.278139f **FLOATING
C1983 XOR2X1_8/a_13_43# 0 7.836241f **FLOATING
C1984 DFFNEGX1_3/a_66_6# 0 6.40992f **FLOATING
C1985 DFFNEGX1_3/a_23_6# 0 6.85692f **FLOATING
C1986 DFFNEGX1_3/a_34_4# 0 4.93023f **FLOATING
C1987 DFFNEGX1_3/a_2_6# 0 9.33504f **FLOATING
C1988 INVX2_65/Y 0 28.982275f **FLOATING
C1989 OAI22X1_62/a_2_6# 0 4.25172f **FLOATING
C1990 OAI22X1_84/a_2_6# 0 4.25172f **FLOATING
C1991 OAI22X1_73/a_2_6# 0 4.25172f **FLOATING
C1992 OAI22X1_40/a_2_6# 0 4.25172f **FLOATING
C1993 OAI22X1_51/a_2_6# 0 4.25172f **FLOATING
C1994 OAI21X1_5/a_2_6# 0 2.78652f **FLOATING
C1995 HAX1_35/a_38_6# 0 2.442f **FLOATING
C1996 HAX1_35/YS 0 8.247f **FLOATING
C1997 HAX1_35/a_41_74# 0 5.99325f **FLOATING
C1998 HAX1_35/a_2_74# 0 7.65318f **FLOATING
C1999 HAX1_24/a_38_6# 0 2.442f **FLOATING
C2000 HAX1_23/B 0 13.55931f **FLOATING
C2001 HAX1_24/a_41_74# 0 5.99325f **FLOATING
C2002 HAX1_24/a_2_74# 0 7.65318f **FLOATING
C2003 HAX1_46/a_38_6# 0 2.442f **FLOATING
C2004 HAX1_46/a_41_74# 0 5.99325f **FLOATING
C2005 HAX1_46/a_2_74# 0 7.65318f **FLOATING
C2006 AOI21X1_21/a_2_54# 0 4.3068f **FLOATING
C2007 HAX1_13/a_38_6# 0 2.442f **FLOATING
C2008 HAX1_12/B 0 12.215281f **FLOATING
C2009 HAX1_13/a_41_74# 0 5.99325f **FLOATING
C2010 HAX1_13/a_2_74# 0 7.65318f **FLOATING
C2011 AOI21X1_10/a_2_54# 0 4.3068f **FLOATING
C2012 BUFX2_20/a_2_6# 0 5.63946f **FLOATING
C2013 XNOR2X1_21/a_2_6# 0 6.77121f **FLOATING
C2014 XNOR2X1_21/a_12_41# 0 7.905991f **FLOATING
C2015 MUX2X1_8/A 0 11.525189f **FLOATING
C2016 XNOR2X1_10/a_2_6# 0 6.77121f **FLOATING
C2017 XNOR2X1_10/a_12_41# 0 7.905991f **FLOATING
C2018 INVX2_218/A 0 6.53484f **FLOATING
C2019 AOI21X1_2/a_2_54# 0 4.3068f **FLOATING
C2020 INVX2_99/Y 0 10.78374f **FLOATING
C2021 out_temp_index[1] 0 15.579152f **FLOATING
C2022 FAX1_0/a_46_6# 0 2.442f **FLOATING
C2023 FAX1_0/a_2_6# 0 2.5308f **FLOATING
C2024 FAX1_0/a_46_54# 0 4.1292f **FLOATING
C2025 FAX1_0/a_2_54# 0 4.3068f **FLOATING
C2026 FAX1_0/a_70_6# 0 6.54516f **FLOATING
C2027 FAX1_0/a_25_6# 0 9.36792f **FLOATING
C2028 in_incr[4] 0 6.02205f **FLOATING
C2029 OAI22X1_51/D 0 39.06087f **FLOATING
C2030 BUFX2_2/a_2_6# 0 5.63946f **FLOATING
C2031 OAI21X1_148/a_2_6# 0 2.78652f **FLOATING
C2032 OAI21X1_159/a_2_6# 0 2.78652f **FLOATING
C2033 OAI21X1_126/a_2_6# 0 2.78652f **FLOATING
C2034 AOI21X1_11/A 0 7.4559f **FLOATING
C2035 OAI21X1_115/a_2_6# 0 2.78652f **FLOATING
C2036 INVX2_43/A 0 14.651371f **FLOATING
C2037 OAI21X1_137/a_2_6# 0 2.78652f **FLOATING
C2038 OAI21X1_104/a_2_6# 0 2.78652f **FLOATING
C2039 NOR2X1_63/Y 0 8.522281f **FLOATING
C2040 XOR2X1_29/Y 0 16.277882f **FLOATING
C2041 XOR2X1_29/a_2_6# 0 8.278139f **FLOATING
C2042 XOR2X1_29/a_13_43# 0 7.836241f **FLOATING
C2043 NOR2X1_43/Y 0 14.61706f **FLOATING
C2044 XOR2X1_18/a_2_6# 0 8.278139f **FLOATING
C2045 XOR2X1_18/a_13_43# 0 7.836241f **FLOATING
C2046 FAX1_10/a_46_6# 0 2.442f **FLOATING
C2047 FAX1_10/a_2_6# 0 2.5308f **FLOATING
C2048 FAX1_10/a_46_54# 0 4.1292f **FLOATING
C2049 FAX1_10/a_2_54# 0 4.3068f **FLOATING
C2050 FAX1_10/a_70_6# 0 6.54516f **FLOATING
C2051 FAX1_10/a_25_6# 0 9.36792f **FLOATING
C2052 MUX2X1_8/a_2_10# 0 6.0456f **FLOATING
C2053 XOR2X1_7/a_2_6# 0 8.278139f **FLOATING
C2054 XOR2X1_7/a_13_43# 0 7.836241f **FLOATING
C2055 DFFNEGX1_2/a_66_6# 0 6.40992f **FLOATING
C2056 DFFNEGX1_2/a_23_6# 0 6.85692f **FLOATING
C2057 DFFNEGX1_2/a_34_4# 0 4.93023f **FLOATING
C2058 DFFNEGX1_2/a_2_6# 0 9.33504f **FLOATING
C2059 INVX2_55/Y 0 12.94968f **FLOATING
C2060 OAI22X1_83/a_2_6# 0 4.25172f **FLOATING
C2061 OAI22X1_72/a_2_6# 0 4.25172f **FLOATING
C2062 OAI22X1_61/a_2_6# 0 4.25172f **FLOATING
C2063 OAI22X1_63/B 0 35.285812f **FLOATING
C2064 OAI22X1_50/a_2_6# 0 4.25172f **FLOATING
C2065 OAI21X1_4/a_2_6# 0 2.78652f **FLOATING
C2066 HAX1_34/a_38_6# 0 2.442f **FLOATING
C2067 HAX1_34/a_41_74# 0 5.99325f **FLOATING
C2068 HAX1_34/a_2_74# 0 7.65318f **FLOATING
C2069 HAX1_45/a_38_6# 0 2.442f **FLOATING
C2070 HAX1_45/a_41_74# 0 5.99325f **FLOATING
C2071 HAX1_45/a_2_74# 0 7.65318f **FLOATING
C2072 AOI21X1_20/a_2_54# 0 4.3068f **FLOATING
C2073 HAX1_23/a_38_6# 0 2.442f **FLOATING
C2074 HAX1_23/a_41_74# 0 5.99325f **FLOATING
C2075 HAX1_23/a_2_74# 0 7.65318f **FLOATING
C2076 HAX1_12/a_38_6# 0 2.442f **FLOATING
C2077 HAX1_12/a_41_74# 0 5.99325f **FLOATING
C2078 HAX1_12/a_2_74# 0 7.65318f **FLOATING
C2079 out_global_score[18] 0 19.270409f **FLOATING
C2080 XNOR2X1_20/a_2_6# 0 6.77121f **FLOATING
C2081 XNOR2X1_20/a_12_41# 0 7.905991f **FLOATING
C2082 INVX2_245/A 0 6.54867f **FLOATING
C2083 AOI21X1_1/a_2_54# 0 4.3068f **FLOATING
C2084 INVX2_1/Y 0 38.82282f **FLOATING
C2085 BUFX2_1/a_2_6# 0 5.63946f **FLOATING
C2086 OAI21X1_158/a_2_6# 0 2.78652f **FLOATING
C2087 OAI21X1_136/a_2_6# 0 2.78652f **FLOATING
C2088 OAI21X1_147/a_2_6# 0 2.78652f **FLOATING
C2089 OAI21X1_114/a_2_6# 0 2.78652f **FLOATING
C2090 OAI21X1_125/a_2_6# 0 2.78652f **FLOATING
C2091 OAI21X1_103/a_2_6# 0 2.78652f **FLOATING
C2092 DFFNEGX1_109/a_66_6# 0 6.40992f **FLOATING
C2093 DFFNEGX1_109/a_23_6# 0 6.85692f **FLOATING
C2094 DFFNEGX1_109/a_34_4# 0 4.93023f **FLOATING
C2095 DFFNEGX1_109/a_2_6# 0 9.33504f **FLOATING
C2096 XOR2X1_28/Y 0 15.35805f **FLOATING
C2097 XOR2X1_28/a_2_6# 0 8.278139f **FLOATING
C2098 XOR2X1_28/a_13_43# 0 7.836241f **FLOATING
C2099 XOR2X1_17/a_2_6# 0 8.278139f **FLOATING
C2100 XOR2X1_17/a_13_43# 0 7.836241f **FLOATING
C2101 NOR2X1_42/Y 0 9.14616f **FLOATING
C2102 DFFNEGX1_19/a_66_6# 0 6.40992f **FLOATING
C2103 DFFNEGX1_19/a_23_6# 0 6.85692f **FLOATING
C2104 DFFNEGX1_19/a_34_4# 0 4.93023f **FLOATING
C2105 DFFNEGX1_19/a_2_6# 0 9.33504f **FLOATING
C2106 INVX2_179/Y 0 9.24252f **FLOATING
C2107 OR2X1_3/A 0 8.47428f **FLOATING
C2108 INVX2_124/A 0 17.16477f **FLOATING
C2109 OAI21X1_74/C 0 9.4167f **FLOATING
C2110 OAI22X1_14/Y 0 9.9711f **FLOATING
C2111 MUX2X1_7/a_2_10# 0 6.0456f **FLOATING
C2112 XOR2X1_6/a_2_6# 0 8.278139f **FLOATING
C2113 XOR2X1_6/a_13_43# 0 7.836241f **FLOATING
C2114 DFFNEGX1_1/a_66_6# 0 6.40992f **FLOATING
C2115 DFFNEGX1_1/a_23_6# 0 6.85692f **FLOATING
C2116 DFFNEGX1_1/a_34_4# 0 4.93023f **FLOATING
C2117 DFFNEGX1_1/a_2_6# 0 9.33504f **FLOATING
C2118 OAI22X1_82/a_2_6# 0 4.25172f **FLOATING
C2119 OAI22X1_71/a_2_6# 0 4.25172f **FLOATING
C2120 OAI22X1_60/a_2_6# 0 4.25172f **FLOATING
C2121 OAI21X1_3/a_2_6# 0 2.78652f **FLOATING
C2122 HAX1_33/a_38_6# 0 2.442f **FLOATING
C2123 HAX1_33/a_41_74# 0 5.99325f **FLOATING
C2124 HAX1_33/a_2_74# 0 7.65318f **FLOATING
C2125 HAX1_44/a_38_6# 0 2.442f **FLOATING
C2126 HAX1_44/a_41_74# 0 5.99325f **FLOATING
C2127 HAX1_44/a_2_74# 0 7.65318f **FLOATING
C2128 HAX1_11/a_38_6# 0 2.442f **FLOATING
C2129 HAX1_11/a_41_74# 0 5.99325f **FLOATING
C2130 HAX1_11/a_2_74# 0 7.65318f **FLOATING
C2131 HAX1_11/B 0 13.37475f **FLOATING
C2132 HAX1_22/a_38_6# 0 2.442f **FLOATING
C2133 HAX1_22/a_41_74# 0 5.99325f **FLOATING
C2134 HAX1_22/a_2_74# 0 7.65318f **FLOATING
C2135 XNOR2X1_30/a_2_6# 0 6.77121f **FLOATING
C2136 XNOR2X1_30/a_12_41# 0 7.905991f **FLOATING
C2137 AOI21X1_0/a_2_54# 0 4.3068f **FLOATING
C2138 OAI21X1_0/A 0 16.80111f **FLOATING
C2139 AOI22X1_19/a_2_54# 0 6.66f **FLOATING
C2140 out_global_score[14] 0 19.335508f **FLOATING
C2141 INVX2_117/Y 0 37.60511f **FLOATING
C2142 BUFX2_0/a_2_6# 0 5.63946f **FLOATING
C2143 OAI21X1_157/a_2_6# 0 2.78652f **FLOATING
C2144 OAI21X1_157/B 0 6.4515f **FLOATING
C2145 OAI21X1_124/a_2_6# 0 2.78652f **FLOATING
C2146 OAI21X1_124/Y 0 9.92004f **FLOATING
C2147 OAI21X1_135/a_2_6# 0 2.78652f **FLOATING
C2148 OAI21X1_146/a_2_6# 0 2.78652f **FLOATING
C2149 OAI21X1_113/a_2_6# 0 2.78652f **FLOATING
C2150 OAI21X1_102/a_2_6# 0 2.78652f **FLOATING
C2151 DFFNEGX1_119/a_66_6# 0 6.40992f **FLOATING
C2152 DFFNEGX1_119/a_23_6# 0 6.85692f **FLOATING
C2153 DFFNEGX1_119/a_34_4# 0 4.93023f **FLOATING
C2154 DFFNEGX1_119/a_2_6# 0 9.33504f **FLOATING
C2155 INVX2_191/Y 0 10.468379f **FLOATING
C2156 NAND3X1_6/Y 0 8.276759f **FLOATING
C2157 DFFNEGX1_108/a_66_6# 0 6.40992f **FLOATING
C2158 DFFNEGX1_108/a_23_6# 0 6.85692f **FLOATING
C2159 DFFNEGX1_108/a_34_4# 0 4.93023f **FLOATING
C2160 DFFNEGX1_108/a_2_6# 0 9.33504f **FLOATING
C2161 XOR2X1_27/a_2_6# 0 8.278139f **FLOATING
C2162 XOR2X1_27/a_13_43# 0 7.836241f **FLOATING
C2163 XOR2X1_16/Y 0 17.176739f **FLOATING
C2164 XOR2X1_16/a_2_6# 0 8.278139f **FLOATING
C2165 XOR2X1_16/a_13_43# 0 7.836241f **FLOATING
C2166 DFFNEGX1_29/a_66_6# 0 6.40992f **FLOATING
C2167 DFFNEGX1_29/a_23_6# 0 6.85692f **FLOATING
C2168 DFFNEGX1_29/a_34_4# 0 4.93023f **FLOATING
C2169 DFFNEGX1_29/a_2_6# 0 9.33504f **FLOATING
C2170 OAI21X1_45/Y 0 10.456441f **FLOATING
C2171 DFFNEGX1_18/a_66_6# 0 6.40992f **FLOATING
C2172 DFFNEGX1_18/a_23_6# 0 6.85692f **FLOATING
C2173 DFFNEGX1_18/a_34_4# 0 4.93023f **FLOATING
C2174 DFFNEGX1_18/a_2_6# 0 9.33504f **FLOATING
C2175 INVX2_243/Y 0 18.30606f **FLOATING
C2176 OR2X1_1/A 0 8.47428f **FLOATING
C2177 out_temp_cleared[1] 0 11.899351f **FLOATING
C2178 OAI21X1_73/C 0 11.68416f **FLOATING
C2179 NOR2X1_84/Y 0 11.236442f **FLOATING
C2180 OAI21X1_88/Y 0 13.05648f **FLOATING
C2181 MUX2X1_6/Y 0 6.36198f **FLOATING
C2182 MUX2X1_6/a_2_10# 0 6.0456f **FLOATING
C2183 XOR2X1_5/Y 0 19.305897f **FLOATING
C2184 XOR2X1_5/a_2_6# 0 8.278139f **FLOATING
C2185 XOR2X1_5/a_13_43# 0 7.836241f **FLOATING
C2186 out_mines[14] 0 0.117649p **FLOATING
C2187 DFFNEGX1_0/a_66_6# 0 6.40992f **FLOATING
C2188 DFFNEGX1_0/a_23_6# 0 6.85692f **FLOATING
C2189 DFFNEGX1_0/a_34_4# 0 4.93023f **FLOATING
C2190 DFFNEGX1_0/a_2_6# 0 9.33504f **FLOATING
C2191 OAI22X1_81/a_2_6# 0 4.25172f **FLOATING
C2192 OAI22X1_70/a_2_6# 0 4.25172f **FLOATING
C2193 OAI21X1_2/a_2_6# 0 2.78652f **FLOATING
C2194 OAI21X1_2/Y 0 8.56716f **FLOATING
C2195 HAX1_43/a_38_6# 0 2.442f **FLOATING
C2196 HAX1_43/YS 0 8.10309f **FLOATING
C2197 HAX1_43/a_41_74# 0 5.99325f **FLOATING
C2198 HAX1_43/a_2_74# 0 7.65318f **FLOATING
C2199 HAX1_10/a_38_6# 0 2.442f **FLOATING
C2200 HAX1_10/YS 0 6.99546f **FLOATING
C2201 HAX1_10/a_41_74# 0 5.99325f **FLOATING
C2202 HAX1_10/a_2_74# 0 7.65318f **FLOATING
C2203 HAX1_32/a_38_6# 0 2.442f **FLOATING
C2204 HAX1_32/a_41_74# 0 5.99325f **FLOATING
C2205 HAX1_32/a_2_74# 0 7.65318f **FLOATING
C2206 HAX1_21/a_38_6# 0 2.442f **FLOATING
C2207 HAX1_20/B 0 11.520601f **FLOATING
C2208 HAX1_21/a_41_74# 0 5.99325f **FLOATING
C2209 HAX1_21/a_2_74# 0 7.65318f **FLOATING
C2210 AOI22X1_29/a_2_54# 0 6.66f **FLOATING
C2211 AOI22X1_18/a_2_54# 0 6.66f **FLOATING
C2212 HAX1_15/YS 0 7.00383f **FLOATING
C2213 OAI21X1_4/A 0 34.205532f **FLOATING
C2214 OAI21X1_123/a_2_6# 0 2.78652f **FLOATING
C2215 OAI21X1_134/a_2_6# 0 2.78652f **FLOATING
C2216 OAI21X1_156/a_2_6# 0 2.78652f **FLOATING
C2217 OAI21X1_145/a_2_6# 0 2.78652f **FLOATING
C2218 OAI21X1_112/a_2_6# 0 2.78652f **FLOATING
C2219 AOI22X1_54/B 0 11.84886f **FLOATING
C2220 OAI21X1_101/a_2_6# 0 2.78652f **FLOATING
C2221 DFFNEGX1_129/a_66_6# 0 6.40992f **FLOATING
C2222 DFFNEGX1_129/a_23_6# 0 6.85692f **FLOATING
C2223 DFFNEGX1_129/a_34_4# 0 4.93023f **FLOATING
C2224 DFFNEGX1_129/a_2_6# 0 9.33504f **FLOATING
C2225 DFFNEGX1_118/a_66_6# 0 6.40992f **FLOATING
C2226 DFFNEGX1_118/a_23_6# 0 6.85692f **FLOATING
C2227 DFFNEGX1_118/a_34_4# 0 4.93023f **FLOATING
C2228 DFFNEGX1_118/a_2_6# 0 9.33504f **FLOATING
C2229 DFFNEGX1_107/a_66_6# 0 6.40992f **FLOATING
C2230 DFFNEGX1_107/a_23_6# 0 6.85692f **FLOATING
C2231 DFFNEGX1_107/a_34_4# 0 4.93023f **FLOATING
C2232 DFFNEGX1_107/a_2_6# 0 9.33504f **FLOATING
C2233 XOR2X1_26/a_2_6# 0 8.278139f **FLOATING
C2234 XOR2X1_26/a_13_43# 0 7.836241f **FLOATING
C2235 XOR2X1_15/Y 0 8.300611f **FLOATING
C2236 XOR2X1_15/a_2_6# 0 8.278139f **FLOATING
C2237 XOR2X1_15/a_13_43# 0 7.836241f **FLOATING
C2238 DFFNEGX1_39/a_66_6# 0 6.40992f **FLOATING
C2239 DFFNEGX1_39/a_23_6# 0 6.85692f **FLOATING
C2240 DFFNEGX1_39/a_34_4# 0 4.93023f **FLOATING
C2241 DFFNEGX1_39/a_2_6# 0 9.33504f **FLOATING
C2242 OAI21X1_109/Y 0 12.32802f **FLOATING
C2243 DFFNEGX1_28/a_66_6# 0 6.40992f **FLOATING
C2244 DFFNEGX1_28/a_23_6# 0 6.85692f **FLOATING
C2245 DFFNEGX1_28/a_34_4# 0 4.93023f **FLOATING
C2246 DFFNEGX1_28/a_2_6# 0 9.33504f **FLOATING
C2247 DFFNEGX1_17/a_66_6# 0 6.40992f **FLOATING
C2248 DFFNEGX1_17/a_23_6# 0 6.85692f **FLOATING
C2249 DFFNEGX1_17/a_34_4# 0 4.93023f **FLOATING
C2250 DFFNEGX1_17/a_2_6# 0 9.33504f **FLOATING
C2251 AOI21X1_14/B 0 9.1689f **FLOATING
C2252 NOR2X1_64/B 0 8.653501f **FLOATING
C2253 INVX2_199/Y 0 11.78586f **FLOATING
C2254 INVX2_199/A 0 11.234819f **FLOATING
C2255 HAX1_40/A 0 19.924139f **FLOATING
C2256 INVX2_122/Y 0 7.11246f **FLOATING
C2257 INVX2_100/Y 0 5.84082f **FLOATING
C2258 OAI21X1_82/Y 0 10.50996f **FLOATING
C2259 OAI21X1_93/Y 0 11.123521f **FLOATING
C2260 NOR2X1_85/A 0 11.121961f **FLOATING
C2261 NOR2X1_84/A 0 24.507868f **FLOATING
C2262 MUX2X1_5/a_2_10# 0 6.0456f **FLOATING
C2263 XOR2X1_4/Y 0 26.854088f **FLOATING
C2264 XOR2X1_4/a_2_6# 0 8.278139f **FLOATING
C2265 XOR2X1_4/a_13_43# 0 7.836241f **FLOATING
C2266 OAI22X1_80/a_2_6# 0 4.25172f **FLOATING
C2267 OAI21X1_1/a_2_6# 0 2.78652f **FLOATING
C2268 AND2X2_6/B 0 10.14165f **FLOATING
C2269 HAX1_31/a_38_6# 0 2.442f **FLOATING
C2270 FAX1_14/A 0 17.60424f **FLOATING
C2271 HAX1_31/a_41_74# 0 5.99325f **FLOATING
C2272 HAX1_31/a_2_74# 0 7.65318f **FLOATING
C2273 HAX1_42/a_38_6# 0 2.442f **FLOATING
C2274 HAX1_42/YS 0 7.77249f **FLOATING
C2275 HAX1_42/a_41_74# 0 5.99325f **FLOATING
C2276 HAX1_42/a_2_74# 0 7.65318f **FLOATING
C2277 HAX1_20/a_38_6# 0 2.442f **FLOATING
C2278 HAX1_20/YS 0 6.99546f **FLOATING
C2279 HAX1_20/a_41_74# 0 5.99325f **FLOATING
C2280 HAX1_20/a_2_74# 0 7.65318f **FLOATING
C2281 out_n_nearby[1] 0 11.525549f **FLOATING
C2282 AOI22X1_39/a_2_54# 0 6.66f **FLOATING
C2283 AOI22X1_28/a_2_54# 0 6.66f **FLOATING
C2284 out_global_score[5] 0 16.232399f **FLOATING
C2285 AOI22X1_17/a_2_54# 0 6.66f **FLOATING
C2286 INVX2_234/Y 0 12.08631f **FLOATING
C2287 OAI21X1_133/a_2_6# 0 2.78652f **FLOATING
C2288 OAI21X1_155/a_2_6# 0 2.78652f **FLOATING
C2289 OAI21X1_144/a_2_6# 0 2.78652f **FLOATING
C2290 AOI22X1_9/a_2_54# 0 6.66f **FLOATING
C2291 OAI21X1_111/a_2_6# 0 2.78652f **FLOATING
C2292 OAI21X1_111/C 0 6.86169f **FLOATING
C2293 OAI21X1_122/a_2_6# 0 2.78652f **FLOATING
C2294 OAI21X1_100/a_2_6# 0 2.78652f **FLOATING
C2295 DFFNEGX1_128/a_66_6# 0 6.40992f **FLOATING
C2296 DFFNEGX1_128/a_23_6# 0 6.85692f **FLOATING
C2297 DFFNEGX1_128/a_34_4# 0 4.93023f **FLOATING
C2298 DFFNEGX1_128/a_2_6# 0 9.33504f **FLOATING
C2299 DFFNEGX1_139/a_66_6# 0 6.40992f **FLOATING
C2300 DFFNEGX1_139/a_23_6# 0 6.85692f **FLOATING
C2301 DFFNEGX1_139/a_34_4# 0 4.93023f **FLOATING
C2302 DFFNEGX1_139/a_2_6# 0 9.33504f **FLOATING
C2303 DFFNEGX1_117/a_66_6# 0 6.40992f **FLOATING
C2304 DFFNEGX1_117/a_23_6# 0 6.85692f **FLOATING
C2305 DFFNEGX1_117/a_34_4# 0 4.93023f **FLOATING
C2306 DFFNEGX1_117/a_2_6# 0 9.33504f **FLOATING
C2307 DFFNEGX1_106/a_66_6# 0 6.40992f **FLOATING
C2308 DFFNEGX1_106/a_23_6# 0 6.85692f **FLOATING
C2309 DFFNEGX1_106/a_34_4# 0 4.93023f **FLOATING
C2310 DFFNEGX1_106/a_2_6# 0 9.33504f **FLOATING
C2311 XOR2X1_25/a_2_6# 0 8.278139f **FLOATING
C2312 XOR2X1_25/a_13_43# 0 7.836241f **FLOATING
C2313 XOR2X1_14/a_2_6# 0 8.278139f **FLOATING
C2314 XOR2X1_14/a_13_43# 0 7.836241f **FLOATING
C2315 DFFNEGX1_38/a_66_6# 0 6.40992f **FLOATING
C2316 DFFNEGX1_38/a_23_6# 0 6.85692f **FLOATING
C2317 DFFNEGX1_38/a_34_4# 0 4.93023f **FLOATING
C2318 DFFNEGX1_38/a_2_6# 0 9.33504f **FLOATING
C2319 DFFNEGX1_49/a_66_6# 0 6.40992f **FLOATING
C2320 DFFNEGX1_49/a_23_6# 0 6.85692f **FLOATING
C2321 DFFNEGX1_49/a_34_4# 0 4.93023f **FLOATING
C2322 DFFNEGX1_49/a_2_6# 0 9.33504f **FLOATING
C2323 OAI21X1_99/Y 0 12.263939f **FLOATING
C2324 DFFNEGX1_27/a_66_6# 0 6.40992f **FLOATING
C2325 DFFNEGX1_27/a_23_6# 0 6.85692f **FLOATING
C2326 DFFNEGX1_27/a_34_4# 0 4.93023f **FLOATING
C2327 DFFNEGX1_27/a_2_6# 0 9.33504f **FLOATING
C2328 DFFNEGX1_16/a_66_6# 0 6.40992f **FLOATING
C2329 DFFNEGX1_16/a_23_6# 0 6.85692f **FLOATING
C2330 DFFNEGX1_16/a_34_4# 0 4.93023f **FLOATING
C2331 DFFNEGX1_16/a_2_6# 0 9.33504f **FLOATING
C2332 NOR2X1_4/A 0 22.252586f **FLOATING
C2333 out_temp_cleared[3] 0 11.608049f **FLOATING
C2334 MUX2X1_4/Y 0 9.10782f **FLOATING
C2335 MUX2X1_4/A 0 6.07278f **FLOATING
C2336 MUX2X1_4/a_2_10# 0 6.0456f **FLOATING
C2337 XOR2X1_3/a_2_6# 0 8.278139f **FLOATING
C2338 XOR2X1_3/a_13_43# 0 7.836241f **FLOATING
C2339 INVX2_66/Y 0 29.999945f **FLOATING
C2340 OAI21X1_0/a_2_6# 0 2.78652f **FLOATING
C2341 HAX1_30/a_38_6# 0 2.442f **FLOATING
C2342 FAX1_3/A 0 17.3973f **FLOATING
C2343 HAX1_30/a_41_74# 0 5.99325f **FLOATING
C2344 HAX1_30/a_2_74# 0 7.65318f **FLOATING
C2345 HAX1_41/a_38_6# 0 2.442f **FLOATING
C2346 HAX1_41/a_41_74# 0 5.99325f **FLOATING
C2347 HAX1_41/a_2_74# 0 7.65318f **FLOATING
C2348 AOI22X1_49/a_2_54# 0 6.66f **FLOATING
C2349 AOI22X1_38/a_2_54# 0 6.66f **FLOATING
C2350 AOI22X1_27/a_2_54# 0 6.66f **FLOATING
C2351 AOI22X1_16/a_2_54# 0 6.66f **FLOATING
C2352 out_global_score[17] 0 19.5105f **FLOATING
C2353 OAI21X1_27/C 0 8.08944f **FLOATING
C2354 OAI21X1_9/C 0 8.684041f **FLOATING
C2355 NOR2X1_66/A 0 30.446938f **FLOATING
C2356 OAI21X1_132/a_2_6# 0 2.78652f **FLOATING
C2357 OAI21X1_132/Y 0 9.02916f **FLOATING
C2358 OAI21X1_154/a_2_6# 0 2.78652f **FLOATING
C2359 AOI22X1_8/a_2_54# 0 6.66f **FLOATING
C2360 OAI21X1_143/a_2_6# 0 2.78652f **FLOATING
C2361 INVX2_38/Y 0 16.11543f **FLOATING
C2362 OAI21X1_121/a_2_6# 0 2.78652f **FLOATING
C2363 OAI21X1_110/a_2_6# 0 2.78652f **FLOATING
C2364 NAND2X1_99/Y 0 6.86169f **FLOATING
C2365 DFFNEGX1_127/a_66_6# 0 6.40992f **FLOATING
C2366 DFFNEGX1_127/a_23_6# 0 6.85692f **FLOATING
C2367 DFFNEGX1_127/a_34_4# 0 4.93023f **FLOATING
C2368 DFFNEGX1_127/a_2_6# 0 9.33504f **FLOATING
C2369 DFFNEGX1_138/a_66_6# 0 6.40992f **FLOATING
C2370 DFFNEGX1_138/a_23_6# 0 6.85692f **FLOATING
C2371 DFFNEGX1_138/a_34_4# 0 4.93023f **FLOATING
C2372 DFFNEGX1_138/a_2_6# 0 9.33504f **FLOATING
C2373 DFFNEGX1_116/a_66_6# 0 6.40992f **FLOATING
C2374 DFFNEGX1_116/a_23_6# 0 6.85692f **FLOATING
C2375 DFFNEGX1_116/a_34_4# 0 4.93023f **FLOATING
C2376 DFFNEGX1_116/a_2_6# 0 9.33504f **FLOATING
C2377 INVX2_194/Y 0 11.164379f **FLOATING
C2378 DFFNEGX1_105/a_66_6# 0 6.40992f **FLOATING
C2379 DFFNEGX1_105/a_23_6# 0 6.85692f **FLOATING
C2380 DFFNEGX1_105/a_34_4# 0 4.93023f **FLOATING
C2381 DFFNEGX1_105/a_2_6# 0 9.33504f **FLOATING
C2382 XOR2X1_24/a_2_6# 0 8.278139f **FLOATING
C2383 XOR2X1_24/a_13_43# 0 7.836241f **FLOATING
C2384 XOR2X1_13/Y 0 13.407301f **FLOATING
C2385 XOR2X1_13/a_2_6# 0 8.278139f **FLOATING
C2386 XOR2X1_13/a_13_43# 0 7.836241f **FLOATING
C2387 DFFNEGX1_37/a_66_6# 0 6.40992f **FLOATING
C2388 DFFNEGX1_37/a_23_6# 0 6.85692f **FLOATING
C2389 DFFNEGX1_37/a_34_4# 0 4.93023f **FLOATING
C2390 DFFNEGX1_37/a_2_6# 0 9.33504f **FLOATING
C2391 DFFNEGX1_48/a_66_6# 0 6.40992f **FLOATING
C2392 out_temp_decoded[18] 0 14.404171f **FLOATING
C2393 DFFNEGX1_48/a_23_6# 0 6.85692f **FLOATING
C2394 DFFNEGX1_48/a_34_4# 0 4.93023f **FLOATING
C2395 DFFNEGX1_48/a_2_6# 0 9.33504f **FLOATING
C2396 DFFNEGX1_59/a_66_6# 0 6.40992f **FLOATING
C2397 DFFNEGX1_59/a_23_6# 0 6.85692f **FLOATING
C2398 DFFNEGX1_59/a_34_4# 0 4.93023f **FLOATING
C2399 DFFNEGX1_59/a_2_6# 0 9.33504f **FLOATING
C2400 DFFNEGX1_26/a_66_6# 0 6.40992f **FLOATING
C2401 DFFNEGX1_26/a_23_6# 0 6.85692f **FLOATING
C2402 DFFNEGX1_26/a_34_4# 0 4.93023f **FLOATING
C2403 DFFNEGX1_26/a_2_6# 0 9.33504f **FLOATING
C2404 OAI21X1_15/Y 0 14.933821f **FLOATING
C2405 DFFNEGX1_15/a_66_6# 0 6.40992f **FLOATING
C2406 DFFNEGX1_15/a_23_6# 0 6.85692f **FLOATING
C2407 DFFNEGX1_15/a_34_4# 0 4.93023f **FLOATING
C2408 DFFNEGX1_15/a_2_6# 0 9.33504f **FLOATING
C2409 OAI22X1_75/B 0 37.43322f **FLOATING
C2410 BUFX2_10/Y 0 0.169818p **FLOATING
C2411 INVX2_186/Y 0 12.119221f **FLOATING
C2412 BUFX2_9/Y 0 0.169961p **FLOATING
C2413 INVX2_236/A 0 8.71374f **FLOATING
C2414 MUX2X1_3/Y 0 21.083282f **FLOATING
C2415 MUX2X1_3/a_2_10# 0 6.0456f **FLOATING
C2416 XOR2X1_2/a_2_6# 0 8.278139f **FLOATING
C2417 XOR2X1_2/a_13_43# 0 7.836241f **FLOATING
C2418 HAX1_40/a_38_6# 0 2.442f **FLOATING
C2419 HAX1_40/a_41_74# 0 5.99325f **FLOATING
C2420 HAX1_40/a_2_74# 0 7.65318f **FLOATING
C2421 OAI22X1_46/Y 0 12.03336f **FLOATING
C2422 AOI21X1_11/B 0 16.460398f **FLOATING
C2423 INVX2_120/Y 0 17.99601f **FLOATING
C2424 AOI22X1_59/a_2_54# 0 6.66f **FLOATING
C2425 AOI22X1_66/D 0 21.60222f **FLOATING
C2426 AOI22X1_48/a_2_54# 0 6.66f **FLOATING
C2427 AOI22X1_37/a_2_54# 0 6.66f **FLOATING
C2428 AOI22X1_26/a_2_54# 0 6.66f **FLOATING
C2429 out_global_score[7] 0 16.232399f **FLOATING
C2430 AOI22X1_15/a_2_54# 0 6.66f **FLOATING
C2431 HAX1_12/YS 0 7.00383f **FLOATING
C2432 OAI21X1_142/a_2_6# 0 2.78652f **FLOATING
C2433 OAI21X1_153/a_2_6# 0 2.78652f **FLOATING
C2434 AOI22X1_7/a_2_54# 0 6.66f **FLOATING
C2435 OAI21X1_131/a_2_6# 0 2.78652f **FLOATING
C2436 XOR2X1_29/B 0 31.720526f **FLOATING
C2437 OAI21X1_120/a_2_6# 0 2.78652f **FLOATING
C2438 INVX2_33/A 0 20.924698f **FLOATING
C2439 DFFNEGX1_137/a_66_6# 0 6.40992f **FLOATING
C2440 DFFNEGX1_137/a_23_6# 0 6.85692f **FLOATING
C2441 DFFNEGX1_137/a_34_4# 0 4.93023f **FLOATING
C2442 DFFNEGX1_137/a_2_6# 0 9.33504f **FLOATING
C2443 DFFNEGX1_126/a_66_6# 0 6.40992f **FLOATING
C2444 DFFNEGX1_126/a_23_6# 0 6.85692f **FLOATING
C2445 DFFNEGX1_126/a_34_4# 0 4.93023f **FLOATING
C2446 DFFNEGX1_126/a_2_6# 0 9.33504f **FLOATING
C2447 DFFNEGX1_115/a_66_6# 0 6.40992f **FLOATING
C2448 DFFNEGX1_115/a_23_6# 0 6.85692f **FLOATING
C2449 DFFNEGX1_115/a_34_4# 0 4.93023f **FLOATING
C2450 DFFNEGX1_115/a_2_6# 0 9.33504f **FLOATING
C2451 INVX2_195/Y 0 12.84738f **FLOATING
C2452 DFFNEGX1_104/a_66_6# 0 6.40992f **FLOATING
C2453 DFFNEGX1_104/a_23_6# 0 6.85692f **FLOATING
C2454 DFFNEGX1_104/a_34_4# 0 4.93023f **FLOATING
C2455 DFFNEGX1_104/a_2_6# 0 9.33504f **FLOATING
C2456 OAI21X1_1/A 0 42.823555f **FLOATING
C2457 XOR2X1_23/a_2_6# 0 8.278139f **FLOATING
C2458 XOR2X1_23/a_13_43# 0 7.836241f **FLOATING
C2459 XOR2X1_23/A 0 12.575009f **FLOATING
C2460 XOR2X1_12/Y 0 13.74456f **FLOATING
C2461 XOR2X1_12/a_2_6# 0 8.278139f **FLOATING
C2462 XOR2X1_12/a_13_43# 0 7.836241f **FLOATING
C2463 DFFNEGX1_69/a_66_6# 0 6.40992f **FLOATING
C2464 out_temp_cleared[22] 0 18.345211f **FLOATING
C2465 DFFNEGX1_69/a_23_6# 0 6.85692f **FLOATING
C2466 DFFNEGX1_69/a_34_4# 0 4.93023f **FLOATING
C2467 DFFNEGX1_69/a_2_6# 0 9.33504f **FLOATING
C2468 OAI22X1_6/Y 0 13.223941f **FLOATING
C2469 DFFNEGX1_36/a_66_6# 0 6.40992f **FLOATING
C2470 DFFNEGX1_36/a_23_6# 0 6.85692f **FLOATING
C2471 DFFNEGX1_36/a_34_4# 0 4.93023f **FLOATING
C2472 DFFNEGX1_36/a_2_6# 0 9.33504f **FLOATING
C2473 DFFNEGX1_47/a_66_6# 0 6.40992f **FLOATING
C2474 DFFNEGX1_47/a_23_6# 0 6.85692f **FLOATING
C2475 DFFNEGX1_47/a_34_4# 0 4.93023f **FLOATING
C2476 DFFNEGX1_47/a_2_6# 0 9.33504f **FLOATING
C2477 DFFNEGX1_58/a_66_6# 0 6.40992f **FLOATING
C2478 DFFNEGX1_58/a_23_6# 0 6.85692f **FLOATING
C2479 DFFNEGX1_58/a_34_4# 0 4.93023f **FLOATING
C2480 DFFNEGX1_58/a_2_6# 0 9.33504f **FLOATING
C2481 DFFNEGX1_14/a_66_6# 0 6.40992f **FLOATING
C2482 DFFNEGX1_14/a_23_6# 0 6.85692f **FLOATING
C2483 DFFNEGX1_14/a_34_4# 0 4.93023f **FLOATING
C2484 DFFNEGX1_14/a_2_6# 0 9.33504f **FLOATING
C2485 DFFNEGX1_25/a_66_6# 0 6.40992f **FLOATING
C2486 DFFNEGX1_25/a_23_6# 0 6.85692f **FLOATING
C2487 DFFNEGX1_25/a_34_4# 0 4.93023f **FLOATING
C2488 DFFNEGX1_25/a_2_6# 0 9.33504f **FLOATING
C2489 OAI21X1_13/Y 0 11.813461f **FLOATING
C2490 NOR2X1_79/Y 0 29.309278f **FLOATING
C2491 OR2X1_4/A 0 11.55048f **FLOATING
C2492 MUX2X1_19/A 0 6.05058f **FLOATING
C2493 OAI22X1_22/Y 0 10.309978f **FLOATING
C2494 MUX2X1_2/a_2_10# 0 6.0456f **FLOATING
C2495 XOR2X1_1/a_2_6# 0 8.278139f **FLOATING
C2496 XOR2X1_1/a_13_43# 0 7.836241f **FLOATING
C2497 OAI22X1_9/a_2_6# 0 4.25172f **FLOATING
C2498 AOI22X1_69/a_2_54# 0 6.66f **FLOATING
C2499 NOR2X1_113/Y 0 26.48169f **FLOATING
C2500 AOI22X1_58/a_2_54# 0 6.66f **FLOATING
C2501 AOI22X1_47/a_2_54# 0 6.66f **FLOATING
C2502 AOI22X1_36/a_2_54# 0 6.66f **FLOATING
C2503 AOI22X1_25/a_2_54# 0 6.66f **FLOATING
C2504 out_global_score[8] 0 16.232399f **FLOATING
C2505 AOI22X1_14/a_2_54# 0 6.66f **FLOATING
C2506 HAX1_11/YS 0 7.00383f **FLOATING
C2507 OAI21X1_54/C 0 8.08944f **FLOATING
C2508 OAI21X1_152/a_2_6# 0 2.78652f **FLOATING
C2509 AOI22X1_6/a_2_54# 0 6.66f **FLOATING
C2510 OAI21X1_141/a_2_6# 0 2.78652f **FLOATING
C2511 OAI21X1_130/a_2_6# 0 2.78652f **FLOATING
C2512 OAI21X1_130/Y 0 12.11796f **FLOATING
C2513 DFFNEGX1_136/a_66_6# 0 6.40992f **FLOATING
C2514 DFFNEGX1_136/a_23_6# 0 6.85692f **FLOATING
C2515 DFFNEGX1_136/a_34_4# 0 4.93023f **FLOATING
C2516 DFFNEGX1_136/a_2_6# 0 9.33504f **FLOATING
C2517 DFFNEGX1_125/a_66_6# 0 6.40992f **FLOATING
C2518 DFFNEGX1_125/a_23_6# 0 6.85692f **FLOATING
C2519 DFFNEGX1_125/a_34_4# 0 4.93023f **FLOATING
C2520 DFFNEGX1_125/a_2_6# 0 9.33504f **FLOATING
C2521 INVX2_185/Y 0 13.04382f **FLOATING
C2522 DFFNEGX1_114/a_66_6# 0 6.40992f **FLOATING
C2523 DFFNEGX1_114/a_23_6# 0 6.85692f **FLOATING
C2524 DFFNEGX1_114/a_34_4# 0 4.93023f **FLOATING
C2525 DFFNEGX1_114/a_2_6# 0 9.33504f **FLOATING
C2526 DFFNEGX1_103/a_66_6# 0 6.40992f **FLOATING
C2527 DFFNEGX1_103/a_23_6# 0 6.85692f **FLOATING
C2528 DFFNEGX1_103/a_34_4# 0 4.93023f **FLOATING
C2529 DFFNEGX1_103/a_2_6# 0 9.33504f **FLOATING
C2530 INVX2_207/Y 0 13.04382f **FLOATING
C2531 NOR2X1_65/A 0 25.310246f **FLOATING
C2532 XOR2X1_22/a_2_6# 0 8.278139f **FLOATING
C2533 XOR2X1_22/a_13_43# 0 7.836241f **FLOATING
C2534 XOR2X1_11/a_2_6# 0 8.278139f **FLOATING
C2535 XOR2X1_11/a_13_43# 0 7.836241f **FLOATING
C2536 DFFNEGX1_79/a_66_6# 0 6.40992f **FLOATING
C2537 DFFNEGX1_79/a_23_6# 0 6.85692f **FLOATING
C2538 DFFNEGX1_79/a_34_4# 0 4.93023f **FLOATING
C2539 DFFNEGX1_79/a_2_6# 0 9.33504f **FLOATING
C2540 DFFNEGX1_46/a_66_6# 0 6.40992f **FLOATING
C2541 DFFNEGX1_46/a_23_6# 0 6.85692f **FLOATING
C2542 DFFNEGX1_46/a_34_4# 0 4.93023f **FLOATING
C2543 DFFNEGX1_46/a_2_6# 0 9.33504f **FLOATING
C2544 DFFNEGX1_57/a_66_6# 0 6.40992f **FLOATING
C2545 DFFNEGX1_57/a_23_6# 0 6.85692f **FLOATING
C2546 DFFNEGX1_57/a_34_4# 0 4.93023f **FLOATING
C2547 DFFNEGX1_57/a_2_6# 0 9.33504f **FLOATING
C2548 DFFNEGX1_68/a_66_6# 0 6.40992f **FLOATING
C2549 out_temp_cleared[23] 0 24.599731f **FLOATING
C2550 DFFNEGX1_68/a_23_6# 0 6.85692f **FLOATING
C2551 DFFNEGX1_68/a_34_4# 0 4.93023f **FLOATING
C2552 DFFNEGX1_68/a_2_6# 0 9.33504f **FLOATING
C2553 DFFNEGX1_35/a_66_6# 0 6.40992f **FLOATING
C2554 DFFNEGX1_35/a_23_6# 0 6.85692f **FLOATING
C2555 DFFNEGX1_35/a_34_4# 0 4.93023f **FLOATING
C2556 DFFNEGX1_35/a_2_6# 0 9.33504f **FLOATING
C2557 DFFNEGX1_24/a_66_6# 0 6.40992f **FLOATING
C2558 DFFNEGX1_24/a_23_6# 0 6.85692f **FLOATING
C2559 DFFNEGX1_24/a_34_4# 0 4.93023f **FLOATING
C2560 DFFNEGX1_24/a_2_6# 0 9.33504f **FLOATING
C2561 DFFNEGX1_13/a_66_6# 0 6.40992f **FLOATING
C2562 DFFNEGX1_13/a_23_6# 0 6.85692f **FLOATING
C2563 DFFNEGX1_13/a_34_4# 0 4.93023f **FLOATING
C2564 DFFNEGX1_13/a_2_6# 0 9.33504f **FLOATING
C2565 NOR2X1_5/A 0 19.771889f **FLOATING
C2566 OR2X1_2/A 0 9.031079f **FLOATING
C2567 OAI21X1_102/Y 0 10.471021f **FLOATING
C2568 MUX2X1_1/Y 0 7.2063f **FLOATING
C2569 MUX2X1_1/a_2_10# 0 6.0456f **FLOATING
C2570 XOR2X1_0/Y 0 10.83774f **FLOATING
C2571 XOR2X1_0/a_2_6# 0 8.278139f **FLOATING
C2572 XOR2X1_0/a_13_43# 0 7.836241f **FLOATING
C2573 OAI22X1_8/a_2_6# 0 4.25172f **FLOATING
C2574 AOI21X1_12/A 0 11.354759f **FLOATING
C2575 OAI22X1_51/Y 0 8.5758f **FLOATING
C2576 AOI22X1_68/a_2_54# 0 6.66f **FLOATING
C2577 AOI22X1_57/a_2_54# 0 6.66f **FLOATING
C2578 AOI22X1_57/A 0 6.59574f **FLOATING
C2579 AOI22X1_35/a_2_54# 0 6.66f **FLOATING
C2580 AOI22X1_46/a_2_54# 0 6.66f **FLOATING
C2581 AOI22X1_13/a_2_54# 0 6.66f **FLOATING
C2582 AOI22X1_24/a_2_54# 0 6.66f **FLOATING
C2583 OAI21X1_62/C 0 6.87006f **FLOATING
C2584 OAI21X1_21/C 0 8.08944f **FLOATING
C2585 OAI21X1_3/A 0 18.061888f **FLOATING
C2586 OAI21X1_162/a_2_6# 0 2.78652f **FLOATING
C2587 OAI21X1_151/a_2_6# 0 2.78652f **FLOATING
C2588 OAI21X1_140/a_2_6# 0 2.78652f **FLOATING
C2589 AOI22X1_5/a_2_54# 0 6.66f **FLOATING
C2590 out_global_score[28] 0 18.439949f **FLOATING
C2591 DFFNEGX1_124/a_66_6# 0 6.40992f **FLOATING
C2592 DFFNEGX1_124/a_23_6# 0 6.85692f **FLOATING
C2593 DFFNEGX1_124/a_34_4# 0 4.93023f **FLOATING
C2594 DFFNEGX1_124/a_2_6# 0 9.33504f **FLOATING
C2595 DFFNEGX1_135/a_66_6# 0 6.40992f **FLOATING
C2596 DFFNEGX1_135/a_23_6# 0 6.85692f **FLOATING
C2597 DFFNEGX1_135/a_34_4# 0 4.93023f **FLOATING
C2598 DFFNEGX1_135/a_2_6# 0 9.33504f **FLOATING
C2599 DFFNEGX1_113/a_66_6# 0 6.40992f **FLOATING
C2600 DFFNEGX1_113/a_23_6# 0 6.85692f **FLOATING
C2601 DFFNEGX1_113/a_34_4# 0 4.93023f **FLOATING
C2602 DFFNEGX1_113/a_2_6# 0 9.33504f **FLOATING
C2603 DFFNEGX1_102/a_66_6# 0 6.40992f **FLOATING
C2604 DFFNEGX1_102/a_23_6# 0 6.85692f **FLOATING
C2605 DFFNEGX1_102/a_34_4# 0 4.93023f **FLOATING
C2606 DFFNEGX1_102/a_2_6# 0 9.33504f **FLOATING
C2607 INVX2_208/Y 0 10.975981f **FLOATING
C2608 gnd 0 4.69506p **FLOATING
C2609 XOR2X1_21/a_2_6# 0 8.278139f **FLOATING
C2610 XOR2X1_21/a_13_43# 0 7.836241f **FLOATING
C2611 NOR2X1_0/B 0 21.81033f **FLOATING
C2612 XOR2X1_10/a_2_6# 0 8.278139f **FLOATING
C2613 XOR2X1_10/a_13_43# 0 7.836241f **FLOATING
C2614 DFFNEGX1_89/a_66_6# 0 6.40992f **FLOATING
C2615 DFFNEGX1_89/a_23_6# 0 6.85692f **FLOATING
C2616 DFFNEGX1_89/a_34_4# 0 4.93023f **FLOATING
C2617 DFFNEGX1_89/a_2_6# 0 9.33504f **FLOATING
C2618 DFFNEGX1_78/a_66_6# 0 6.40992f **FLOATING
C2619 DFFNEGX1_78/a_23_6# 0 6.85692f **FLOATING
C2620 DFFNEGX1_78/a_34_4# 0 4.93023f **FLOATING
C2621 DFFNEGX1_78/a_2_6# 0 9.33504f **FLOATING
C2622 OAI22X1_15/Y 0 11.28756f **FLOATING
C2623 DFFNEGX1_67/a_66_6# 0 6.40992f **FLOATING
C2624 DFFNEGX1_67/a_23_6# 0 6.85692f **FLOATING
C2625 DFFNEGX1_67/a_34_4# 0 4.93023f **FLOATING
C2626 DFFNEGX1_67/a_2_6# 0 9.33504f **FLOATING
C2627 OAI22X1_4/Y 0 10.71954f **FLOATING
C2628 DFFNEGX1_45/a_66_6# 0 6.40992f **FLOATING
C2629 DFFNEGX1_45/a_23_6# 0 6.85692f **FLOATING
C2630 DFFNEGX1_45/a_34_4# 0 4.93023f **FLOATING
C2631 DFFNEGX1_45/a_2_6# 0 9.33504f **FLOATING
C2632 DFFNEGX1_56/a_66_6# 0 6.40992f **FLOATING
C2633 out_temp_decoded[10] 0 18.316711f **FLOATING
C2634 DFFNEGX1_56/a_23_6# 0 6.85692f **FLOATING
C2635 DFFNEGX1_56/a_34_4# 0 4.93023f **FLOATING
C2636 DFFNEGX1_56/a_2_6# 0 9.33504f **FLOATING
C2637 DFFNEGX1_34/a_66_6# 0 6.40992f **FLOATING
C2638 DFFNEGX1_34/a_23_6# 0 6.85692f **FLOATING
C2639 DFFNEGX1_34/a_34_4# 0 4.93023f **FLOATING
C2640 DFFNEGX1_34/a_2_6# 0 9.33504f **FLOATING
C2641 AND2X2_10/Y 0 12.385349f **FLOATING
C2642 DFFNEGX1_12/a_66_6# 0 6.40992f **FLOATING
C2643 DFFNEGX1_12/a_23_6# 0 6.85692f **FLOATING
C2644 DFFNEGX1_12/a_34_4# 0 4.93023f **FLOATING
C2645 DFFNEGX1_12/a_2_6# 0 9.33504f **FLOATING
C2646 DFFNEGX1_23/a_66_6# 0 6.40992f **FLOATING
C2647 DFFNEGX1_23/a_23_6# 0 6.85692f **FLOATING
C2648 DFFNEGX1_23/a_34_4# 0 4.93023f **FLOATING
C2649 DFFNEGX1_23/a_2_6# 0 9.33504f **FLOATING
C2650 HAX1_42/A 0 22.18134f **FLOATING
C2651 MUX2X1_25/Y 0 6.36198f **FLOATING
C2652 NAND3X1_39/A 0 7.812f **FLOATING
C2653 OAI21X1_91/Y 0 10.0662f **FLOATING
C2654 INVX2_221/A 0 9.369361f **FLOATING
C2655 MUX2X1_0/Y 0 6.36198f **FLOATING
C2656 MUX2X1_0/a_2_10# 0 6.0456f **FLOATING
C2657 INVX2_49/Y 0 7.36035f **FLOATING
C2658 out_mines[9] 0 80.68047f **FLOATING
C2659 OAI22X1_7/a_2_6# 0 4.25172f **FLOATING
C2660 AOI22X1_67/a_2_54# 0 6.66f **FLOATING
C2661 AOI22X1_78/a_2_54# 0 6.66f **FLOATING
C2662 NOR2X1_121/Y 0 22.712698f **FLOATING
C2663 AOI22X1_56/a_2_54# 0 6.66f **FLOATING
C2664 INVX2_47/A 0 13.21332f **FLOATING
C2665 AOI22X1_34/a_2_54# 0 6.66f **FLOATING
C2666 AOI22X1_45/a_2_54# 0 6.66f **FLOATING
C2667 AOI22X1_12/a_2_54# 0 6.66f **FLOATING
C2668 HAX1_9/YS 0 7.00383f **FLOATING
C2669 AOI22X1_23/a_2_54# 0 6.66f **FLOATING
C2670 OAI21X1_82/C 0 11.319602f **FLOATING
C2671 OAI21X1_60/A 0 7.9392f **FLOATING
C2672 NAND2X1_14/Y 0 13.240861f **FLOATING
C2673 OAI21X1_19/C 0 8.507041f **FLOATING
C2674 OAI21X1_161/a_2_6# 0 2.78652f **FLOATING
C2675 OAI21X1_150/a_2_6# 0 2.78652f **FLOATING
C2676 AOI22X1_4/a_2_54# 0 6.66f **FLOATING
C2677 INVX2_258/Y 0 0.130294p **FLOATING
C2678 HAX1_1/YS 0 7.00383f **FLOATING
C2679 DFFNEGX1_123/a_66_6# 0 6.40992f **FLOATING
C2680 DFFNEGX1_123/a_23_6# 0 6.85692f **FLOATING
C2681 DFFNEGX1_123/a_34_4# 0 4.93023f **FLOATING
C2682 DFFNEGX1_123/a_2_6# 0 9.33504f **FLOATING
C2683 DFFNEGX1_134/a_66_6# 0 6.40992f **FLOATING
C2684 DFFNEGX1_134/a_23_6# 0 6.85692f **FLOATING
C2685 DFFNEGX1_134/a_34_4# 0 4.93023f **FLOATING
C2686 DFFNEGX1_134/a_2_6# 0 9.33504f **FLOATING
C2687 DFFNEGX1_112/a_66_6# 0 6.40992f **FLOATING
C2688 DFFNEGX1_112/a_23_6# 0 6.85692f **FLOATING
C2689 DFFNEGX1_112/a_34_4# 0 4.93023f **FLOATING
C2690 DFFNEGX1_112/a_2_6# 0 9.33504f **FLOATING
C2691 INVX2_198/Y 0 12.20658f **FLOATING
C2692 DFFNEGX1_101/a_66_6# 0 6.40992f **FLOATING
C2693 DFFNEGX1_101/a_23_6# 0 6.85692f **FLOATING
C2694 DFFNEGX1_101/a_34_4# 0 4.93023f **FLOATING
C2695 DFFNEGX1_101/a_2_6# 0 9.33504f **FLOATING
C2696 INVX2_209/Y 0 10.173361f **FLOATING
C2697 XOR2X1_20/a_2_6# 0 8.278139f **FLOATING
C2698 XOR2X1_20/a_13_43# 0 7.836241f **FLOATING
C2699 AND2X2_9/a_2_6# 0 6.03567f **FLOATING
C2700 DFFNEGX1_88/a_66_6# 0 6.40992f **FLOATING
C2701 DFFNEGX1_88/a_23_6# 0 6.85692f **FLOATING
C2702 DFFNEGX1_88/a_34_4# 0 4.93023f **FLOATING
C2703 DFFNEGX1_88/a_2_6# 0 9.33504f **FLOATING
C2704 DFFNEGX1_99/a_66_6# 0 6.40992f **FLOATING
C2705 DFFNEGX1_99/a_23_6# 0 6.85692f **FLOATING
C2706 DFFNEGX1_99/a_34_4# 0 4.93023f **FLOATING
C2707 DFFNEGX1_99/a_2_6# 0 9.33504f **FLOATING
C2708 INVX2_211/Y 0 10.975981f **FLOATING
C2709 DFFNEGX1_66/a_66_6# 0 6.40992f **FLOATING
C2710 out_temp_decoded[0] 0 8.23572f **FLOATING
C2711 DFFNEGX1_66/a_23_6# 0 6.85692f **FLOATING
C2712 DFFNEGX1_66/a_34_4# 0 4.93023f **FLOATING
C2713 DFFNEGX1_66/a_2_6# 0 9.33504f **FLOATING
C2714 DFFNEGX1_77/a_66_6# 0 6.40992f **FLOATING
C2715 DFFNEGX1_77/a_23_6# 0 6.85692f **FLOATING
C2716 DFFNEGX1_77/a_34_4# 0 4.93023f **FLOATING
C2717 DFFNEGX1_77/a_2_6# 0 9.33504f **FLOATING
C2718 DFFNEGX1_55/a_66_6# 0 6.40992f **FLOATING
C2719 out_temp_decoded[11] 0 17.65266f **FLOATING
C2720 DFFNEGX1_55/a_23_6# 0 6.85692f **FLOATING
C2721 DFFNEGX1_55/a_34_4# 0 4.93023f **FLOATING
C2722 DFFNEGX1_55/a_2_6# 0 9.33504f **FLOATING
C2723 DFFNEGX1_44/a_66_6# 0 6.40992f **FLOATING
C2724 DFFNEGX1_44/a_23_6# 0 6.85692f **FLOATING
C2725 DFFNEGX1_44/a_34_4# 0 4.93023f **FLOATING
C2726 DFFNEGX1_44/a_2_6# 0 9.33504f **FLOATING
C2727 DFFNEGX1_11/a_66_6# 0 6.40992f **FLOATING
C2728 DFFNEGX1_11/a_23_6# 0 6.85692f **FLOATING
C2729 DFFNEGX1_11/a_34_4# 0 4.93023f **FLOATING
C2730 DFFNEGX1_11/a_2_6# 0 9.33504f **FLOATING
C2731 DFFNEGX1_22/a_66_6# 0 6.40992f **FLOATING
C2732 DFFNEGX1_22/a_23_6# 0 6.85692f **FLOATING
C2733 DFFNEGX1_22/a_34_4# 0 4.93023f **FLOATING
C2734 DFFNEGX1_22/a_2_6# 0 9.33504f **FLOATING
C2735 DFFNEGX1_33/a_66_6# 0 6.40992f **FLOATING
C2736 DFFNEGX1_33/a_23_6# 0 6.85692f **FLOATING
C2737 DFFNEGX1_33/a_34_4# 0 4.93023f **FLOATING
C2738 DFFNEGX1_33/a_2_6# 0 9.33504f **FLOATING
C2739 INVX2_72/Y 0 30.400656f **FLOATING
C2740 XNOR2X1_9/Y 0 9.938669f **FLOATING
C2741 XNOR2X1_9/a_2_6# 0 6.77121f **FLOATING
C2742 XNOR2X1_9/a_12_41# 0 7.905991f **FLOATING
C2743 INVX2_241/Y 0 12.69708f **FLOATING
C2744 NAND3X1_7/C 0 9.33078f **FLOATING
C2745 OAI21X1_72/B 0 9.99078f **FLOATING
C2746 OAI22X1_26/Y 0 9.78018f **FLOATING
C2747 OAI21X1_90/Y 0 11.521741f **FLOATING
C2748 INVX2_48/Y 0 22.640278f **FLOATING
C2749 out_mines[8] 0 0.119332p **FLOATING
C2750 OAI22X1_6/a_2_6# 0 4.25172f **FLOATING
C2751 OAI22X1_52/B 0 36.735878f **FLOATING
C2752 AOI22X1_77/a_2_54# 0 6.66f **FLOATING
C2753 AOI22X1_66/a_2_54# 0 6.66f **FLOATING
C2754 NOR2X1_111/Y 0 20.573608f **FLOATING
C2755 AOI22X1_55/a_2_54# 0 6.66f **FLOATING
C2756 INVX2_41/Y 0 5.8155f **FLOATING
C2757 AOI22X1_44/a_2_54# 0 6.66f **FLOATING
C2758 AOI22X1_11/a_2_54# 0 6.66f **FLOATING
C2759 AOI22X1_33/a_2_54# 0 6.66f **FLOATING
C2760 AOI22X1_22/a_2_54# 0 6.66f **FLOATING
C2761 out_global_score[11] 0 21.624811f **FLOATING
C2762 OAI21X1_35/C 0 6.87006f **FLOATING
C2763 OAI21X1_160/a_2_6# 0 2.78652f **FLOATING
C2764 AOI22X1_3/a_2_54# 0 6.66f **FLOATING
C2765 DFFNEGX1_122/a_66_6# 0 6.40992f **FLOATING
C2766 DFFNEGX1_122/a_23_6# 0 6.85692f **FLOATING
C2767 DFFNEGX1_122/a_34_4# 0 4.93023f **FLOATING
C2768 DFFNEGX1_122/a_2_6# 0 9.33504f **FLOATING
C2769 DFFNEGX1_133/a_66_6# 0 6.40992f **FLOATING
C2770 DFFNEGX1_133/a_23_6# 0 6.85692f **FLOATING
C2771 DFFNEGX1_133/a_34_4# 0 4.93023f **FLOATING
C2772 DFFNEGX1_133/a_2_6# 0 9.33504f **FLOATING
C2773 NOR2X1_118/Y 0 12.576301f **FLOATING
C2774 DFFNEGX1_100/a_66_6# 0 6.40992f **FLOATING
C2775 DFFNEGX1_100/a_23_6# 0 6.85692f **FLOATING
C2776 DFFNEGX1_100/a_34_4# 0 4.93023f **FLOATING
C2777 DFFNEGX1_100/a_2_6# 0 9.33504f **FLOATING
C2778 INVX2_210/Y 0 13.888141f **FLOATING
C2779 DFFNEGX1_111/a_66_6# 0 6.40992f **FLOATING
C2780 DFFNEGX1_111/a_23_6# 0 6.85692f **FLOATING
C2781 DFFNEGX1_111/a_34_4# 0 4.93023f **FLOATING
C2782 DFFNEGX1_111/a_2_6# 0 9.33504f **FLOATING
C2783 AND2X2_8/a_2_6# 0 6.03567f **FLOATING
C2784 DFFNEGX1_87/a_66_6# 0 6.40992f **FLOATING
C2785 out_temp_cleared[4] 0 8.23572f **FLOATING
C2786 DFFNEGX1_87/a_23_6# 0 6.85692f **FLOATING
C2787 DFFNEGX1_87/a_34_4# 0 4.93023f **FLOATING
C2788 DFFNEGX1_87/a_2_6# 0 9.33504f **FLOATING
C2789 DFFNEGX1_98/a_66_6# 0 6.40992f **FLOATING
C2790 DFFNEGX1_98/a_23_6# 0 6.85692f **FLOATING
C2791 DFFNEGX1_98/a_34_4# 0 4.93023f **FLOATING
C2792 DFFNEGX1_98/a_2_6# 0 9.33504f **FLOATING
C2793 INVX2_212/Y 0 13.465981f **FLOATING
C2794 DFFNEGX1_65/a_66_6# 0 6.40992f **FLOATING
C2795 DFFNEGX1_65/a_23_6# 0 6.85692f **FLOATING
C2796 DFFNEGX1_65/a_34_4# 0 4.93023f **FLOATING
C2797 DFFNEGX1_65/a_2_6# 0 9.33504f **FLOATING
C2798 DFFNEGX1_76/a_66_6# 0 6.40992f **FLOATING
C2799 out_temp_cleared[15] 0 8.23572f **FLOATING
C2800 DFFNEGX1_76/a_23_6# 0 6.85692f **FLOATING
C2801 DFFNEGX1_76/a_34_4# 0 4.93023f **FLOATING
C2802 DFFNEGX1_76/a_2_6# 0 9.33504f **FLOATING
C2803 DFFNEGX1_54/a_66_6# 0 6.40992f **FLOATING
C2804 DFFNEGX1_54/a_23_6# 0 6.85692f **FLOATING
C2805 DFFNEGX1_54/a_34_4# 0 4.93023f **FLOATING
C2806 DFFNEGX1_54/a_2_6# 0 9.33504f **FLOATING
C2807 OAI21X1_94/Y 0 11.833501f **FLOATING
C2808 DFFNEGX1_43/a_66_6# 0 6.40992f **FLOATING
C2809 DFFNEGX1_43/a_23_6# 0 6.85692f **FLOATING
C2810 DFFNEGX1_43/a_34_4# 0 4.93023f **FLOATING
C2811 DFFNEGX1_43/a_2_6# 0 9.33504f **FLOATING
C2812 OAI21X1_105/Y 0 12.550261f **FLOATING
C2813 DFFNEGX1_21/a_66_6# 0 6.40992f **FLOATING
C2814 DFFNEGX1_21/a_23_6# 0 6.85692f **FLOATING
C2815 DFFNEGX1_21/a_34_4# 0 4.93023f **FLOATING
C2816 DFFNEGX1_21/a_2_6# 0 9.33504f **FLOATING
C2817 DFFNEGX1_10/a_66_6# 0 6.40992f **FLOATING
C2818 DFFNEGX1_10/a_23_6# 0 6.85692f **FLOATING
C2819 DFFNEGX1_10/a_34_4# 0 4.93023f **FLOATING
C2820 DFFNEGX1_10/a_2_6# 0 9.33504f **FLOATING
C2821 DFFNEGX1_32/a_66_6# 0 6.40992f **FLOATING
C2822 DFFNEGX1_32/a_23_6# 0 6.85692f **FLOATING
C2823 DFFNEGX1_32/a_34_4# 0 4.93023f **FLOATING
C2824 DFFNEGX1_32/a_2_6# 0 9.33504f **FLOATING
C2825 INVX2_75/Y 0 22.01316f **FLOATING
C2826 XNOR2X1_8/Y 0 12.390629f **FLOATING
C2827 XNOR2X1_8/a_2_6# 0 6.77121f **FLOATING
C2828 XNOR2X1_8/a_12_41# 0 7.905991f **FLOATING
C2829 INVX2_192/Y 0 10.626481f **FLOATING
C2830 INVX2_40/A 0 58.128586f **FLOATING
C2831 OAI22X1_5/a_2_6# 0 4.25172f **FLOATING
C2832 AOI22X1_76/a_2_54# 0 6.66f **FLOATING
C2833 AOI22X1_65/a_2_54# 0 6.66f **FLOATING
C2834 AOI22X1_54/a_2_54# 0 6.66f **FLOATING
C2835 AOI22X1_43/a_2_54# 0 6.66f **FLOATING
C2836 AOI22X1_10/a_2_54# 0 6.66f **FLOATING
C2837 AOI22X1_32/a_2_54# 0 6.66f **FLOATING
C2838 AOI22X1_21/a_2_54# 0 6.66f **FLOATING
C2839 NOR2X1_47/Y 0 6.2739f **FLOATING
C2840 OAI21X1_59/B 0 8.598122f **FLOATING
C2841 OAI21X1_79/B 0 7.384621f **FLOATING
C2842 OAI21X1_33/C 0 6.87006f **FLOATING
C2843 AOI22X1_2/a_2_54# 0 6.66f **FLOATING
C2844 MUX2X1_19/a_2_10# 0 6.0456f **FLOATING
C2845 DFFNEGX1_132/a_66_6# 0 6.40992f **FLOATING
C2846 DFFNEGX1_132/a_23_6# 0 6.85692f **FLOATING
C2847 DFFNEGX1_132/a_34_4# 0 4.93023f **FLOATING
C2848 DFFNEGX1_132/a_2_6# 0 9.33504f **FLOATING
C2849 DFFNEGX1_121/a_66_6# 0 6.40992f **FLOATING
C2850 DFFNEGX1_121/a_23_6# 0 6.85692f **FLOATING
C2851 DFFNEGX1_121/a_34_4# 0 4.93023f **FLOATING
C2852 DFFNEGX1_121/a_2_6# 0 9.33504f **FLOATING
C2853 INVX2_189/Y 0 12.078781f **FLOATING
C2854 DFFNEGX1_110/a_66_6# 0 6.40992f **FLOATING
C2855 DFFNEGX1_110/a_23_6# 0 6.85692f **FLOATING
C2856 DFFNEGX1_110/a_34_4# 0 4.93023f **FLOATING
C2857 DFFNEGX1_110/a_2_6# 0 9.33504f **FLOATING
C2858 INVX2_25/Y 0 10.67082f **FLOATING
C2859 AND2X2_7/a_2_6# 0 6.03567f **FLOATING
C2860 DFFNEGX1_97/a_66_6# 0 6.40992f **FLOATING
C2861 DFFNEGX1_97/a_23_6# 0 6.85692f **FLOATING
C2862 DFFNEGX1_97/a_34_4# 0 4.93023f **FLOATING
C2863 DFFNEGX1_97/a_2_6# 0 9.33504f **FLOATING
C2864 DFFNEGX1_86/a_66_6# 0 6.40992f **FLOATING
C2865 DFFNEGX1_86/a_23_6# 0 6.85692f **FLOATING
C2866 DFFNEGX1_86/a_34_4# 0 4.93023f **FLOATING
C2867 DFFNEGX1_86/a_2_6# 0 9.33504f **FLOATING
C2868 OAI22X1_23/Y 0 14.187271f **FLOATING
C2869 DFFNEGX1_64/a_66_6# 0 6.40992f **FLOATING
C2870 DFFNEGX1_64/a_23_6# 0 6.85692f **FLOATING
C2871 DFFNEGX1_64/a_34_4# 0 4.93023f **FLOATING
C2872 DFFNEGX1_64/a_2_6# 0 9.33504f **FLOATING
C2873 DFFNEGX1_75/a_66_6# 0 6.40992f **FLOATING
C2874 out_temp_cleared[16] 0 19.11243f **FLOATING
C2875 DFFNEGX1_75/a_23_6# 0 6.85692f **FLOATING
C2876 DFFNEGX1_75/a_34_4# 0 4.93023f **FLOATING
C2877 DFFNEGX1_75/a_2_6# 0 9.33504f **FLOATING
C2878 OAI22X1_12/Y 0 13.30176f **FLOATING
C2879 DFFNEGX1_53/a_66_6# 0 6.40992f **FLOATING
C2880 DFFNEGX1_53/a_23_6# 0 6.85692f **FLOATING
C2881 DFFNEGX1_53/a_34_4# 0 4.93023f **FLOATING
C2882 DFFNEGX1_53/a_2_6# 0 9.33504f **FLOATING
C2883 DFFNEGX1_42/a_66_6# 0 6.40992f **FLOATING
C2884 DFFNEGX1_42/a_23_6# 0 6.85692f **FLOATING
C2885 DFFNEGX1_42/a_34_4# 0 4.93023f **FLOATING
C2886 DFFNEGX1_42/a_2_6# 0 9.33504f **FLOATING
C2887 DFFNEGX1_20/a_66_6# 0 6.40992f **FLOATING
C2888 DFFNEGX1_20/a_23_6# 0 6.85692f **FLOATING
C2889 DFFNEGX1_20/a_34_4# 0 4.93023f **FLOATING
C2890 DFFNEGX1_20/a_2_6# 0 9.33504f **FLOATING
C2891 DFFNEGX1_31/a_66_6# 0 6.40992f **FLOATING
C2892 DFFNEGX1_31/a_23_6# 0 6.85692f **FLOATING
C2893 DFFNEGX1_31/a_34_4# 0 4.93023f **FLOATING
C2894 DFFNEGX1_31/a_2_6# 0 9.33504f **FLOATING
C2895 XNOR2X1_7/Y 0 10.897471f **FLOATING
C2896 XNOR2X1_7/a_2_6# 0 6.77121f **FLOATING
C2897 XNOR2X1_7/a_12_41# 0 7.905991f **FLOATING
C2898 BUFX2_5/Y 0 0.169899p **FLOATING
C2899 INVX2_46/Y 0 9.781441f **FLOATING
C2900 out_temp_decoded[22] 0 23.30919f **FLOATING
C2901 INVX2_35/Y 0 14.799479f **FLOATING
C2902 OAI22X1_4/a_2_6# 0 4.25172f **FLOATING
C2903 OAI22X1_44/Y 0 9.545579f **FLOATING
C2904 OAI22X1_41/Y 0 10.683782f **FLOATING
C2905 AOI22X1_64/a_2_54# 0 6.66f **FLOATING
C2906 AOI22X1_53/a_2_54# 0 6.66f **FLOATING
C2907 XOR2X1_27/Y 0 17.427149f **FLOATING
C2908 AOI22X1_75/a_2_54# 0 6.66f **FLOATING
C2909 AOI22X1_42/a_2_54# 0 6.66f **FLOATING
C2910 AOI22X1_31/a_2_54# 0 6.66f **FLOATING
C2911 AOI22X1_20/a_2_54# 0 6.66f **FLOATING
C2912 HAX1_17/YS 0 7.00383f **FLOATING
C2913 NOR2X1_63/B 0 45.838127f **FLOATING
C2914 AOI22X1_1/a_2_54# 0 6.66f **FLOATING
C2915 MUX2X1_29/Y 0 8.313899f **FLOATING
C2916 MUX2X1_29/A 0 6.05058f **FLOATING
C2917 MUX2X1_29/a_2_10# 0 6.0456f **FLOATING
C2918 DFFNEGX1_131/a_66_6# 0 6.40992f **FLOATING
C2919 DFFNEGX1_131/a_23_6# 0 6.85692f **FLOATING
C2920 DFFNEGX1_131/a_34_4# 0 4.93023f **FLOATING
C2921 DFFNEGX1_131/a_2_6# 0 9.33504f **FLOATING
C2922 DFFNEGX1_142/a_66_6# 0 6.40992f **FLOATING
C2923 DFFNEGX1_142/a_23_6# 0 6.85692f **FLOATING
C2924 DFFNEGX1_142/a_34_4# 0 4.93023f **FLOATING
C2925 DFFNEGX1_142/a_2_6# 0 9.33504f **FLOATING
C2926 MUX2X1_18/a_2_10# 0 6.0456f **FLOATING
C2927 DFFNEGX1_120/a_66_6# 0 6.40992f **FLOATING
C2928 DFFNEGX1_120/a_23_6# 0 6.85692f **FLOATING
C2929 DFFNEGX1_120/a_34_4# 0 4.93023f **FLOATING
C2930 DFFNEGX1_120/a_2_6# 0 9.33504f **FLOATING
C2931 AND2X2_6/a_2_6# 0 6.03567f **FLOATING
C2932 DFFNEGX1_96/a_66_6# 0 6.40992f **FLOATING
C2933 DFFNEGX1_96/a_23_6# 0 6.85692f **FLOATING
C2934 DFFNEGX1_96/a_34_4# 0 4.93023f **FLOATING
C2935 DFFNEGX1_96/a_2_6# 0 9.33504f **FLOATING
C2936 DFFNEGX1_63/a_66_6# 0 6.40992f **FLOATING
C2937 DFFNEGX1_63/a_23_6# 0 6.85692f **FLOATING
C2938 DFFNEGX1_63/a_34_4# 0 4.93023f **FLOATING
C2939 DFFNEGX1_63/a_2_6# 0 9.33504f **FLOATING
C2940 DFFNEGX1_85/a_66_6# 0 6.40992f **FLOATING
C2941 DFFNEGX1_85/a_23_6# 0 6.85692f **FLOATING
C2942 DFFNEGX1_85/a_34_4# 0 4.93023f **FLOATING
C2943 DFFNEGX1_85/a_2_6# 0 9.33504f **FLOATING
C2944 DFFNEGX1_74/a_66_6# 0 6.40992f **FLOATING
C2945 DFFNEGX1_74/a_23_6# 0 6.85692f **FLOATING
C2946 DFFNEGX1_74/a_34_4# 0 4.93023f **FLOATING
C2947 DFFNEGX1_74/a_2_6# 0 9.33504f **FLOATING
C2948 OAI22X1_11/Y 0 12.16164f **FLOATING
C2949 DFFNEGX1_41/a_66_6# 0 6.40992f **FLOATING
C2950 DFFNEGX1_41/a_23_6# 0 6.85692f **FLOATING
C2951 DFFNEGX1_41/a_34_4# 0 4.93023f **FLOATING
C2952 DFFNEGX1_41/a_2_6# 0 9.33504f **FLOATING
C2953 OAI21X1_107/Y 0 12.616739f **FLOATING
C2954 DFFNEGX1_52/a_66_6# 0 6.40992f **FLOATING
C2955 DFFNEGX1_52/a_23_6# 0 6.85692f **FLOATING
C2956 DFFNEGX1_52/a_34_4# 0 4.93023f **FLOATING
C2957 DFFNEGX1_52/a_2_6# 0 9.33504f **FLOATING
C2958 OAI21X1_96/Y 0 11.105461f **FLOATING
C2959 DFFNEGX1_30/a_66_6# 0 6.40992f **FLOATING
C2960 DFFNEGX1_30/a_23_6# 0 6.85692f **FLOATING
C2961 DFFNEGX1_30/a_34_4# 0 4.93023f **FLOATING
C2962 DFFNEGX1_30/a_2_6# 0 9.33504f **FLOATING
C2963 INVX2_74/Y 0 34.153152f **FLOATING
C2964 INVX2_69/Y 0 14.88096f **FLOATING
C2965 XNOR2X1_6/a_2_6# 0 6.77121f **FLOATING
C2966 XNOR2X1_6/a_12_41# 0 7.905991f **FLOATING
C2967 NOR2X1_91/A 0 12.053729f **FLOATING
C2968 OAI21X1_51/C 0 8.146441f **FLOATING
C2969 OAI21X1_25/C 0 10.930439f **FLOATING
C2970 OAI21X1_19/a_2_6# 0 2.78652f **FLOATING
C2971 out_temp_decoded[23] 0 30.223349f **FLOATING
C2972 OAI22X1_3/a_2_6# 0 4.25172f **FLOATING
C2973 AOI21X1_14/Y 0 13.423109f **FLOATING
C2974 AOI22X1_63/a_2_54# 0 6.66f **FLOATING
C2975 AOI22X1_52/a_2_54# 0 6.66f **FLOATING
C2976 XOR2X1_17/Y 0 15.560282f **FLOATING
C2977 AOI22X1_74/a_2_54# 0 6.66f **FLOATING
C2978 INVX2_39/Y 0 12.184021f **FLOATING
C2979 AOI22X1_74/A 0 14.501282f **FLOATING
C2980 AOI22X1_41/a_2_54# 0 6.66f **FLOATING
C2981 AOI22X1_30/a_2_54# 0 6.66f **FLOATING
C2982 NAND2X1_98/Y 0 6.87006f **FLOATING
C2983 NAND2X1_87/Y 0 6.87006f **FLOATING
C2984 OAI21X1_58/C 0 6.87006f **FLOATING
C2985 OAI21X1_76/B 0 10.49256f **FLOATING
C2986 OAI21X1_89/C 0 18.502602f **FLOATING
C2987 NOR2X1_43/A 0 7.25151f **FLOATING
C2988 AOI22X1_0/a_2_54# 0 6.66f **FLOATING
C2989 MUX2X1_28/a_2_10# 0 6.0456f **FLOATING
C2990 DFFNEGX1_130/a_66_6# 0 6.40992f **FLOATING
C2991 DFFNEGX1_130/a_23_6# 0 6.85692f **FLOATING
C2992 DFFNEGX1_130/a_34_4# 0 4.93023f **FLOATING
C2993 DFFNEGX1_130/a_2_6# 0 9.33504f **FLOATING
C2994 DFFNEGX1_141/a_66_6# 0 6.40992f **FLOATING
C2995 out_alu 0 19.745338f **FLOATING
C2996 DFFNEGX1_141/a_23_6# 0 6.85692f **FLOATING
C2997 DFFNEGX1_141/a_34_4# 0 4.93023f **FLOATING
C2998 DFFNEGX1_141/a_2_6# 0 9.33504f **FLOATING
C2999 OAI21X1_157/Y 0 13.775221f **FLOATING
C3000 MUX2X1_17/Y 0 10.32702f **FLOATING
C3001 MUX2X1_17/a_2_10# 0 6.0456f **FLOATING
C3002 AND2X2_5/a_2_6# 0 6.03567f **FLOATING
C3003 HAX1_9/a_38_6# 0 2.442f **FLOATING
C3004 HAX1_9/a_41_74# 0 5.99325f **FLOATING
C3005 HAX1_9/a_2_74# 0 7.65318f **FLOATING
C3006 DFFNEGX1_62/a_66_6# 0 6.40992f **FLOATING
C3007 DFFNEGX1_62/a_23_6# 0 6.85692f **FLOATING
C3008 DFFNEGX1_62/a_34_4# 0 4.93023f **FLOATING
C3009 DFFNEGX1_62/a_2_6# 0 9.33504f **FLOATING
C3010 DFFNEGX1_73/a_66_6# 0 6.40992f **FLOATING
C3011 DFFNEGX1_73/a_23_6# 0 6.85692f **FLOATING
C3012 DFFNEGX1_73/a_34_4# 0 4.93023f **FLOATING
C3013 DFFNEGX1_73/a_2_6# 0 9.33504f **FLOATING
C3014 DFFNEGX1_84/a_66_6# 0 6.40992f **FLOATING
C3015 DFFNEGX1_84/a_23_6# 0 6.85692f **FLOATING
C3016 DFFNEGX1_84/a_34_4# 0 4.93023f **FLOATING
C3017 DFFNEGX1_84/a_2_6# 0 9.33504f **FLOATING
C3018 DFFNEGX1_95/a_66_6# 0 6.40992f **FLOATING
C3019 DFFNEGX1_95/a_23_6# 0 6.85692f **FLOATING
C3020 DFFNEGX1_95/a_34_4# 0 4.93023f **FLOATING
C3021 DFFNEGX1_95/a_2_6# 0 9.33504f **FLOATING
C3022 DFFNEGX1_40/a_66_6# 0 6.40992f **FLOATING
C3023 DFFNEGX1_40/a_23_6# 0 6.85692f **FLOATING
C3024 DFFNEGX1_40/a_34_4# 0 4.93023f **FLOATING
C3025 DFFNEGX1_40/a_2_6# 0 9.33504f **FLOATING
C3026 DFFNEGX1_51/a_66_6# 0 6.40992f **FLOATING
C3027 out_temp_decoded[15] 0 19.35801f **FLOATING
C3028 DFFNEGX1_51/a_23_6# 0 6.85692f **FLOATING
C3029 DFFNEGX1_51/a_34_4# 0 4.93023f **FLOATING
C3030 DFFNEGX1_51/a_2_6# 0 9.33504f **FLOATING
C3031 OAI21X1_97/Y 0 11.97402f **FLOATING
