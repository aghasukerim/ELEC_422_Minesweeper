magic
tech scmos
timestamp 1710899220
<< metal1 >>
rect 14 2607 2730 2627
rect 38 2583 2706 2603
rect 38 2567 2706 2573
rect 156 2533 165 2536
rect 204 2533 220 2536
rect 380 2533 389 2536
rect 508 2533 524 2536
rect 684 2533 693 2536
rect 812 2533 821 2536
rect 1004 2533 1013 2536
rect 1132 2533 1141 2536
rect 1276 2533 1285 2536
rect 1484 2533 1493 2536
rect 1612 2533 1621 2536
rect 1804 2533 1820 2536
rect 1946 2533 1956 2536
rect 2138 2533 2156 2536
rect 2178 2533 2188 2536
rect 108 2523 125 2526
rect 130 2523 140 2526
rect 266 2503 269 2533
rect 1170 2526 1173 2533
rect 1986 2526 1989 2533
rect 338 2523 348 2526
rect 466 2523 476 2526
rect 642 2523 652 2526
rect 770 2523 780 2526
rect 836 2523 845 2526
rect 884 2523 893 2526
rect 332 2513 341 2516
rect 420 2513 429 2516
rect 460 2513 469 2516
rect 636 2513 645 2516
rect 724 2513 733 2516
rect 764 2513 773 2516
rect 898 2503 901 2525
rect 962 2523 972 2526
rect 1090 2523 1100 2526
rect 1138 2523 1156 2526
rect 1162 2523 1173 2526
rect 1204 2523 1229 2526
rect 1300 2523 1309 2526
rect 1442 2523 1452 2526
rect 1498 2523 1508 2526
rect 1570 2523 1580 2526
rect 1636 2523 1645 2526
rect 1690 2523 1700 2526
rect 1762 2523 1772 2526
rect 1810 2523 1828 2526
rect 1868 2523 1893 2526
rect 1930 2523 1940 2526
rect 1980 2523 1989 2526
rect 2058 2523 2076 2526
rect 2138 2523 2148 2526
rect 2404 2523 2421 2526
rect 2588 2523 2605 2526
rect 956 2513 965 2516
rect 1084 2513 1093 2516
rect 1162 2515 1165 2523
rect 2138 2516 2141 2523
rect 1436 2513 1445 2516
rect 1524 2513 1533 2516
rect 1564 2513 1573 2516
rect 1756 2513 1765 2516
rect 2012 2513 2021 2516
rect 2132 2513 2141 2516
rect 14 2467 2730 2473
rect 100 2413 133 2416
rect 140 2413 157 2416
rect 178 2413 188 2416
rect 260 2413 269 2416
rect 284 2413 293 2416
rect 298 2413 324 2416
rect 356 2413 365 2416
rect 402 2413 412 2416
rect 418 2406 421 2425
rect 1570 2423 1605 2426
rect 1620 2423 1629 2426
rect 1660 2423 1677 2426
rect 2228 2423 2237 2426
rect 2268 2423 2277 2426
rect 2548 2423 2557 2426
rect 468 2413 501 2416
rect 508 2413 517 2416
rect 570 2413 596 2416
rect 628 2413 637 2416
rect 652 2413 685 2416
rect 692 2413 709 2416
rect 740 2413 765 2416
rect 772 2413 781 2416
rect 844 2413 861 2416
rect 876 2413 885 2416
rect 890 2413 900 2416
rect 932 2413 941 2416
rect 980 2413 1004 2416
rect 1052 2413 1061 2416
rect 1076 2413 1093 2416
rect 1124 2413 1149 2416
rect 1194 2413 1212 2416
rect 1244 2413 1268 2416
rect 1282 2413 1333 2416
rect 1348 2413 1357 2416
rect 1404 2413 1429 2416
rect 1436 2413 1477 2416
rect 1564 2413 1597 2416
rect 1602 2415 1605 2423
rect 2274 2416 2277 2423
rect 2554 2416 2557 2423
rect 1666 2413 1684 2416
rect 1852 2413 1877 2416
rect 1914 2413 1924 2416
rect 1964 2413 1973 2416
rect 124 2403 132 2406
rect 220 2403 252 2406
rect 266 2403 276 2406
rect 356 2403 397 2406
rect 418 2403 436 2406
rect 490 2403 500 2406
rect 564 2403 589 2406
rect 698 2403 708 2406
rect 820 2403 836 2406
rect 850 2403 868 2406
rect 980 2403 989 2406
rect 1010 2403 1044 2406
rect 1058 2395 1061 2413
rect 1074 2403 1092 2406
rect 1188 2403 1205 2406
rect 1244 2403 1253 2406
rect 1274 2403 1300 2406
rect 1330 2395 1333 2413
rect 1594 2407 1597 2413
rect 1970 2407 1973 2413
rect 2186 2413 2212 2416
rect 2274 2413 2284 2416
rect 2396 2413 2405 2416
rect 2474 2413 2492 2416
rect 2554 2413 2564 2416
rect 2602 2413 2612 2416
rect 1340 2403 1365 2406
rect 1420 2403 1428 2406
rect 1442 2403 1476 2406
rect 1524 2403 1556 2406
rect 1716 2403 1732 2406
rect 2186 2403 2189 2413
rect 2402 2407 2405 2413
rect 2314 2403 2324 2406
rect 2338 2403 2372 2406
rect 2554 2403 2572 2406
rect 2594 2403 2604 2406
rect 38 2367 2706 2373
rect 74 2326 77 2346
rect 474 2343 484 2346
rect 138 2333 148 2336
rect 274 2333 300 2336
rect 306 2333 316 2336
rect 412 2333 421 2336
rect 442 2333 460 2336
rect 74 2323 132 2326
rect 138 2315 141 2333
rect 180 2323 221 2326
rect 306 2325 309 2333
rect 474 2326 477 2343
rect 1938 2336 1941 2346
rect 498 2333 508 2336
rect 684 2333 693 2336
rect 714 2333 748 2336
rect 906 2333 916 2336
rect 964 2333 981 2336
rect 1372 2333 1389 2336
rect 1434 2333 1444 2336
rect 1458 2333 1492 2336
rect 1540 2333 1548 2336
rect 1562 2333 1580 2336
rect 1628 2333 1637 2336
rect 1692 2333 1709 2336
rect 1738 2333 1756 2336
rect 1898 2333 2012 2336
rect 2034 2333 2044 2336
rect 2058 2333 2068 2336
rect 2234 2333 2260 2336
rect 2282 2333 2292 2336
rect 2554 2333 2564 2336
rect 554 2326 557 2333
rect 348 2323 373 2326
rect 412 2323 436 2326
rect 468 2323 477 2326
rect 500 2323 509 2326
rect 538 2323 557 2326
rect 620 2323 645 2326
rect 684 2323 708 2326
rect 756 2323 781 2326
rect 948 2323 973 2326
rect 1316 2323 1333 2326
rect 1378 2323 1396 2326
rect 1428 2323 1452 2326
rect 1524 2323 1549 2326
rect 1556 2323 1573 2326
rect 1650 2323 1660 2326
rect 1692 2323 1701 2326
rect 1754 2323 1764 2326
rect 2036 2323 2045 2326
rect 2052 2323 2069 2326
rect 2138 2323 2164 2326
rect 2242 2323 2252 2326
rect 2300 2323 2317 2326
rect 2514 2323 2524 2326
rect 2242 2316 2245 2323
rect 2514 2316 2517 2323
rect 1780 2313 1789 2316
rect 2092 2313 2101 2316
rect 2180 2313 2189 2316
rect 2220 2313 2245 2316
rect 2508 2313 2517 2316
rect 14 2267 2730 2273
rect 676 2223 685 2226
rect 716 2223 725 2226
rect 1748 2223 1757 2226
rect 1970 2223 1981 2226
rect 2388 2223 2397 2226
rect 2468 2223 2477 2226
rect 2508 2223 2517 2226
rect 100 2213 125 2216
rect 458 2213 477 2216
rect 850 2213 860 2216
rect 1418 2213 1445 2216
rect 1500 2213 1524 2216
rect 1546 2213 1572 2216
rect 1684 2213 1725 2216
rect 1852 2213 1877 2216
rect 1964 2213 1973 2216
rect 1978 2215 1981 2223
rect 2514 2216 2517 2223
rect 2188 2213 2213 2216
rect 2300 2213 2309 2216
rect 474 2207 477 2213
rect 306 2203 316 2206
rect 418 2203 428 2206
rect 476 2203 485 2206
rect 722 2203 732 2206
rect 1210 2203 1236 2206
rect 1442 2195 1445 2213
rect 1970 2207 1973 2213
rect 2306 2207 2309 2213
rect 2354 2206 2357 2214
rect 2442 2213 2452 2216
rect 2514 2213 2524 2216
rect 2596 2213 2621 2216
rect 2658 2213 2668 2216
rect 1500 2203 1509 2206
rect 1604 2203 1629 2206
rect 1690 2203 1724 2206
rect 1930 2203 1940 2206
rect 2266 2203 2276 2206
rect 2322 2203 2332 2206
rect 2354 2203 2364 2206
rect 38 2167 2706 2173
rect 650 2136 653 2146
rect 658 2143 684 2146
rect 1050 2143 1076 2146
rect 1090 2136 1093 2146
rect 98 2133 108 2136
rect 226 2133 236 2136
rect 650 2133 692 2136
rect 698 2133 716 2136
rect 1084 2133 1093 2136
rect 1194 2133 1220 2136
rect 522 2126 525 2133
rect 1250 2126 1253 2144
rect 1260 2133 1285 2136
rect 1426 2133 1436 2136
rect 1556 2133 1573 2136
rect 1580 2133 1597 2136
rect 1642 2133 1652 2136
rect 1666 2133 1676 2136
rect 1724 2133 1732 2136
rect 1916 2133 1933 2136
rect 2138 2133 2148 2136
rect 2346 2133 2388 2136
rect 498 2123 525 2126
rect 1244 2123 1253 2126
rect 1282 2123 1285 2133
rect 1938 2126 1941 2133
rect 2178 2126 2181 2133
rect 1348 2123 1381 2126
rect 1420 2123 1444 2126
rect 1500 2123 1517 2126
rect 1642 2123 1660 2126
rect 1796 2123 1821 2126
rect 1858 2123 1884 2126
rect 1924 2123 1941 2126
rect 2060 2123 2085 2126
rect 2172 2123 2181 2126
rect 2250 2123 2284 2126
rect 2396 2123 2405 2126
rect 1148 2113 1157 2116
rect 1188 2113 1205 2116
rect 1964 2113 1973 2116
rect 14 2067 2730 2073
rect 492 2023 501 2026
rect 98 2006 101 2016
rect 252 2013 268 2016
rect 692 2013 701 2016
rect 746 2013 756 2016
rect 980 2013 989 2016
rect 1010 2013 1020 2016
rect 1186 2013 1221 2016
rect 1260 2013 1285 2016
rect 1316 2013 1325 2016
rect 1332 2013 1349 2016
rect 1378 2013 1388 2016
rect 1436 2013 1453 2016
rect 1498 2013 1516 2016
rect 1532 2013 1549 2016
rect 1852 2013 1877 2016
rect 1914 2013 1924 2016
rect 1964 2013 1973 2016
rect 2324 2013 2333 2016
rect 2450 2015 2453 2036
rect 2508 2023 2517 2026
rect 2514 2016 2517 2023
rect 2514 2013 2524 2016
rect 1970 2007 1973 2013
rect 98 2003 244 2006
rect 498 2003 516 2006
rect 644 2003 653 2006
rect 674 2003 684 2006
rect 708 2003 717 2006
rect 738 2003 748 2006
rect 818 2003 844 2006
rect 850 2003 868 2006
rect 882 2003 892 2006
rect 906 2003 916 2006
rect 946 2003 972 2006
rect 978 2003 996 2006
rect 1044 2003 1060 2006
rect 1130 2003 1148 2006
rect 1154 2003 1172 2006
rect 1572 2003 1589 2006
rect 1956 2003 1965 2006
rect 2074 2003 2084 2006
rect 2266 2003 2284 2006
rect 2306 2003 2316 2006
rect 2514 2003 2532 2006
rect 2554 2003 2564 2006
rect 218 1993 236 1996
rect 690 1993 700 1996
rect 738 1993 741 2003
rect 826 1993 836 1996
rect 850 1993 860 1996
rect 874 1993 884 1996
rect 946 1993 964 1996
rect 978 1993 988 1996
rect 1026 1993 1036 1996
rect 1154 1993 1164 1996
rect 2074 1993 2077 2003
rect 38 1967 2706 1973
rect 1562 1943 1580 1946
rect 250 1933 260 1936
rect 274 1933 284 1936
rect 426 1933 436 1936
rect 450 1933 468 1936
rect 474 1933 492 1936
rect 658 1933 668 1936
rect 1364 1933 1373 1936
rect 1378 1933 1404 1936
rect 1418 1933 1428 1936
rect 1508 1933 1525 1936
rect 1570 1933 1613 1936
rect 1634 1933 1644 1936
rect 2138 1933 2172 1936
rect 2194 1933 2204 1936
rect 642 1926 645 1933
rect 1314 1926 1317 1933
rect 476 1923 485 1926
rect 500 1923 517 1926
rect 564 1923 589 1926
rect 620 1923 645 1926
rect 652 1923 669 1926
rect 690 1923 716 1926
rect 804 1923 829 1926
rect 890 1923 908 1926
rect 972 1923 997 1926
rect 1028 1923 1037 1926
rect 1058 1923 1076 1926
rect 1114 1923 1132 1926
rect 1154 1923 1164 1926
rect 1228 1923 1253 1926
rect 1284 1923 1317 1926
rect 1324 1923 1341 1926
rect 1412 1923 1429 1926
rect 890 1915 893 1923
rect 1058 1915 1061 1923
rect 1114 1916 1117 1923
rect 1084 1913 1117 1916
rect 1364 1913 1381 1916
rect 1522 1906 1525 1933
rect 1570 1923 1581 1926
rect 1602 1923 1612 1926
rect 1634 1925 1637 1933
rect 1652 1923 1669 1926
rect 2020 1923 2045 1926
rect 2082 1923 2100 1926
rect 2196 1923 2205 1926
rect 2212 1923 2237 1926
rect 2276 1923 2285 1926
rect 2498 1923 2508 1926
rect 2546 1923 2549 1933
rect 2658 1923 2668 1926
rect 1570 1916 1573 1923
rect 2498 1916 2501 1923
rect 1532 1913 1541 1916
rect 1556 1913 1573 1916
rect 2452 1913 2461 1916
rect 2492 1913 2501 1916
rect 1522 1903 1548 1906
rect 14 1867 2730 1873
rect 1538 1833 1556 1836
rect 1642 1833 1660 1836
rect 1002 1816 1005 1825
rect 1026 1816 1029 1825
rect 500 1813 525 1816
rect 556 1813 605 1816
rect 612 1813 629 1816
rect 650 1813 668 1816
rect 724 1813 749 1816
rect 780 1813 789 1816
rect 804 1813 821 1816
rect 842 1813 860 1816
rect 908 1813 933 1816
rect 1002 1813 1020 1816
rect 1026 1813 1044 1816
rect 1058 1813 1076 1816
rect 1186 1813 1212 1816
rect 1226 1813 1244 1816
rect 1258 1813 1276 1816
rect 1282 1813 1292 1816
rect 602 1807 605 1813
rect 786 1806 789 1813
rect 1298 1806 1301 1825
rect 1540 1823 1549 1826
rect 1588 1823 1597 1826
rect 1668 1823 1677 1826
rect 2404 1823 2413 1826
rect 2524 1823 2533 1826
rect 1594 1816 1597 1823
rect 1674 1816 1677 1823
rect 2530 1816 2533 1823
rect 1306 1813 1316 1816
rect 1412 1813 1421 1816
rect 1436 1813 1461 1816
rect 1468 1813 1477 1816
rect 1508 1813 1517 1816
rect 1594 1813 1605 1816
rect 1612 1813 1621 1816
rect 1628 1813 1637 1816
rect 1674 1813 1685 1816
rect 1692 1813 1701 1816
rect 1708 1813 1725 1816
rect 1866 1813 1884 1816
rect 1900 1813 1908 1816
rect 2164 1813 2189 1816
rect 2260 1813 2285 1816
rect 2322 1813 2332 1816
rect 2372 1813 2381 1816
rect 2458 1813 2468 1816
rect 2530 1813 2540 1816
rect 2612 1813 2637 1816
rect 618 1803 628 1806
rect 786 1803 796 1806
rect 810 1803 820 1806
rect 1298 1803 1308 1806
rect 1410 1803 1428 1806
rect 1434 1803 1444 1806
rect 1474 1795 1477 1813
rect 1514 1795 1517 1813
rect 1602 1807 1605 1813
rect 1618 1807 1621 1813
rect 1634 1803 1637 1813
rect 2378 1807 2381 1813
rect 1674 1803 1684 1806
rect 1714 1803 1724 1806
rect 1748 1803 1757 1806
rect 2530 1803 2548 1806
rect 210 1783 421 1786
rect 38 1767 2706 1773
rect 1210 1736 1213 1756
rect 482 1733 508 1736
rect 546 1733 555 1736
rect 620 1733 629 1736
rect 714 1733 732 1736
rect 922 1733 932 1736
rect 956 1733 965 1736
rect 986 1733 996 1736
rect 1020 1733 1029 1736
rect 1034 1733 1044 1736
rect 1106 1733 1124 1736
rect 1210 1733 1220 1736
rect 1250 1733 1260 1736
rect 1314 1733 1324 1736
rect 1338 1733 1364 1736
rect 1404 1733 1412 1736
rect 1498 1733 1508 1736
rect 1522 1733 1532 1736
rect 1546 1733 1556 1736
rect 1612 1733 1621 1736
rect 1746 1733 1756 1736
rect 1780 1733 1789 1736
rect 2186 1733 2196 1736
rect 2530 1733 2548 1736
rect 754 1726 757 1733
rect 130 1723 196 1726
rect 250 1723 268 1726
rect 354 1723 364 1726
rect 442 1723 452 1726
rect 594 1723 604 1726
rect 626 1723 644 1726
rect 714 1723 740 1726
rect 754 1723 765 1726
rect 772 1723 789 1726
rect 844 1723 869 1726
rect 916 1723 933 1726
rect 980 1723 997 1726
rect 1042 1723 1052 1726
rect 1058 1723 1068 1726
rect 1074 1723 1084 1726
rect 1090 1723 1100 1726
rect 1194 1723 1204 1726
rect 1210 1723 1228 1726
rect 1250 1723 1261 1726
rect 1290 1723 1308 1726
rect 1322 1723 1332 1726
rect 1346 1723 1388 1726
rect 1492 1723 1509 1726
rect 1516 1723 1533 1726
rect 1540 1723 1564 1726
rect 1578 1723 1596 1726
rect 1610 1723 1645 1726
rect 1674 1723 1692 1726
rect 1724 1723 1733 1726
rect 1740 1723 1757 1726
rect 1924 1723 1949 1726
rect 2018 1723 2028 1726
rect 2034 1723 2044 1726
rect 2106 1723 2124 1726
rect 250 1716 253 1723
rect 1250 1716 1253 1723
rect 2186 1716 2189 1733
rect 2378 1726 2381 1733
rect 2260 1723 2285 1726
rect 2322 1723 2332 1726
rect 2372 1723 2381 1726
rect 2450 1723 2468 1726
rect 2530 1723 2540 1726
rect 2530 1716 2533 1723
rect 236 1713 253 1716
rect 1244 1713 1253 1716
rect 1284 1713 1301 1716
rect 1340 1713 1357 1716
rect 2060 1713 2069 1716
rect 2100 1713 2125 1716
rect 2180 1713 2189 1716
rect 2404 1713 2413 1716
rect 2524 1713 2533 1716
rect 1354 1693 1357 1713
rect 14 1667 2730 1673
rect 260 1623 277 1626
rect 706 1616 709 1625
rect 866 1616 869 1625
rect 1394 1616 1397 1625
rect 1618 1616 1621 1625
rect 338 1613 356 1616
rect 442 1613 460 1616
rect 514 1613 524 1616
rect 554 1613 580 1616
rect 610 1613 644 1616
rect 674 1613 692 1616
rect 706 1613 733 1616
rect 780 1613 805 1616
rect 866 1613 884 1616
rect 948 1613 973 1616
rect 1044 1613 1069 1616
rect 1100 1613 1109 1616
rect 1116 1613 1133 1616
rect 1154 1613 1172 1616
rect 1178 1613 1188 1616
rect 1250 1613 1268 1616
rect 1282 1613 1300 1616
rect 1322 1613 1332 1616
rect 1346 1613 1364 1616
rect 1394 1613 1412 1616
rect 1530 1613 1540 1616
rect 1554 1613 1572 1616
rect 1618 1613 1636 1616
rect 1650 1613 1668 1616
rect 1690 1613 1700 1616
rect 1714 1613 1732 1616
rect 1780 1613 1789 1616
rect 1796 1613 1805 1616
rect 380 1603 397 1606
rect 484 1603 501 1606
rect 506 1603 516 1606
rect 554 1603 572 1606
rect 674 1603 684 1606
rect 1106 1605 1109 1613
rect 1122 1603 1132 1606
rect 1348 1603 1356 1606
rect 1748 1603 1772 1606
rect 1810 1605 1813 1636
rect 2138 1625 2141 1636
rect 1826 1616 1829 1623
rect 1826 1613 1837 1616
rect 2116 1613 2133 1616
rect 2204 1613 2237 1616
rect 2252 1613 2269 1616
rect 1834 1605 1837 1613
rect 1860 1603 1869 1606
rect 1986 1603 2004 1606
rect 2058 1603 2084 1606
rect 2170 1603 2180 1606
rect 506 1596 509 1603
rect 490 1593 509 1596
rect 2234 1595 2237 1613
rect 2554 1606 2557 1616
rect 2610 1613 2620 1616
rect 2258 1603 2276 1606
rect 2554 1603 2612 1606
rect 2482 1583 2557 1586
rect 38 1567 2706 1573
rect 770 1536 773 1545
rect 146 1533 156 1536
rect 172 1533 181 1536
rect 364 1533 381 1536
rect 490 1533 516 1536
rect 724 1533 756 1536
rect 770 1533 788 1536
rect 810 1533 820 1536
rect 946 1533 956 1536
rect 1250 1533 1260 1536
rect 1506 1533 1516 1536
rect 1714 1533 1724 1536
rect 2194 1533 2220 1536
rect 2322 1533 2332 1536
rect 2618 1533 2636 1536
rect 186 1526 189 1533
rect 930 1526 933 1533
rect 130 1523 148 1526
rect 180 1523 189 1526
rect 378 1523 404 1526
rect 514 1523 524 1526
rect 562 1523 580 1526
rect 610 1523 619 1526
rect 642 1523 668 1526
rect 698 1523 707 1526
rect 722 1523 747 1526
rect 818 1523 828 1526
rect 868 1523 893 1526
rect 924 1523 933 1526
rect 308 1513 325 1516
rect 636 1513 645 1516
rect 724 1513 733 1516
rect 946 1515 949 1533
rect 1082 1526 1085 1533
rect 1234 1526 1237 1533
rect 1020 1523 1045 1526
rect 1076 1523 1085 1526
rect 1092 1523 1109 1526
rect 1172 1523 1197 1526
rect 1228 1523 1237 1526
rect 1244 1523 1261 1526
rect 1282 1523 1300 1526
rect 1330 1523 1340 1526
rect 1354 1523 1372 1526
rect 1500 1523 1517 1526
rect 1538 1523 1556 1526
rect 1612 1523 1621 1526
rect 1708 1523 1725 1526
rect 1874 1523 1892 1526
rect 1972 1523 1989 1526
rect 1354 1515 1357 1523
rect 1874 1515 1877 1523
rect 2194 1516 2197 1533
rect 2330 1523 2340 1526
rect 2498 1523 2508 1526
rect 2618 1523 2628 1526
rect 2498 1516 2501 1523
rect 2618 1516 2621 1523
rect 2148 1513 2157 1516
rect 2188 1513 2197 1516
rect 2492 1513 2501 1516
rect 2612 1513 2621 1516
rect 14 1467 2730 1473
rect 858 1453 877 1456
rect 172 1423 181 1426
rect 212 1423 221 1426
rect 402 1416 405 1426
rect 98 1413 156 1416
rect 268 1413 277 1416
rect 402 1413 427 1416
rect 434 1406 437 1425
rect 524 1423 534 1426
rect 442 1413 453 1416
rect 522 1413 540 1416
rect 402 1403 420 1406
rect 434 1403 445 1406
rect 450 1405 453 1413
rect 546 1406 549 1425
rect 852 1423 877 1426
rect 874 1416 877 1423
rect 1346 1416 1349 1425
rect 564 1413 581 1416
rect 602 1413 612 1416
rect 626 1413 644 1416
rect 674 1413 692 1416
rect 722 1413 739 1416
rect 490 1403 508 1406
rect 522 1403 531 1406
rect 546 1403 555 1406
rect 578 1405 581 1413
rect 778 1406 781 1414
rect 804 1413 836 1416
rect 874 1413 892 1416
rect 1060 1413 1085 1416
rect 1116 1413 1133 1416
rect 1140 1413 1157 1416
rect 1252 1413 1277 1416
rect 1314 1413 1332 1416
rect 1346 1413 1364 1416
rect 1556 1413 1565 1416
rect 594 1403 604 1406
rect 756 1403 781 1406
rect 802 1403 828 1406
rect 852 1403 877 1406
rect 908 1403 1005 1406
rect 1130 1405 1133 1413
rect 1578 1406 1581 1425
rect 1586 1413 1596 1416
rect 1770 1413 1780 1416
rect 2044 1413 2053 1416
rect 2058 1413 2108 1416
rect 2204 1413 2229 1416
rect 2308 1413 2333 1416
rect 2444 1413 2469 1416
rect 2506 1413 2516 1416
rect 2564 1413 2589 1416
rect 2626 1413 2636 1416
rect 1146 1403 1156 1406
rect 1578 1403 1588 1406
rect 1612 1403 1629 1406
rect 804 1393 821 1396
rect 38 1367 2706 1373
rect 738 1353 749 1356
rect 306 1343 316 1346
rect 402 1336 405 1346
rect 538 1336 541 1345
rect 124 1333 133 1336
rect 402 1333 427 1336
rect 482 1333 524 1336
rect 538 1333 573 1336
rect 708 1333 717 1336
rect 724 1333 741 1336
rect 426 1326 429 1333
rect 746 1326 749 1353
rect 834 1336 837 1356
rect 2074 1343 2124 1346
rect 820 1333 845 1336
rect 874 1333 885 1336
rect 908 1333 917 1336
rect 922 1333 940 1336
rect 962 1333 972 1336
rect 1026 1333 1044 1336
rect 1106 1333 1116 1336
rect 1164 1333 1172 1336
rect 1186 1333 1196 1336
rect 1348 1333 1356 1336
rect 1554 1333 1564 1336
rect 1684 1333 1692 1336
rect 1956 1333 1981 1336
rect 2034 1333 2044 1336
rect 2074 1333 2132 1336
rect 2154 1333 2180 1336
rect 2234 1333 2252 1336
rect 2314 1333 2324 1336
rect 2442 1333 2516 1336
rect 2538 1333 2548 1336
rect 842 1326 845 1333
rect 882 1326 885 1333
rect 1258 1326 1261 1333
rect 1618 1326 1621 1333
rect 1634 1326 1637 1333
rect 2074 1326 2077 1333
rect 2370 1326 2373 1333
rect 156 1323 165 1326
rect 196 1323 213 1326
rect 276 1323 309 1326
rect 380 1323 429 1326
rect 436 1323 445 1326
rect 452 1323 461 1326
rect 570 1323 587 1326
rect 588 1323 597 1326
rect 618 1323 661 1326
rect 692 1323 717 1326
rect 746 1323 757 1326
rect 788 1323 805 1326
rect 964 1323 973 1326
rect 980 1323 997 1326
rect 1002 1323 1012 1326
rect 1018 1323 1036 1326
rect 1074 1323 1100 1326
rect 1140 1323 1173 1326
rect 1180 1323 1197 1326
rect 1226 1323 1261 1326
rect 1324 1323 1357 1326
rect 1394 1323 1404 1326
rect 1436 1323 1477 1326
rect 1530 1323 1548 1326
rect 1594 1323 1621 1326
rect 1628 1323 1637 1326
rect 1666 1323 1700 1326
rect 1850 1323 1916 1326
rect 1962 1323 2012 1326
rect 2068 1323 2077 1326
rect 2148 1323 2181 1326
rect 2250 1323 2260 1326
rect 2276 1323 2285 1326
rect 2290 1323 2308 1326
rect 2348 1323 2373 1326
rect 2556 1323 2573 1326
rect 460 1313 469 1316
rect 618 1315 621 1323
rect 14 1267 2730 1273
rect 402 1216 405 1226
rect 1106 1216 1109 1218
rect 1514 1216 1517 1246
rect 2218 1233 2228 1236
rect 1764 1223 1773 1226
rect 1802 1216 1805 1225
rect 1986 1216 1989 1225
rect 2404 1223 2413 1226
rect 2444 1223 2453 1226
rect 2524 1223 2533 1226
rect 2450 1216 2453 1223
rect 116 1213 181 1216
rect 202 1213 213 1216
rect 316 1213 325 1216
rect 402 1213 413 1216
rect 450 1213 459 1216
rect 522 1213 533 1216
rect 578 1213 595 1216
rect 730 1213 739 1216
rect 754 1213 765 1216
rect 202 1207 205 1213
rect 410 1207 413 1213
rect 522 1207 525 1213
rect 754 1207 757 1213
rect 818 1206 821 1214
rect 1028 1213 1037 1216
rect 1044 1213 1053 1216
rect 1074 1213 1084 1216
rect 1098 1213 1109 1216
rect 1130 1213 1141 1216
rect 1204 1213 1237 1216
rect 1324 1213 1365 1216
rect 1388 1213 1420 1216
rect 1514 1213 1525 1216
rect 1554 1213 1573 1216
rect 1588 1213 1597 1216
rect 1676 1213 1685 1216
rect 1802 1213 1820 1216
rect 1954 1213 1965 1216
rect 1986 1213 2004 1216
rect 2146 1213 2164 1216
rect 1098 1207 1101 1213
rect 1130 1207 1133 1213
rect 1362 1207 1365 1213
rect 1522 1207 1525 1213
rect 1570 1207 1573 1213
rect 1954 1207 1957 1213
rect 2258 1206 2261 1214
rect 2266 1213 2276 1216
rect 2450 1213 2460 1216
rect 2498 1213 2508 1216
rect 2650 1213 2669 1216
rect 2666 1207 2669 1213
rect 74 1203 92 1206
rect 140 1203 149 1206
rect 236 1203 253 1206
rect 402 1203 412 1206
rect 490 1203 499 1206
rect 722 1203 732 1206
rect 778 1203 796 1206
rect 818 1203 853 1206
rect 890 1203 900 1206
rect 916 1203 933 1206
rect 996 1203 1020 1206
rect 1060 1203 1076 1206
rect 1250 1203 1260 1206
rect 1450 1203 1460 1206
rect 1650 1203 1668 1206
rect 1724 1203 1740 1206
rect 1764 1203 1780 1206
rect 2170 1203 2188 1206
rect 2242 1203 2252 1206
rect 2258 1203 2268 1206
rect 2450 1203 2468 1206
rect 2570 1203 2588 1206
rect 316 1193 333 1196
rect 402 1183 405 1203
rect 778 1193 781 1203
rect 38 1167 2706 1173
rect 82 1143 108 1146
rect 282 1143 333 1146
rect 258 1133 268 1136
rect 172 1123 205 1126
rect 258 1125 261 1133
rect 282 1126 285 1143
rect 386 1136 389 1146
rect 786 1143 804 1146
rect 818 1143 845 1146
rect 890 1143 908 1146
rect 818 1136 821 1143
rect 978 1136 981 1145
rect 386 1133 396 1136
rect 450 1133 474 1136
rect 508 1133 541 1136
rect 636 1133 653 1136
rect 722 1133 739 1136
rect 764 1133 797 1136
rect 812 1133 821 1136
rect 826 1133 860 1136
rect 882 1133 916 1136
rect 922 1133 957 1136
rect 978 1133 988 1136
rect 1002 1133 1028 1136
rect 1194 1133 1204 1136
rect 266 1123 285 1126
rect 378 1123 402 1126
rect 434 1123 483 1126
rect 546 1123 555 1126
rect 586 1123 612 1126
rect 650 1113 653 1133
rect 730 1123 747 1126
rect 842 1123 852 1126
rect 882 1125 885 1133
rect 954 1125 957 1133
rect 1258 1126 1261 1135
rect 1298 1133 1308 1136
rect 1362 1126 1365 1135
rect 1458 1133 1468 1136
rect 1588 1133 1605 1136
rect 1682 1126 1685 1135
rect 1708 1133 1725 1136
rect 1802 1126 1805 1135
rect 1010 1123 1020 1126
rect 1132 1123 1157 1126
rect 1228 1123 1261 1126
rect 1332 1123 1365 1126
rect 1388 1123 1420 1126
rect 1500 1123 1524 1126
rect 1556 1123 1564 1126
rect 1660 1123 1685 1126
rect 1740 1123 1749 1126
rect 1764 1123 1805 1126
rect 1826 1126 1829 1135
rect 2060 1133 2069 1136
rect 1826 1123 1837 1126
rect 2002 1123 2044 1126
rect 2282 1116 2285 1135
rect 2292 1123 2325 1126
rect 2596 1123 2621 1126
rect 2658 1123 2668 1126
rect 1708 1113 1717 1116
rect 1828 1113 1837 1116
rect 2242 1113 2252 1116
rect 2276 1113 2285 1116
rect 2300 1113 2309 1116
rect 1834 1103 1837 1113
rect 14 1067 2730 1073
rect 330 1053 349 1056
rect 2426 1033 2460 1036
rect 538 1023 557 1026
rect 116 1013 180 1016
rect 242 1013 284 1016
rect 354 1013 363 1016
rect 450 1013 468 1016
rect 74 1003 92 1006
rect 140 1003 157 1006
rect 324 1003 333 1006
rect 338 1003 354 1006
rect 450 1003 459 1006
rect 154 993 157 1003
rect 538 996 541 1023
rect 658 1016 661 1024
rect 1170 1016 1173 1025
rect 1346 1016 1349 1025
rect 2580 1023 2589 1026
rect 546 1013 564 1016
rect 570 1006 573 1016
rect 578 1013 587 1016
rect 602 1013 626 1016
rect 642 1013 652 1016
rect 658 1013 683 1016
rect 690 1013 700 1016
rect 738 1013 747 1016
rect 770 1013 788 1016
rect 858 1013 868 1016
rect 882 1013 893 1016
rect 956 1013 965 1016
rect 882 1006 885 1013
rect 570 1003 580 1006
rect 602 1003 619 1006
rect 666 1003 675 1006
rect 698 1003 707 1006
rect 730 1003 739 1006
rect 764 1003 781 1006
rect 906 1003 916 1006
rect 962 1005 965 1013
rect 994 1006 997 1014
rect 1052 1013 1068 1016
rect 1098 1013 1108 1016
rect 1170 1013 1188 1016
rect 1252 1013 1277 1016
rect 1314 1013 1332 1016
rect 1346 1013 1364 1016
rect 1436 1013 1485 1016
rect 1546 1013 1556 1016
rect 1596 1013 1613 1016
rect 1700 1013 1725 1016
rect 1756 1013 1765 1016
rect 1796 1013 1805 1016
rect 1844 1013 1853 1016
rect 1914 1013 1933 1016
rect 988 1003 997 1006
rect 1034 1003 1043 1006
rect 1138 1003 1148 1006
rect 1498 1003 1508 1006
rect 1762 1005 1765 1013
rect 1818 1003 1829 1006
rect 1836 1003 1845 1006
rect 530 993 541 996
rect 1826 995 1829 1003
rect 1850 995 1853 1013
rect 1930 1005 1933 1013
rect 2002 1006 2005 1014
rect 2034 1006 2037 1014
rect 2282 1013 2292 1016
rect 1946 1003 1964 1006
rect 1978 1003 1988 1006
rect 2002 1003 2013 1006
rect 2034 1003 2044 1006
rect 2276 1003 2284 1006
rect 2474 1003 2484 1006
rect 2586 996 2589 1023
rect 2594 1003 2612 1006
rect 2500 993 2525 996
rect 2586 993 2604 996
rect 38 967 2706 973
rect 2242 936 2245 946
rect 130 933 140 936
rect 242 933 253 936
rect 594 933 604 936
rect 682 933 700 936
rect 778 933 787 936
rect 802 933 812 936
rect 836 933 845 936
rect 898 933 908 936
rect 1010 933 1018 936
rect 1580 933 1597 936
rect 108 923 125 926
rect 242 925 245 933
rect 314 926 317 933
rect 306 923 317 926
rect 346 923 354 926
rect 386 923 396 926
rect 466 923 474 926
rect 506 923 516 926
rect 538 923 548 926
rect 578 923 587 926
rect 666 913 669 933
rect 1010 926 1013 933
rect 772 923 789 926
rect 810 923 820 926
rect 876 923 892 926
rect 1002 923 1013 926
rect 1034 923 1043 926
rect 1098 923 1108 926
rect 1114 923 1132 926
rect 1170 923 1188 926
rect 1236 923 1261 926
rect 1322 923 1340 926
rect 1388 923 1413 926
rect 1474 923 1492 926
rect 1564 923 1573 926
rect 1594 925 1597 933
rect 2194 933 2252 936
rect 1626 923 1636 926
rect 1676 923 1685 926
rect 1786 923 1796 926
rect 1802 923 1820 926
rect 1850 923 1860 926
rect 1890 923 1900 926
rect 2194 923 2197 933
rect 2266 926 2269 945
rect 2282 943 2292 946
rect 2356 943 2365 946
rect 2276 933 2300 936
rect 2330 933 2340 936
rect 2354 933 2380 936
rect 2498 926 2501 935
rect 2260 923 2269 926
rect 2322 923 2332 926
rect 2490 923 2501 926
rect 1116 913 1125 916
rect 1170 915 1173 923
rect 1322 915 1325 923
rect 1474 915 1477 923
rect 1716 913 1725 916
rect 1506 903 1524 906
rect 1714 903 1732 906
rect 2514 903 2517 935
rect 2546 933 2556 936
rect 2572 933 2589 936
rect 2618 933 2628 936
rect 2530 923 2548 926
rect 2586 925 2589 933
rect 2626 923 2636 926
rect 14 867 2730 873
rect 1010 833 1018 836
rect 1042 833 1052 836
rect 1250 833 1276 836
rect 1290 833 1301 836
rect 1418 833 1436 836
rect 1522 833 1532 836
rect 1842 833 1868 836
rect 1930 833 1940 836
rect 2610 833 2628 836
rect 220 823 229 826
rect 258 816 261 825
rect 644 823 661 826
rect 124 813 133 816
rect 164 813 173 816
rect 186 813 212 816
rect 258 813 269 816
rect 276 813 285 816
rect 362 813 372 816
rect 442 813 451 816
rect 530 813 540 816
rect 578 813 595 816
rect 676 813 693 816
rect 708 813 724 816
rect 130 803 140 806
rect 266 805 269 813
rect 477 803 485 806
rect 690 795 693 813
rect 730 806 733 825
rect 834 813 852 816
rect 874 813 884 816
rect 906 813 916 816
rect 986 813 996 816
rect 730 803 748 806
rect 804 803 813 806
rect 820 803 837 806
rect 858 803 876 806
rect 946 803 956 806
rect 1010 783 1013 814
rect 1066 813 1084 816
rect 1090 813 1100 816
rect 1114 813 1125 816
rect 1146 813 1173 816
rect 1298 815 1301 833
rect 1658 816 1661 825
rect 1842 816 1845 833
rect 2186 816 2189 825
rect 2242 823 2268 826
rect 2292 823 2317 826
rect 2498 823 2508 826
rect 1484 813 1500 816
rect 1612 813 1621 816
rect 1658 813 1669 816
rect 1682 813 1692 816
rect 1738 813 1748 816
rect 1780 813 1789 816
rect 1826 813 1845 816
rect 1954 813 1972 816
rect 2002 813 2012 816
rect 2140 813 2157 816
rect 2186 813 2204 816
rect 2442 813 2452 816
rect 2484 813 2493 816
rect 1114 805 1117 813
rect 1146 805 1149 813
rect 1380 803 1397 806
rect 1476 803 1485 806
rect 1660 803 1668 806
rect 1708 803 1717 806
rect 1754 803 1772 806
rect 2322 803 2332 806
rect 2642 803 2652 806
rect 38 767 2706 773
rect 442 733 468 736
rect 506 733 531 736
rect 554 733 564 736
rect 578 733 588 736
rect 690 726 693 734
rect 764 733 781 736
rect 866 733 876 736
rect 907 726 910 744
rect 916 733 933 736
rect 956 733 973 736
rect 346 723 476 726
rect 477 723 517 726
rect 562 723 572 726
rect 660 723 693 726
rect 738 723 748 726
rect 770 723 780 726
rect 810 723 820 726
rect 842 723 852 726
rect 858 723 868 726
rect 900 723 910 726
rect 924 723 932 726
rect 1002 725 1005 736
rect 1068 733 1077 736
rect 1316 733 1325 736
rect 1332 733 1341 736
rect 1362 733 1372 736
rect 1690 733 1700 736
rect 1009 723 1018 726
rect 1092 723 1101 726
rect 1140 723 1165 726
rect 1356 723 1365 726
rect 1380 723 1397 726
rect 1516 723 1525 726
rect 1722 725 1725 756
rect 2346 743 2364 746
rect 1820 733 1837 736
rect 1866 733 1892 736
rect 2106 733 2148 736
rect 2162 733 2172 736
rect 2362 733 2372 736
rect 2378 733 2388 736
rect 2412 733 2429 736
rect 1834 723 1844 726
rect 2132 723 2149 726
rect 2156 723 2173 726
rect 2186 723 2196 726
rect 2210 723 2228 726
rect 2276 723 2293 726
rect 2380 723 2389 726
rect 2396 723 2405 726
rect 2420 723 2437 726
rect 2482 723 2492 726
rect 2580 723 2589 726
rect 2626 723 2636 726
rect 764 713 773 716
rect 1028 713 1037 716
rect 1364 713 1373 716
rect 1716 713 1725 716
rect 1932 713 1941 716
rect 2210 715 2213 723
rect 2586 716 2589 723
rect 2586 713 2597 716
rect 770 693 773 713
rect 1026 703 1043 706
rect 14 667 2730 673
rect 748 623 757 626
rect 1378 616 1381 636
rect 1642 633 1660 636
rect 2130 633 2141 636
rect 2226 633 2244 636
rect 2266 633 2276 636
rect 2124 623 2132 626
rect 212 613 237 616
rect 268 613 277 616
rect 314 605 317 616
rect 386 613 396 616
rect 468 613 477 616
rect 484 613 493 616
rect 514 606 517 614
rect 546 606 549 614
rect 620 613 645 616
rect 778 613 788 616
rect 948 613 973 616
rect 1004 613 1013 616
rect 1084 613 1093 616
rect 1276 613 1285 616
rect 1300 613 1309 616
rect 1316 613 1333 616
rect 1372 613 1381 616
rect 1388 613 1405 616
rect 1412 613 1429 616
rect 1548 613 1557 616
rect 388 603 397 606
rect 466 603 476 606
rect 500 603 517 606
rect 538 603 549 606
rect 1036 603 1045 606
rect 1098 603 1108 606
rect 1258 603 1268 606
rect 1292 603 1308 606
rect 1340 603 1357 606
rect 1370 603 1380 606
rect 1394 603 1404 606
rect 1554 605 1557 613
rect 1586 606 1589 614
rect 1604 613 1620 616
rect 1730 613 1740 616
rect 1930 613 1940 616
rect 1946 613 1964 616
rect 1994 613 2004 616
rect 2138 615 2141 633
rect 2228 623 2237 626
rect 2172 613 2181 616
rect 2324 613 2341 616
rect 2420 613 2429 616
rect 1586 603 1596 606
rect 1722 603 1732 606
rect 1780 603 1789 606
rect 1274 593 1284 596
rect 38 567 2706 573
rect 1626 536 1629 546
rect 1634 543 1652 546
rect 1666 536 1669 546
rect 2258 536 2261 546
rect 274 533 308 536
rect 378 526 381 535
rect 410 533 420 536
rect 714 533 724 536
rect 834 526 837 535
rect 946 526 949 535
rect 962 526 965 535
rect 1066 533 1076 536
rect 1082 533 1092 536
rect 1316 533 1325 536
rect 1332 533 1348 536
rect 1362 533 1380 536
rect 1620 533 1629 536
rect 1660 533 1669 536
rect 204 523 229 526
rect 260 523 301 526
rect 306 523 316 526
rect 346 523 381 526
rect 410 523 428 526
rect 476 523 501 526
rect 538 523 548 526
rect 604 523 629 526
rect 666 523 676 526
rect 690 523 708 526
rect 714 523 732 526
rect 772 523 797 526
rect 828 523 837 526
rect 884 523 901 526
rect 940 523 949 526
rect 956 523 965 526
rect 1356 523 1373 526
rect 1394 523 1404 526
rect 1522 523 1532 526
rect 1668 523 1677 526
rect 1684 523 1693 526
rect 1714 525 1717 536
rect 1748 533 1757 536
rect 1794 533 1804 536
rect 2258 533 2276 536
rect 1812 523 1829 526
rect 1842 523 1852 526
rect 1922 523 1932 526
rect 1986 523 1996 526
rect 2026 523 2036 526
rect 2284 523 2325 526
rect 2420 523 2429 526
rect 2564 523 2573 526
rect 2620 523 2637 526
rect 410 516 413 523
rect 396 513 413 516
rect 690 515 693 523
rect 1034 503 1037 515
rect 1764 513 1773 516
rect 1938 513 1965 516
rect 1714 503 1724 506
rect 1762 503 1780 506
rect 1946 503 1972 506
rect 14 467 2730 473
rect 2522 453 2573 456
rect 554 433 564 436
rect 1370 433 1396 436
rect 1650 433 1668 436
rect 1682 433 1700 436
rect 1786 433 1804 436
rect 2346 433 2365 436
rect 2346 426 2349 433
rect 572 423 581 426
rect 628 423 661 426
rect 850 416 853 425
rect 1068 423 1077 426
rect 1434 416 1437 426
rect 1452 423 1469 426
rect 1676 423 1684 426
rect 1788 423 1797 426
rect 1956 423 1965 426
rect 2332 423 2349 426
rect 268 413 293 416
rect 324 413 333 416
rect 378 413 388 416
rect 436 413 461 416
rect 578 413 605 416
rect 626 413 668 416
rect 682 413 692 416
rect 706 413 716 416
rect 756 413 765 416
rect 810 413 836 416
rect 850 413 868 416
rect 930 413 956 416
rect 1034 413 1052 416
rect 1130 413 1196 416
rect 1434 413 1444 416
rect 1450 413 1484 416
rect 498 403 516 406
rect 602 405 605 413
rect 1538 406 1541 414
rect 1732 413 1741 416
rect 1818 413 1844 416
rect 1924 413 1933 416
rect 2124 413 2149 416
rect 2228 413 2253 416
rect 2474 413 2516 416
rect 722 403 748 406
rect 754 403 772 406
rect 778 403 796 406
rect 874 403 892 406
rect 906 403 948 406
rect 972 403 988 406
rect 1002 403 1044 406
rect 1092 403 1108 406
rect 1234 403 1244 406
rect 1332 403 1341 406
rect 1356 403 1373 406
rect 1426 403 1436 406
rect 1538 403 1557 406
rect 1906 403 1916 406
rect 1922 403 1932 406
rect 2290 403 2308 406
rect 2386 403 2444 406
rect 730 393 740 396
rect 1226 393 1236 396
rect 38 367 2706 373
rect 426 336 429 345
rect 1306 343 1316 346
rect 1330 343 1340 346
rect 274 333 300 336
rect 354 326 357 335
rect 420 333 429 336
rect 436 333 453 336
rect 458 333 468 336
rect 682 333 700 336
rect 706 333 724 336
rect 754 333 772 336
rect 796 333 812 336
rect 890 333 900 336
rect 922 333 940 336
rect 986 333 996 336
rect 1018 333 1036 336
rect 1210 333 1228 336
rect 1252 333 1268 336
rect 1300 333 1317 336
rect 1324 333 1341 336
rect 1348 333 1357 336
rect 1362 326 1365 345
rect 2444 343 2453 346
rect 1378 333 1388 336
rect 1402 333 1412 336
rect 1426 333 1436 336
rect 1450 333 1460 336
rect 1610 326 1613 335
rect 2330 333 2340 336
rect 2370 333 2380 336
rect 2386 333 2428 336
rect 204 323 229 326
rect 260 323 301 326
rect 348 323 357 326
rect 364 323 404 326
rect 580 323 605 326
rect 642 323 652 326
rect 708 323 717 326
rect 748 323 765 326
rect 780 323 789 326
rect 1100 323 1125 326
rect 1186 323 1204 326
rect 1210 323 1221 326
rect 1276 323 1293 326
rect 1356 323 1365 326
rect 1386 323 1396 326
rect 1444 323 1461 326
rect 1468 323 1485 326
rect 1604 323 1613 326
rect 1658 323 1668 326
rect 1698 323 1708 326
rect 1810 323 1820 326
rect 2164 323 2189 326
rect 2220 323 2237 326
rect 2386 325 2389 333
rect 2586 326 2589 335
rect 2394 323 2420 326
rect 2570 323 2589 326
rect 500 313 509 316
rect 1186 315 1189 323
rect 1210 315 1213 323
rect 2234 316 2237 323
rect 1628 313 1637 316
rect 2234 313 2244 316
rect 2564 313 2573 316
rect 498 303 516 306
rect 1634 303 1644 306
rect 2458 303 2484 306
rect 14 267 2730 273
rect 546 233 564 236
rect 834 233 852 236
rect 2402 233 2421 236
rect 2490 233 2516 236
rect 2402 226 2405 233
rect 636 223 645 226
rect 860 223 885 226
rect 2236 223 2253 226
rect 2332 223 2349 226
rect 2396 223 2405 226
rect 268 213 293 216
rect 324 213 333 216
rect 340 213 356 216
rect 418 213 428 216
rect 442 213 460 216
rect 500 213 516 216
rect 578 213 613 216
rect 634 213 660 216
rect 674 213 692 216
rect 788 213 797 216
rect 866 213 899 216
rect 914 213 932 216
rect 1010 213 1020 216
rect 1068 213 1077 216
rect 1084 213 1100 216
rect 1130 213 1140 216
rect 1186 213 1196 216
rect 1202 213 1236 216
rect 1330 213 1372 216
rect 1386 213 1404 216
rect 1418 213 1436 216
rect 1548 213 1557 216
rect 1618 213 1628 216
rect 1634 213 1668 216
rect 1698 213 1708 216
rect 1762 213 1772 216
rect 1786 213 1797 216
rect 1994 213 2004 216
rect 2108 213 2133 216
rect 2164 213 2189 216
rect 2196 213 2220 216
rect 2372 213 2388 216
rect 2418 215 2421 233
rect 2500 223 2509 226
rect 2554 213 2565 216
rect 330 205 333 213
rect 610 205 613 213
rect 794 206 797 213
rect 698 203 716 206
rect 794 203 804 206
rect 954 203 972 206
rect 1026 203 1036 206
rect 1050 203 1060 206
rect 1074 205 1077 213
rect 1202 203 1228 206
rect 1242 203 1252 206
rect 1298 203 1308 206
rect 1410 203 1428 206
rect 1554 205 1557 213
rect 1650 203 1660 206
rect 1794 205 1797 213
rect 1946 203 1956 206
rect 2186 205 2189 213
rect 2242 203 2252 206
rect 2354 203 2364 206
rect 2562 205 2565 213
rect 1202 193 1205 203
rect 2338 193 2356 196
rect 38 167 2706 173
rect 476 123 501 126
rect 588 123 613 126
rect 788 123 813 126
rect 844 123 853 126
rect 892 123 917 126
rect 1084 123 1109 126
rect 1292 123 1317 126
rect 1588 123 1597 126
rect 1796 123 1805 126
rect 14 67 2730 73
rect 38 37 2706 57
rect 14 13 2730 33
<< metal2 >>
rect 14 13 34 2627
rect 38 37 58 2603
rect 1282 2563 1325 2566
rect 122 2553 157 2556
rect 74 2503 77 2536
rect 122 2533 125 2553
rect 146 2536 149 2546
rect 130 2533 149 2536
rect 122 2513 125 2526
rect 130 2503 133 2526
rect 74 2343 77 2416
rect 130 2413 133 2426
rect 122 2333 125 2356
rect 130 2316 133 2406
rect 122 2313 133 2316
rect 122 2213 125 2313
rect 74 2193 77 2206
rect 122 2156 125 2206
rect 130 2193 133 2226
rect 138 2213 141 2533
rect 154 2526 157 2553
rect 530 2553 573 2556
rect 162 2533 173 2536
rect 154 2523 165 2526
rect 146 2413 149 2426
rect 154 2413 157 2523
rect 170 2466 173 2533
rect 234 2526 237 2546
rect 178 2503 181 2526
rect 202 2513 205 2526
rect 226 2523 237 2526
rect 242 2516 245 2536
rect 266 2533 269 2546
rect 258 2523 269 2526
rect 274 2523 277 2536
rect 330 2523 341 2526
rect 354 2523 357 2546
rect 378 2516 381 2526
rect 242 2513 293 2516
rect 338 2513 381 2516
rect 170 2463 181 2466
rect 178 2386 181 2463
rect 194 2393 197 2416
rect 218 2413 221 2426
rect 266 2413 269 2506
rect 386 2496 389 2536
rect 378 2493 389 2496
rect 378 2436 381 2493
rect 378 2433 389 2436
rect 290 2413 293 2426
rect 178 2383 205 2386
rect 146 2333 149 2346
rect 194 2333 197 2356
rect 202 2333 205 2383
rect 218 2353 245 2356
rect 218 2336 221 2353
rect 210 2333 221 2336
rect 210 2306 213 2333
rect 218 2316 221 2326
rect 226 2323 229 2346
rect 234 2323 237 2336
rect 242 2323 245 2353
rect 266 2333 269 2406
rect 274 2333 277 2356
rect 290 2343 293 2356
rect 298 2333 301 2416
rect 330 2356 333 2416
rect 362 2376 365 2416
rect 386 2413 389 2433
rect 394 2423 397 2546
rect 402 2496 405 2526
rect 426 2513 429 2536
rect 458 2523 469 2526
rect 482 2523 485 2546
rect 506 2516 509 2526
rect 530 2523 533 2553
rect 466 2513 509 2516
rect 402 2493 413 2496
rect 410 2436 413 2493
rect 538 2436 541 2546
rect 546 2516 549 2536
rect 562 2523 565 2536
rect 570 2533 573 2553
rect 850 2553 893 2556
rect 578 2523 581 2536
rect 634 2523 645 2526
rect 658 2523 661 2546
rect 682 2516 685 2526
rect 690 2523 693 2536
rect 546 2513 597 2516
rect 642 2513 685 2516
rect 402 2433 413 2436
rect 514 2433 541 2436
rect 402 2413 405 2433
rect 394 2386 397 2406
rect 402 2393 405 2406
rect 418 2386 421 2406
rect 394 2383 421 2386
rect 362 2373 373 2376
rect 314 2353 333 2356
rect 266 2316 269 2326
rect 218 2313 269 2316
rect 210 2303 229 2306
rect 146 2156 149 2226
rect 178 2213 189 2216
rect 194 2213 197 2226
rect 226 2213 229 2303
rect 314 2236 317 2353
rect 362 2316 365 2356
rect 370 2323 373 2373
rect 482 2356 485 2406
rect 490 2403 493 2416
rect 498 2413 501 2426
rect 514 2413 517 2433
rect 522 2423 541 2426
rect 522 2413 525 2423
rect 530 2406 533 2416
rect 538 2413 541 2423
rect 562 2413 565 2426
rect 570 2406 573 2506
rect 698 2496 701 2546
rect 690 2493 701 2496
rect 690 2416 693 2493
rect 514 2383 517 2406
rect 530 2403 573 2406
rect 418 2343 445 2346
rect 474 2343 477 2356
rect 482 2353 493 2356
rect 378 2323 381 2336
rect 418 2333 421 2343
rect 426 2326 429 2336
rect 442 2333 445 2343
rect 490 2333 493 2353
rect 386 2323 453 2326
rect 386 2316 389 2323
rect 362 2313 389 2316
rect 314 2233 341 2236
rect 170 2203 205 2206
rect 122 2153 149 2156
rect 146 2143 149 2153
rect 250 2146 253 2216
rect 282 2213 285 2226
rect 274 2196 277 2206
rect 298 2203 301 2216
rect 306 2196 309 2216
rect 338 2213 341 2233
rect 274 2193 309 2196
rect 362 2166 365 2226
rect 394 2213 397 2226
rect 402 2213 413 2216
rect 450 2213 453 2323
rect 498 2296 501 2336
rect 570 2333 573 2403
rect 586 2393 589 2406
rect 602 2356 605 2416
rect 626 2403 629 2416
rect 586 2353 605 2356
rect 586 2333 589 2353
rect 634 2346 637 2416
rect 682 2413 693 2416
rect 642 2393 645 2406
rect 682 2393 685 2406
rect 698 2403 701 2426
rect 706 2413 709 2526
rect 730 2513 733 2536
rect 762 2523 773 2526
rect 786 2523 789 2546
rect 818 2543 845 2546
rect 818 2533 821 2543
rect 762 2506 765 2523
rect 810 2516 813 2526
rect 826 2523 829 2536
rect 842 2533 845 2543
rect 770 2513 813 2516
rect 842 2516 845 2526
rect 850 2523 853 2553
rect 858 2516 861 2546
rect 842 2513 861 2516
rect 866 2516 869 2536
rect 890 2533 893 2553
rect 890 2523 901 2526
rect 954 2523 965 2526
rect 978 2523 981 2556
rect 1002 2516 1005 2526
rect 866 2513 917 2516
rect 962 2513 1005 2516
rect 762 2503 789 2506
rect 762 2413 765 2426
rect 770 2406 773 2416
rect 754 2393 757 2406
rect 762 2403 773 2406
rect 778 2406 781 2416
rect 786 2413 789 2503
rect 898 2493 901 2506
rect 1010 2503 1013 2536
rect 794 2406 797 2416
rect 818 2413 821 2426
rect 858 2413 861 2466
rect 1018 2463 1021 2536
rect 1026 2513 1029 2526
rect 1090 2523 1093 2536
rect 1138 2533 1141 2556
rect 1106 2523 1117 2526
rect 1130 2516 1133 2526
rect 1042 2493 1045 2516
rect 1090 2513 1133 2516
rect 1138 2513 1141 2526
rect 778 2403 797 2406
rect 850 2393 853 2406
rect 634 2343 645 2346
rect 506 2306 509 2326
rect 530 2306 533 2326
rect 506 2303 533 2306
rect 490 2293 501 2296
rect 458 2213 461 2226
rect 386 2203 421 2206
rect 210 2143 253 2146
rect 338 2163 365 2166
rect 338 2143 341 2163
rect 98 2116 101 2136
rect 210 2133 221 2136
rect 90 2113 101 2116
rect 90 2036 93 2113
rect 90 2033 101 2036
rect 98 2013 101 2033
rect 114 1963 117 2126
rect 122 2103 125 2126
rect 226 2096 229 2136
rect 218 2093 229 2096
rect 218 2016 221 2093
rect 218 2013 229 2016
rect 218 1983 221 1996
rect 226 1986 229 2013
rect 242 1993 245 2126
rect 250 2113 253 2126
rect 346 2103 349 2136
rect 378 2133 381 2146
rect 386 2036 389 2126
rect 394 2123 397 2186
rect 482 2143 485 2206
rect 490 2203 493 2293
rect 538 2226 541 2326
rect 634 2313 637 2336
rect 642 2323 645 2343
rect 690 2343 709 2346
rect 650 2323 653 2336
rect 690 2333 693 2343
rect 706 2336 709 2343
rect 658 2313 661 2326
rect 698 2313 701 2336
rect 706 2333 717 2336
rect 778 2323 781 2356
rect 858 2353 861 2396
rect 882 2376 885 2426
rect 890 2413 893 2436
rect 882 2373 893 2376
rect 890 2343 893 2373
rect 786 2233 789 2336
rect 802 2323 805 2336
rect 898 2323 901 2336
rect 906 2333 909 2416
rect 930 2403 933 2446
rect 938 2356 941 2416
rect 946 2413 949 2436
rect 954 2413 957 2426
rect 994 2416 997 2426
rect 978 2413 997 2416
rect 938 2353 973 2356
rect 970 2323 973 2353
rect 978 2333 981 2413
rect 986 2396 989 2406
rect 994 2403 997 2413
rect 1002 2403 1013 2406
rect 1066 2403 1069 2456
rect 1146 2453 1149 2536
rect 1162 2526 1165 2536
rect 1170 2533 1173 2546
rect 1162 2523 1173 2526
rect 1162 2443 1165 2516
rect 1170 2506 1173 2523
rect 1170 2503 1197 2506
rect 1146 2423 1189 2426
rect 1002 2396 1005 2403
rect 1074 2396 1077 2406
rect 986 2393 1005 2396
rect 1058 2393 1077 2396
rect 1090 2386 1093 2416
rect 1146 2413 1149 2423
rect 1138 2386 1141 2406
rect 1090 2383 1141 2386
rect 1154 2386 1157 2416
rect 1162 2393 1165 2416
rect 1186 2413 1189 2423
rect 1194 2386 1197 2503
rect 1218 2453 1221 2536
rect 1226 2533 1229 2546
rect 1226 2506 1229 2526
rect 1234 2516 1237 2526
rect 1242 2523 1245 2536
rect 1282 2533 1285 2563
rect 1250 2516 1253 2526
rect 1234 2513 1253 2516
rect 1274 2506 1277 2526
rect 1226 2503 1277 2506
rect 1290 2503 1293 2536
rect 1306 2533 1309 2556
rect 1306 2516 1309 2526
rect 1314 2523 1317 2536
rect 1322 2533 1325 2563
rect 1330 2523 1333 2556
rect 1338 2516 1341 2546
rect 1370 2536 1373 2546
rect 1306 2513 1341 2516
rect 1346 2516 1349 2536
rect 1354 2533 1373 2536
rect 1354 2523 1365 2526
rect 1378 2523 1381 2536
rect 1434 2523 1445 2526
rect 1458 2523 1461 2546
rect 1346 2513 1397 2516
rect 1218 2413 1261 2416
rect 1202 2393 1205 2406
rect 1154 2383 1197 2386
rect 1218 2383 1221 2413
rect 1250 2396 1253 2406
rect 1258 2403 1261 2413
rect 1274 2396 1277 2406
rect 1250 2393 1277 2396
rect 1098 2343 1101 2383
rect 1250 2343 1253 2356
rect 994 2243 997 2336
rect 1098 2333 1109 2336
rect 1010 2313 1013 2326
rect 1146 2316 1149 2336
rect 1138 2313 1149 2316
rect 1138 2256 1141 2313
rect 1138 2253 1149 2256
rect 498 2223 541 2226
rect 498 2213 501 2223
rect 514 2203 517 2216
rect 530 2213 533 2223
rect 530 2193 533 2206
rect 538 2173 541 2216
rect 546 2203 549 2216
rect 634 2193 637 2216
rect 642 2183 645 2206
rect 626 2143 629 2176
rect 490 2113 493 2136
rect 634 2133 637 2146
rect 650 2143 653 2206
rect 658 2176 661 2216
rect 682 2206 685 2226
rect 722 2213 725 2226
rect 962 2216 965 2236
rect 682 2203 725 2206
rect 658 2173 701 2176
rect 226 1983 237 1986
rect 234 1943 237 1983
rect 130 1923 133 1936
rect 242 1933 245 1966
rect 250 1943 253 1956
rect 138 1913 141 1926
rect 146 1883 149 1926
rect 250 1913 253 1936
rect 266 1923 269 2016
rect 274 1943 277 1986
rect 282 1976 285 2016
rect 306 2003 309 2036
rect 386 2033 421 2036
rect 314 1983 317 2016
rect 322 2013 325 2026
rect 418 2016 421 2033
rect 410 2013 421 2016
rect 434 2013 437 2066
rect 450 2023 453 2036
rect 498 2023 501 2126
rect 530 2113 533 2126
rect 410 1993 413 2013
rect 418 1993 421 2006
rect 426 2003 437 2006
rect 490 2003 501 2006
rect 458 1993 509 1996
rect 282 1973 293 1976
rect 274 1923 277 1936
rect 290 1923 293 1973
rect 306 1933 309 1946
rect 410 1943 413 1986
rect 426 1943 429 1966
rect 314 1903 317 1926
rect 322 1913 325 1926
rect 418 1883 421 1936
rect 426 1913 429 1936
rect 442 1923 445 1956
rect 458 1943 461 1993
rect 506 1983 509 1993
rect 450 1903 453 1936
rect 474 1933 477 1946
rect 482 1943 485 1976
rect 482 1923 485 1936
rect 514 1923 517 2006
rect 522 1953 525 2046
rect 538 2033 541 2126
rect 658 2103 661 2146
rect 698 2133 701 2173
rect 738 2146 741 2216
rect 746 2183 749 2216
rect 834 2213 853 2216
rect 834 2193 837 2213
rect 842 2193 845 2206
rect 850 2163 853 2206
rect 866 2173 869 2216
rect 954 2213 965 2216
rect 954 2193 957 2213
rect 962 2193 965 2206
rect 970 2203 973 2216
rect 978 2186 981 2216
rect 986 2213 989 2226
rect 1082 2216 1085 2246
rect 1146 2233 1149 2253
rect 1162 2243 1165 2326
rect 1258 2313 1261 2336
rect 1282 2333 1285 2416
rect 1330 2393 1349 2396
rect 1330 2333 1333 2356
rect 1330 2316 1333 2326
rect 1338 2323 1341 2336
rect 1346 2323 1349 2393
rect 1354 2353 1357 2416
rect 1426 2413 1429 2436
rect 1362 2386 1365 2406
rect 1370 2393 1373 2406
rect 1418 2386 1421 2406
rect 1362 2383 1421 2386
rect 1434 2366 1437 2523
rect 1482 2516 1485 2526
rect 1490 2523 1493 2536
rect 1498 2533 1501 2556
rect 1442 2513 1485 2516
rect 1498 2436 1501 2526
rect 1530 2513 1533 2536
rect 1562 2523 1573 2526
rect 1586 2523 1589 2556
rect 1650 2553 1693 2556
rect 1618 2543 1645 2546
rect 1618 2533 1621 2543
rect 1562 2513 1565 2523
rect 1610 2516 1613 2526
rect 1626 2523 1629 2536
rect 1642 2533 1645 2543
rect 1570 2513 1613 2516
rect 1642 2516 1645 2526
rect 1650 2523 1653 2553
rect 1658 2516 1661 2546
rect 1642 2513 1661 2516
rect 1666 2513 1669 2536
rect 1690 2533 1693 2553
rect 1682 2446 1685 2526
rect 1666 2443 1685 2446
rect 1474 2433 1501 2436
rect 1442 2393 1445 2426
rect 1474 2413 1477 2433
rect 1482 2423 1501 2426
rect 1482 2413 1485 2423
rect 1434 2363 1445 2366
rect 1370 2316 1373 2326
rect 1378 2323 1381 2336
rect 1386 2333 1389 2346
rect 1402 2323 1405 2356
rect 1330 2313 1373 2316
rect 1074 2213 1085 2216
rect 1074 2193 1077 2213
rect 706 2136 709 2146
rect 738 2143 749 2146
rect 882 2143 885 2186
rect 978 2183 1037 2186
rect 1034 2143 1037 2183
rect 1082 2173 1085 2206
rect 706 2133 733 2136
rect 666 2123 701 2126
rect 714 2123 725 2126
rect 530 2003 533 2016
rect 538 1993 541 2016
rect 546 2013 549 2056
rect 642 2016 645 2036
rect 634 2013 645 2016
rect 634 1993 637 2013
rect 650 2003 653 2026
rect 650 1963 653 1996
rect 658 1993 661 2006
rect 666 2003 669 2123
rect 682 2086 685 2106
rect 682 2083 693 2086
rect 674 2003 677 2066
rect 690 2036 693 2083
rect 682 2033 693 2036
rect 682 1996 685 2033
rect 698 2013 709 2016
rect 714 2013 717 2123
rect 730 2116 733 2133
rect 726 2113 733 2116
rect 726 2026 729 2113
rect 746 2066 749 2143
rect 738 2063 749 2066
rect 738 2043 741 2063
rect 722 2023 729 2026
rect 738 2023 757 2026
rect 770 2023 773 2056
rect 778 2033 781 2136
rect 674 1993 693 1996
rect 474 1803 477 1856
rect 538 1853 541 1936
rect 586 1923 589 1956
rect 522 1793 525 1816
rect 122 1736 125 1776
rect 106 1733 125 1736
rect 186 1733 189 1746
rect 210 1733 213 1786
rect 66 1626 69 1646
rect 66 1623 85 1626
rect 82 1436 85 1623
rect 106 1516 109 1733
rect 130 1706 133 1726
rect 122 1703 133 1706
rect 122 1546 125 1703
rect 122 1543 133 1546
rect 130 1523 133 1543
rect 106 1513 117 1516
rect 74 1433 85 1436
rect 114 1436 117 1513
rect 138 1506 141 1726
rect 218 1723 221 1736
rect 234 1726 237 1736
rect 258 1733 269 1736
rect 274 1733 277 1756
rect 298 1733 301 1746
rect 314 1733 317 1766
rect 322 1733 333 1736
rect 226 1723 237 1726
rect 226 1716 229 1723
rect 202 1713 229 1716
rect 154 1636 157 1656
rect 154 1633 165 1636
rect 162 1576 165 1633
rect 258 1623 261 1726
rect 266 1706 269 1733
rect 282 1713 285 1726
rect 298 1706 301 1716
rect 266 1703 301 1706
rect 298 1633 301 1703
rect 274 1623 309 1626
rect 234 1583 237 1606
rect 154 1573 165 1576
rect 146 1533 149 1546
rect 134 1503 141 1506
rect 114 1433 125 1436
rect 74 1366 77 1433
rect 66 1363 77 1366
rect 66 1033 69 1363
rect 98 1353 101 1416
rect 66 896 69 1016
rect 74 1003 77 1336
rect 98 1313 101 1326
rect 82 983 85 1306
rect 90 1093 93 1296
rect 122 1213 125 1433
rect 134 1396 137 1503
rect 146 1403 149 1516
rect 154 1496 157 1573
rect 242 1566 245 1616
rect 242 1563 253 1566
rect 178 1533 181 1556
rect 162 1513 165 1526
rect 154 1493 161 1496
rect 158 1396 161 1493
rect 170 1403 173 1466
rect 186 1433 189 1526
rect 194 1523 197 1546
rect 242 1543 253 1546
rect 258 1536 261 1606
rect 282 1603 285 1616
rect 290 1593 293 1616
rect 306 1586 309 1606
rect 226 1523 229 1536
rect 234 1533 261 1536
rect 270 1583 309 1586
rect 270 1526 273 1583
rect 178 1423 205 1426
rect 202 1416 205 1423
rect 186 1403 189 1416
rect 194 1403 197 1416
rect 202 1413 213 1416
rect 210 1403 213 1413
rect 134 1393 141 1396
rect 130 1343 133 1366
rect 138 1346 141 1393
rect 154 1393 161 1396
rect 138 1343 149 1346
rect 154 1343 157 1393
rect 130 1313 133 1336
rect 138 1323 141 1336
rect 98 1103 101 1176
rect 106 1043 109 1186
rect 138 1143 141 1306
rect 146 1296 149 1343
rect 154 1333 165 1336
rect 210 1333 213 1366
rect 218 1353 221 1426
rect 234 1356 237 1436
rect 250 1423 253 1526
rect 266 1523 273 1526
rect 282 1523 285 1536
rect 298 1533 309 1536
rect 242 1413 253 1416
rect 266 1406 269 1523
rect 290 1503 293 1526
rect 306 1426 309 1516
rect 298 1423 309 1426
rect 250 1403 269 1406
rect 274 1403 277 1416
rect 266 1356 269 1396
rect 282 1373 285 1406
rect 290 1393 293 1416
rect 298 1396 301 1423
rect 306 1403 309 1416
rect 298 1393 309 1396
rect 234 1353 269 1356
rect 218 1333 221 1346
rect 154 1323 157 1333
rect 162 1313 165 1326
rect 210 1316 213 1326
rect 218 1323 229 1326
rect 234 1316 237 1353
rect 298 1346 301 1386
rect 306 1353 309 1393
rect 242 1323 245 1336
rect 210 1313 237 1316
rect 250 1313 253 1346
rect 298 1343 309 1346
rect 146 1293 157 1296
rect 146 1173 149 1206
rect 154 1183 157 1293
rect 258 1273 269 1276
rect 202 1233 221 1236
rect 202 1226 205 1233
rect 178 1223 205 1226
rect 178 1213 181 1223
rect 178 1173 181 1206
rect 186 1203 189 1216
rect 114 1133 141 1136
rect 186 1133 189 1156
rect 114 1116 117 1133
rect 114 1113 121 1116
rect 118 1056 121 1113
rect 130 1103 133 1126
rect 114 1053 121 1056
rect 114 1036 117 1053
rect 90 1033 117 1036
rect 90 953 93 1033
rect 130 946 133 986
rect 122 943 133 946
rect 74 923 77 936
rect 122 933 125 943
rect 66 893 77 896
rect 74 776 77 893
rect 98 793 101 806
rect 106 783 109 916
rect 122 913 125 926
rect 130 896 133 936
rect 122 893 133 896
rect 122 836 125 893
rect 138 843 141 1126
rect 154 1106 157 1126
rect 150 1103 157 1106
rect 150 1016 153 1103
rect 146 1013 153 1016
rect 146 923 149 1013
rect 154 923 157 996
rect 162 963 165 1076
rect 194 1073 197 1216
rect 210 1213 213 1226
rect 218 1213 221 1233
rect 226 1223 237 1226
rect 210 1146 213 1206
rect 250 1203 253 1236
rect 258 1213 261 1273
rect 266 1153 269 1206
rect 202 1123 205 1146
rect 210 1143 245 1146
rect 226 1066 229 1126
rect 234 1116 237 1136
rect 242 1123 245 1143
rect 250 1123 253 1136
rect 258 1133 261 1146
rect 266 1116 269 1126
rect 234 1113 269 1116
rect 178 1013 181 1046
rect 186 1016 189 1066
rect 226 1063 245 1066
rect 194 1023 221 1026
rect 226 1023 229 1046
rect 186 1013 197 1016
rect 170 996 173 1006
rect 194 1003 197 1013
rect 170 993 197 996
rect 186 936 189 956
rect 162 913 165 936
rect 170 933 189 936
rect 170 923 173 933
rect 122 833 133 836
rect 130 813 133 833
rect 170 813 173 856
rect 178 836 181 926
rect 194 923 197 993
rect 202 973 205 1006
rect 210 983 213 1016
rect 218 1006 221 1023
rect 218 1003 229 1006
rect 226 976 229 996
rect 210 973 229 976
rect 202 916 205 936
rect 194 913 205 916
rect 210 913 213 973
rect 234 936 237 1056
rect 242 1013 245 1063
rect 274 1053 277 1266
rect 282 1203 285 1216
rect 290 1213 293 1226
rect 298 1216 301 1336
rect 306 1323 309 1336
rect 298 1213 309 1216
rect 282 1143 285 1196
rect 298 1193 301 1206
rect 242 943 245 956
rect 178 833 189 836
rect 186 813 189 833
rect 74 773 85 776
rect 82 496 85 773
rect 130 723 133 806
rect 186 783 189 806
rect 194 743 197 913
rect 218 893 221 926
rect 226 923 229 936
rect 234 933 245 936
rect 250 933 253 976
rect 258 963 261 1036
rect 290 1023 293 1046
rect 298 1033 301 1166
rect 306 1133 309 1213
rect 314 1116 317 1676
rect 322 1656 325 1726
rect 338 1693 341 1726
rect 346 1683 349 1736
rect 354 1733 365 1736
rect 354 1656 357 1726
rect 362 1723 365 1733
rect 370 1713 373 1736
rect 378 1733 389 1736
rect 402 1733 405 1776
rect 418 1733 421 1786
rect 442 1753 485 1756
rect 378 1676 381 1726
rect 322 1653 357 1656
rect 370 1673 381 1676
rect 322 1513 325 1636
rect 322 1293 325 1336
rect 322 1173 325 1216
rect 330 1203 333 1546
rect 338 1513 341 1653
rect 346 1603 349 1646
rect 362 1593 365 1606
rect 346 1533 349 1566
rect 370 1526 373 1673
rect 378 1533 381 1666
rect 354 1523 373 1526
rect 354 1436 357 1523
rect 378 1506 381 1526
rect 346 1433 357 1436
rect 370 1503 381 1506
rect 338 1403 341 1416
rect 346 1413 349 1433
rect 354 1356 357 1426
rect 362 1403 365 1426
rect 370 1413 373 1503
rect 386 1443 389 1733
rect 394 1603 397 1656
rect 410 1613 413 1726
rect 426 1613 429 1726
rect 434 1673 437 1736
rect 442 1733 445 1753
rect 458 1733 461 1746
rect 442 1706 445 1726
rect 442 1703 453 1706
rect 450 1656 453 1703
rect 466 1686 469 1726
rect 474 1723 477 1736
rect 482 1733 485 1753
rect 466 1683 477 1686
rect 442 1653 453 1656
rect 402 1573 405 1606
rect 418 1583 421 1606
rect 434 1586 437 1626
rect 442 1613 445 1653
rect 434 1583 445 1586
rect 450 1583 453 1606
rect 394 1483 397 1536
rect 386 1413 389 1436
rect 402 1423 405 1526
rect 410 1503 413 1536
rect 418 1533 429 1536
rect 410 1416 413 1456
rect 418 1433 421 1526
rect 426 1453 429 1533
rect 378 1393 381 1406
rect 386 1403 397 1406
rect 346 1353 357 1356
rect 338 1313 341 1326
rect 346 1293 349 1353
rect 394 1333 397 1386
rect 402 1343 405 1416
rect 410 1413 417 1416
rect 414 1356 417 1413
rect 410 1353 417 1356
rect 410 1336 413 1353
rect 402 1333 413 1336
rect 402 1263 405 1333
rect 362 1226 365 1246
rect 362 1223 397 1226
rect 402 1223 405 1246
rect 346 1213 357 1216
rect 330 1143 333 1196
rect 338 1173 341 1206
rect 346 1166 349 1206
rect 338 1163 349 1166
rect 310 1113 317 1116
rect 310 1046 313 1113
rect 310 1043 317 1046
rect 274 993 277 1006
rect 282 986 285 1006
rect 258 933 261 956
rect 266 936 269 986
rect 274 983 285 986
rect 298 983 301 1006
rect 306 1003 309 1016
rect 274 943 277 983
rect 266 933 277 936
rect 282 933 285 976
rect 242 866 245 933
rect 250 873 253 926
rect 274 923 277 933
rect 290 923 293 946
rect 306 933 309 956
rect 298 923 309 926
rect 298 913 301 923
rect 226 813 229 826
rect 202 796 205 806
rect 234 803 237 866
rect 242 863 253 866
rect 242 813 245 836
rect 250 823 253 863
rect 258 823 261 856
rect 258 796 261 806
rect 202 793 261 796
rect 266 753 269 906
rect 274 793 277 886
rect 306 826 309 916
rect 282 823 309 826
rect 282 813 285 823
rect 290 813 309 816
rect 282 783 285 806
rect 298 803 309 806
rect 314 763 317 1043
rect 322 1023 325 1136
rect 338 1096 341 1163
rect 354 1133 357 1213
rect 362 1193 365 1206
rect 370 1203 373 1216
rect 378 1213 405 1216
rect 378 1136 381 1206
rect 386 1143 389 1156
rect 394 1143 397 1206
rect 402 1196 405 1213
rect 410 1203 413 1296
rect 426 1293 429 1446
rect 402 1193 413 1196
rect 330 1093 341 1096
rect 330 1053 333 1093
rect 330 1003 333 1046
rect 338 946 341 1086
rect 346 1066 349 1126
rect 362 1103 365 1126
rect 370 1086 373 1136
rect 378 1133 389 1136
rect 378 1113 381 1126
rect 366 1083 373 1086
rect 346 1063 357 1066
rect 330 943 341 946
rect 322 923 325 936
rect 330 916 333 943
rect 338 923 341 936
rect 346 933 349 1056
rect 354 1013 357 1063
rect 366 1026 369 1083
rect 362 1023 369 1026
rect 362 996 365 1023
rect 370 1003 373 1016
rect 378 1013 381 1106
rect 386 1013 389 1133
rect 362 993 381 996
rect 354 933 365 936
rect 378 933 381 993
rect 386 976 389 1006
rect 394 986 397 1096
rect 402 996 405 1186
rect 410 1133 413 1193
rect 418 1146 421 1256
rect 434 1243 437 1576
rect 442 1516 445 1583
rect 450 1533 453 1566
rect 442 1513 449 1516
rect 446 1456 449 1513
rect 446 1453 453 1456
rect 442 1413 445 1446
rect 442 1333 445 1406
rect 442 1313 445 1326
rect 450 1286 453 1453
rect 458 1323 461 1616
rect 466 1603 469 1616
rect 466 1523 469 1536
rect 474 1506 477 1683
rect 490 1583 493 1786
rect 506 1716 509 1736
rect 522 1733 525 1746
rect 502 1713 509 1716
rect 502 1646 505 1713
rect 502 1643 509 1646
rect 482 1523 485 1536
rect 490 1513 493 1566
rect 470 1503 477 1506
rect 470 1436 473 1503
rect 470 1433 477 1436
rect 466 1373 469 1406
rect 466 1333 469 1356
rect 474 1323 477 1433
rect 482 1403 485 1476
rect 490 1393 493 1416
rect 482 1333 485 1386
rect 498 1376 501 1626
rect 494 1373 501 1376
rect 466 1313 485 1316
rect 494 1296 497 1373
rect 442 1283 453 1286
rect 490 1293 497 1296
rect 426 1173 429 1206
rect 434 1156 437 1216
rect 442 1163 445 1283
rect 450 1213 453 1256
rect 450 1193 453 1206
rect 458 1186 461 1266
rect 466 1203 469 1216
rect 450 1183 461 1186
rect 434 1153 445 1156
rect 418 1143 437 1146
rect 418 1103 421 1126
rect 426 1093 429 1136
rect 434 1086 437 1143
rect 418 1083 437 1086
rect 410 1003 413 1076
rect 418 1013 421 1083
rect 434 1073 437 1083
rect 442 1066 445 1153
rect 434 1063 445 1066
rect 426 1013 429 1056
rect 434 1013 437 1063
rect 450 1053 453 1183
rect 402 993 413 996
rect 394 983 405 986
rect 386 973 397 976
rect 386 933 389 966
rect 394 926 397 973
rect 402 966 405 983
rect 410 976 413 993
rect 426 983 429 1006
rect 410 973 429 976
rect 402 963 421 966
rect 402 933 405 946
rect 418 933 421 963
rect 426 933 429 973
rect 434 943 437 1006
rect 442 1003 445 1026
rect 450 1013 453 1046
rect 322 913 333 916
rect 322 703 325 913
rect 338 903 341 916
rect 346 896 349 926
rect 362 896 365 926
rect 346 893 365 896
rect 370 896 373 926
rect 378 923 389 926
rect 394 923 405 926
rect 370 893 389 896
rect 346 866 349 893
rect 330 863 349 866
rect 330 813 333 863
rect 338 803 341 816
rect 346 803 349 816
rect 354 803 357 886
rect 362 816 365 893
rect 386 846 389 893
rect 394 853 397 906
rect 402 883 405 923
rect 410 846 413 926
rect 386 843 413 846
rect 362 813 373 816
rect 362 793 365 806
rect 370 773 373 813
rect 378 803 381 836
rect 386 803 389 843
rect 418 836 421 926
rect 394 833 421 836
rect 266 646 269 686
rect 258 643 269 646
rect 186 566 189 606
rect 234 593 237 616
rect 66 493 85 496
rect 178 563 189 566
rect 66 473 69 493
rect 178 333 181 563
rect 226 523 229 556
rect 258 466 261 643
rect 306 636 309 696
rect 274 633 309 636
rect 346 633 349 726
rect 394 656 397 833
rect 434 826 437 926
rect 442 913 445 936
rect 450 933 453 1006
rect 458 933 461 1166
rect 466 1093 469 1146
rect 474 1123 477 1246
rect 490 1236 493 1293
rect 506 1263 509 1643
rect 514 1413 517 1726
rect 530 1676 533 1726
rect 538 1723 541 1836
rect 546 1713 549 1886
rect 618 1883 621 1926
rect 658 1913 661 1936
rect 666 1933 685 1936
rect 690 1933 693 1956
rect 706 1946 709 2013
rect 714 1986 717 2006
rect 722 1993 725 2023
rect 738 2013 741 2023
rect 746 2006 749 2016
rect 730 2003 749 2006
rect 738 1986 741 1996
rect 714 1983 741 1986
rect 698 1943 709 1946
rect 698 1933 701 1943
rect 682 1926 685 1933
rect 666 1913 669 1926
rect 626 1833 653 1836
rect 554 1753 557 1816
rect 618 1803 621 1826
rect 626 1813 629 1833
rect 634 1813 637 1826
rect 650 1823 653 1833
rect 674 1823 677 1926
rect 682 1923 693 1926
rect 682 1913 693 1916
rect 690 1853 701 1856
rect 706 1853 709 1936
rect 754 1933 757 2023
rect 786 2006 789 2126
rect 794 2096 797 2126
rect 890 2113 893 2136
rect 794 2093 801 2096
rect 798 2016 801 2093
rect 810 2023 813 2046
rect 798 2013 845 2016
rect 850 2013 853 2046
rect 842 2006 845 2013
rect 866 2006 869 2056
rect 874 2023 901 2026
rect 874 2013 877 2023
rect 786 2003 821 2006
rect 842 2003 853 2006
rect 866 2003 877 2006
rect 882 2003 885 2016
rect 898 2013 901 2023
rect 906 2003 909 2036
rect 922 2013 925 2056
rect 930 2006 933 2136
rect 1042 2133 1045 2166
rect 1050 2133 1053 2146
rect 1090 2143 1093 2206
rect 938 2106 941 2126
rect 946 2113 949 2126
rect 938 2103 965 2106
rect 938 2013 941 2046
rect 962 2006 965 2103
rect 1082 2096 1085 2116
rect 1074 2093 1085 2096
rect 1074 2046 1077 2093
rect 1074 2043 1085 2046
rect 1090 2043 1093 2126
rect 1098 2123 1101 2216
rect 1106 2176 1109 2216
rect 1202 2203 1205 2226
rect 1210 2196 1213 2206
rect 1186 2193 1197 2196
rect 1202 2193 1213 2196
rect 1106 2173 1113 2176
rect 1110 2116 1113 2173
rect 1122 2133 1125 2156
rect 1194 2133 1197 2156
rect 1106 2113 1113 2116
rect 994 2033 1013 2036
rect 986 2006 989 2016
rect 994 2006 997 2033
rect 1002 2013 1005 2026
rect 1010 2013 1013 2033
rect 930 2003 949 2006
rect 962 2003 981 2006
rect 986 2003 997 2006
rect 826 1983 829 1996
rect 850 1966 853 1996
rect 834 1963 853 1966
rect 874 1936 877 2003
rect 906 1993 949 1996
rect 946 1983 949 1993
rect 978 1973 981 1996
rect 994 1963 997 2003
rect 1010 1993 1013 2006
rect 1026 1983 1029 1996
rect 1050 1973 1053 2016
rect 1066 2013 1069 2026
rect 1082 2023 1085 2043
rect 1106 2026 1109 2113
rect 1130 2086 1133 2126
rect 1154 2113 1157 2126
rect 1202 2113 1205 2193
rect 1250 2156 1253 2216
rect 1346 2203 1349 2246
rect 1370 2233 1421 2236
rect 1370 2203 1373 2233
rect 1394 2213 1405 2216
rect 1418 2213 1421 2233
rect 1338 2193 1349 2196
rect 1418 2193 1421 2206
rect 1426 2203 1429 2336
rect 1434 2333 1437 2356
rect 1442 2333 1445 2363
rect 1458 2333 1461 2346
rect 1490 2333 1493 2416
rect 1498 2413 1501 2423
rect 1522 2413 1525 2436
rect 1450 2203 1453 2296
rect 1538 2293 1541 2336
rect 1546 2313 1549 2326
rect 1562 2313 1565 2346
rect 1570 2323 1573 2426
rect 1626 2423 1629 2436
rect 1594 2403 1605 2406
rect 1578 2333 1597 2336
rect 1578 2236 1581 2333
rect 1586 2316 1589 2326
rect 1594 2323 1597 2333
rect 1602 2316 1605 2326
rect 1586 2313 1605 2316
rect 1626 2313 1629 2326
rect 1634 2296 1637 2336
rect 1666 2333 1669 2443
rect 1690 2433 1693 2526
rect 1754 2523 1765 2526
rect 1778 2523 1781 2546
rect 1706 2513 1717 2516
rect 1754 2503 1757 2523
rect 1802 2516 1805 2526
rect 1762 2513 1805 2516
rect 1674 2423 1717 2426
rect 1810 2423 1813 2526
rect 1842 2456 1845 2546
rect 1930 2543 1965 2546
rect 1930 2533 1933 2543
rect 1938 2533 1949 2536
rect 1890 2486 1893 2526
rect 1922 2513 1925 2526
rect 1930 2486 1933 2526
rect 1890 2483 1933 2486
rect 1826 2453 1845 2456
rect 1690 2403 1693 2416
rect 1706 2343 1709 2416
rect 1714 2413 1717 2423
rect 1570 2233 1581 2236
rect 1626 2293 1637 2296
rect 1458 2223 1477 2226
rect 1458 2193 1461 2223
rect 1466 2183 1469 2216
rect 1474 2213 1477 2223
rect 1506 2196 1509 2206
rect 1514 2203 1525 2206
rect 1530 2196 1533 2206
rect 1506 2193 1533 2196
rect 1538 2186 1541 2216
rect 1530 2183 1541 2186
rect 1546 2183 1549 2216
rect 1570 2213 1573 2233
rect 1626 2226 1629 2293
rect 1578 2213 1581 2226
rect 1626 2223 1637 2226
rect 1594 2213 1605 2216
rect 1626 2196 1629 2206
rect 1634 2203 1637 2223
rect 1642 2213 1645 2226
rect 1626 2193 1645 2196
rect 1250 2153 1261 2156
rect 1210 2133 1213 2146
rect 1130 2083 1145 2086
rect 1142 2026 1145 2083
rect 1226 2036 1229 2126
rect 1250 2046 1253 2126
rect 1258 2116 1261 2153
rect 1426 2153 1437 2156
rect 1266 2123 1269 2136
rect 1290 2133 1325 2136
rect 1282 2123 1301 2126
rect 1314 2116 1317 2126
rect 1370 2123 1373 2136
rect 1258 2113 1317 2116
rect 1378 2116 1381 2126
rect 1386 2123 1389 2136
rect 1418 2133 1421 2146
rect 1426 2126 1429 2153
rect 1394 2123 1429 2126
rect 1394 2116 1397 2123
rect 1378 2113 1397 2116
rect 1250 2043 1261 2046
rect 1154 2026 1157 2036
rect 1218 2033 1229 2036
rect 1106 2023 1125 2026
rect 1130 2003 1133 2026
rect 1142 2023 1149 2026
rect 1146 2006 1149 2023
rect 1154 2023 1189 2026
rect 1154 2013 1157 2023
rect 1138 1993 1141 2006
rect 1146 2003 1157 2006
rect 1178 2003 1181 2016
rect 1186 2013 1189 2023
rect 1218 2013 1221 2033
rect 1154 1983 1157 1996
rect 1034 1943 1085 1946
rect 778 1863 781 1936
rect 826 1893 829 1926
rect 642 1813 653 1816
rect 642 1806 645 1813
rect 626 1803 645 1806
rect 650 1793 653 1806
rect 658 1803 661 1816
rect 698 1803 701 1853
rect 530 1673 541 1676
rect 530 1593 533 1606
rect 530 1533 533 1566
rect 538 1526 541 1673
rect 546 1603 549 1626
rect 554 1613 557 1676
rect 562 1646 565 1726
rect 570 1716 573 1736
rect 578 1733 589 1736
rect 594 1733 597 1746
rect 626 1733 629 1756
rect 634 1733 637 1776
rect 730 1773 733 1846
rect 746 1773 749 1816
rect 650 1733 653 1746
rect 578 1723 589 1726
rect 594 1716 597 1726
rect 570 1713 597 1716
rect 610 1656 613 1726
rect 618 1666 621 1716
rect 626 1673 629 1726
rect 618 1663 629 1666
rect 610 1653 621 1656
rect 562 1643 613 1646
rect 546 1546 549 1586
rect 554 1573 557 1606
rect 546 1543 557 1546
rect 522 1523 541 1526
rect 522 1413 525 1523
rect 546 1503 549 1536
rect 554 1493 557 1543
rect 562 1523 565 1643
rect 594 1613 597 1636
rect 570 1576 573 1586
rect 586 1583 589 1606
rect 570 1573 589 1576
rect 594 1573 597 1606
rect 602 1603 605 1616
rect 610 1613 613 1643
rect 618 1576 621 1653
rect 602 1573 621 1576
rect 531 1423 549 1426
rect 514 1403 525 1406
rect 514 1323 517 1403
rect 522 1316 525 1336
rect 514 1313 525 1316
rect 490 1233 501 1236
rect 498 1216 501 1233
rect 482 1213 501 1216
rect 482 1203 485 1213
rect 482 1116 485 1196
rect 490 1173 493 1206
rect 490 1133 493 1146
rect 498 1136 501 1213
rect 506 1143 509 1216
rect 498 1133 509 1136
rect 514 1133 517 1313
rect 530 1266 533 1366
rect 538 1323 541 1423
rect 546 1343 549 1386
rect 554 1316 557 1416
rect 562 1393 565 1506
rect 570 1386 573 1536
rect 586 1533 589 1573
rect 602 1546 605 1573
rect 594 1543 605 1546
rect 578 1496 581 1526
rect 594 1506 597 1543
rect 602 1523 605 1536
rect 610 1533 613 1566
rect 626 1563 629 1663
rect 634 1603 637 1646
rect 626 1533 637 1536
rect 594 1503 601 1506
rect 578 1493 585 1496
rect 582 1436 585 1493
rect 598 1446 601 1503
rect 610 1493 613 1526
rect 642 1523 645 1616
rect 650 1603 653 1646
rect 658 1633 661 1726
rect 666 1693 669 1736
rect 674 1733 677 1766
rect 706 1753 725 1756
rect 658 1573 661 1616
rect 666 1603 669 1656
rect 674 1613 677 1646
rect 674 1593 677 1606
rect 682 1586 685 1726
rect 690 1716 693 1736
rect 706 1733 709 1753
rect 714 1733 717 1746
rect 698 1723 709 1726
rect 714 1716 717 1726
rect 690 1713 717 1716
rect 722 1683 725 1753
rect 762 1733 765 1756
rect 762 1716 765 1726
rect 730 1713 757 1716
rect 762 1713 781 1716
rect 666 1583 685 1586
rect 650 1516 653 1566
rect 658 1533 661 1546
rect 642 1513 653 1516
rect 598 1443 605 1446
rect 582 1433 589 1436
rect 586 1413 589 1433
rect 594 1413 597 1426
rect 602 1413 605 1443
rect 578 1403 597 1406
rect 562 1383 573 1386
rect 562 1363 565 1383
rect 562 1323 565 1356
rect 570 1333 573 1376
rect 578 1333 581 1356
rect 570 1316 573 1326
rect 554 1313 573 1316
rect 490 1123 501 1126
rect 474 1113 485 1116
rect 474 1086 477 1113
rect 466 1083 477 1086
rect 466 933 469 1083
rect 474 1003 477 1026
rect 482 1013 485 1106
rect 482 996 485 1006
rect 474 993 485 996
rect 450 916 453 926
rect 450 913 461 916
rect 442 826 445 836
rect 410 823 445 826
rect 410 813 413 823
rect 402 753 405 806
rect 410 776 413 796
rect 418 783 421 806
rect 426 803 429 816
rect 442 813 445 823
rect 410 773 421 776
rect 394 653 405 656
rect 274 613 277 633
rect 282 613 285 626
rect 306 616 309 633
rect 322 623 333 626
rect 354 623 389 626
rect 274 476 277 606
rect 290 593 293 606
rect 298 603 301 616
rect 306 613 317 616
rect 322 613 325 623
rect 306 596 309 606
rect 338 603 341 616
rect 306 593 349 596
rect 298 523 301 536
rect 322 533 325 556
rect 306 513 309 526
rect 330 503 333 526
rect 274 473 281 476
rect 258 463 269 466
rect 242 366 245 406
rect 266 386 269 463
rect 278 406 281 473
rect 338 426 341 593
rect 362 553 365 606
rect 346 533 357 536
rect 370 526 373 616
rect 386 533 389 616
rect 394 583 397 606
rect 402 553 405 653
rect 410 613 413 646
rect 410 533 413 606
rect 418 603 421 773
rect 434 763 437 806
rect 426 623 437 626
rect 346 513 349 526
rect 370 523 389 526
rect 394 503 397 516
rect 426 496 429 623
rect 434 596 437 616
rect 442 603 445 806
rect 450 803 453 913
rect 458 803 461 866
rect 466 833 469 926
rect 466 803 469 816
rect 474 786 477 993
rect 482 933 485 976
rect 490 943 493 1006
rect 498 1003 501 1096
rect 506 1053 509 1133
rect 522 1116 525 1266
rect 530 1263 549 1266
rect 530 1213 533 1226
rect 538 1213 541 1256
rect 546 1213 549 1263
rect 554 1213 557 1246
rect 530 1153 533 1206
rect 538 1146 541 1206
rect 546 1173 549 1205
rect 562 1203 565 1306
rect 586 1303 589 1396
rect 594 1333 597 1376
rect 570 1186 573 1226
rect 578 1196 581 1216
rect 594 1213 597 1326
rect 602 1296 605 1326
rect 610 1303 613 1476
rect 618 1363 621 1426
rect 626 1413 629 1436
rect 618 1323 621 1336
rect 626 1333 629 1356
rect 634 1316 637 1446
rect 642 1323 645 1513
rect 666 1486 669 1583
rect 674 1506 677 1536
rect 682 1523 685 1576
rect 690 1533 693 1666
rect 698 1533 701 1586
rect 698 1506 701 1526
rect 674 1503 701 1506
rect 706 1493 709 1606
rect 714 1563 717 1606
rect 722 1556 725 1576
rect 714 1553 725 1556
rect 714 1486 717 1553
rect 722 1523 725 1536
rect 730 1513 733 1713
rect 786 1706 789 1726
rect 778 1703 789 1706
rect 778 1646 781 1703
rect 794 1693 797 1806
rect 802 1796 805 1866
rect 810 1803 813 1826
rect 818 1813 821 1826
rect 826 1813 829 1876
rect 858 1843 861 1926
rect 866 1923 869 1936
rect 874 1933 885 1936
rect 890 1926 893 1936
rect 874 1836 877 1926
rect 882 1923 893 1926
rect 882 1893 885 1923
rect 898 1846 901 1936
rect 914 1913 917 1926
rect 946 1886 949 1936
rect 1034 1933 1037 1943
rect 1058 1926 1061 1936
rect 994 1903 997 1926
rect 938 1883 949 1886
rect 938 1863 941 1883
rect 898 1843 909 1846
rect 858 1833 877 1836
rect 834 1823 845 1826
rect 834 1813 845 1816
rect 834 1806 837 1813
rect 818 1803 837 1806
rect 802 1793 821 1796
rect 778 1643 789 1646
rect 754 1603 757 1636
rect 738 1496 741 1556
rect 666 1483 677 1486
rect 658 1413 661 1456
rect 650 1393 653 1406
rect 666 1403 669 1476
rect 674 1413 677 1483
rect 706 1483 717 1486
rect 734 1493 741 1496
rect 682 1356 685 1426
rect 650 1353 685 1356
rect 690 1353 693 1476
rect 698 1403 701 1416
rect 706 1413 709 1483
rect 734 1426 737 1493
rect 734 1423 741 1426
rect 714 1413 725 1416
rect 706 1403 717 1406
rect 618 1313 637 1316
rect 602 1293 613 1296
rect 602 1206 605 1276
rect 610 1223 613 1293
rect 586 1203 597 1206
rect 602 1203 613 1206
rect 578 1193 613 1196
rect 570 1183 581 1186
rect 518 1113 525 1116
rect 530 1143 549 1146
rect 518 1046 521 1113
rect 518 1043 525 1046
rect 522 1023 525 1043
rect 506 1013 517 1016
rect 522 993 525 1006
rect 530 1003 533 1143
rect 538 1006 541 1136
rect 546 1133 549 1143
rect 546 1013 549 1126
rect 554 1066 557 1156
rect 562 1133 565 1146
rect 578 1133 581 1183
rect 602 1146 605 1166
rect 610 1156 613 1193
rect 618 1163 621 1313
rect 626 1266 629 1306
rect 642 1273 645 1316
rect 650 1276 653 1353
rect 658 1333 661 1346
rect 658 1313 661 1326
rect 706 1306 709 1403
rect 730 1393 733 1406
rect 714 1343 717 1366
rect 738 1353 741 1423
rect 746 1353 749 1526
rect 754 1423 757 1566
rect 770 1546 773 1596
rect 786 1586 789 1643
rect 762 1543 773 1546
rect 778 1583 789 1586
rect 762 1433 765 1543
rect 770 1506 773 1526
rect 778 1523 781 1583
rect 802 1573 805 1616
rect 818 1596 821 1793
rect 842 1773 845 1806
rect 850 1793 853 1806
rect 858 1786 861 1833
rect 850 1783 861 1786
rect 834 1603 837 1616
rect 850 1613 853 1783
rect 866 1723 869 1746
rect 882 1633 885 1806
rect 906 1746 909 1843
rect 914 1773 917 1796
rect 930 1793 933 1816
rect 890 1743 909 1746
rect 890 1676 893 1743
rect 898 1733 909 1736
rect 898 1723 901 1733
rect 914 1726 917 1766
rect 910 1723 917 1726
rect 890 1673 901 1676
rect 890 1626 893 1646
rect 858 1623 893 1626
rect 858 1606 861 1623
rect 842 1603 861 1606
rect 818 1593 845 1596
rect 786 1563 821 1566
rect 786 1533 789 1563
rect 794 1523 797 1536
rect 802 1533 805 1556
rect 810 1506 813 1536
rect 818 1523 821 1563
rect 770 1503 805 1506
rect 810 1503 821 1506
rect 786 1403 789 1496
rect 802 1403 805 1503
rect 802 1363 805 1396
rect 714 1333 733 1336
rect 738 1333 741 1346
rect 746 1333 757 1336
rect 802 1333 805 1346
rect 690 1303 709 1306
rect 650 1273 661 1276
rect 626 1263 653 1266
rect 626 1215 629 1256
rect 626 1203 637 1206
rect 610 1153 621 1156
rect 594 1136 597 1146
rect 602 1143 613 1146
rect 594 1133 605 1136
rect 554 1063 565 1066
rect 554 1023 557 1056
rect 562 1043 565 1063
rect 570 1056 573 1126
rect 586 1093 589 1126
rect 602 1093 605 1133
rect 570 1053 581 1056
rect 570 1023 573 1036
rect 554 1013 573 1016
rect 578 1013 581 1053
rect 538 1003 549 1006
rect 554 1003 557 1013
rect 586 1006 589 1056
rect 570 1003 589 1006
rect 530 986 533 996
rect 498 983 533 986
rect 498 933 501 983
rect 506 933 509 946
rect 514 933 533 936
rect 538 933 541 976
rect 482 886 485 926
rect 490 913 493 926
rect 498 923 509 926
rect 482 883 493 886
rect 482 803 485 816
rect 466 783 477 786
rect 466 736 469 783
rect 466 733 477 736
rect 474 713 477 733
rect 450 613 453 666
rect 458 603 461 636
rect 466 596 469 606
rect 434 593 469 596
rect 466 553 469 593
rect 394 493 429 496
rect 290 413 293 426
rect 322 423 341 426
rect 346 423 381 426
rect 262 383 269 386
rect 274 403 281 406
rect 274 386 277 403
rect 322 386 325 423
rect 330 393 333 416
rect 346 413 349 423
rect 274 383 285 386
rect 322 383 333 386
rect 338 383 341 406
rect 354 403 357 416
rect 362 413 373 416
rect 378 413 381 423
rect 394 406 397 493
rect 450 456 453 536
rect 242 363 253 366
rect 226 323 229 356
rect 250 286 253 363
rect 262 296 265 383
rect 274 303 277 383
rect 298 323 301 346
rect 322 336 325 356
rect 306 323 309 336
rect 314 333 325 336
rect 330 333 333 383
rect 338 333 341 346
rect 370 336 373 406
rect 378 403 397 406
rect 410 453 453 456
rect 378 393 381 403
rect 410 393 413 453
rect 450 396 453 446
rect 474 416 477 616
rect 482 443 485 786
rect 490 633 493 883
rect 498 863 501 923
rect 514 916 517 933
rect 546 926 549 1003
rect 554 933 565 936
rect 570 933 573 1003
rect 578 993 589 996
rect 578 933 581 986
rect 506 913 517 916
rect 506 873 509 913
rect 514 816 517 896
rect 530 866 533 916
rect 522 863 533 866
rect 538 906 541 926
rect 546 923 557 926
rect 538 903 549 906
rect 522 823 525 863
rect 538 856 541 903
rect 554 896 557 923
rect 530 853 541 856
rect 546 893 557 896
rect 498 783 501 806
rect 506 803 509 816
rect 514 813 525 816
rect 530 813 533 853
rect 546 813 549 893
rect 562 856 565 926
rect 578 903 581 926
rect 554 853 565 856
rect 554 813 557 853
rect 522 803 525 813
rect 498 716 501 756
rect 506 733 509 746
rect 514 723 517 766
rect 522 723 525 736
rect 498 713 505 716
rect 502 646 505 713
rect 530 696 533 806
rect 546 783 549 806
rect 562 803 565 846
rect 570 796 573 836
rect 538 723 541 756
rect 546 713 549 736
rect 554 733 557 796
rect 562 793 573 796
rect 514 693 533 696
rect 554 693 557 726
rect 514 653 517 693
rect 562 686 565 793
rect 578 773 581 816
rect 526 683 565 686
rect 502 643 517 646
rect 490 613 501 616
rect 506 613 509 626
rect 490 423 493 606
rect 498 523 501 536
rect 458 403 461 416
rect 474 413 493 416
rect 498 403 501 506
rect 514 476 517 643
rect 526 626 529 683
rect 578 676 581 736
rect 586 683 589 993
rect 594 933 597 1026
rect 602 1013 605 1076
rect 594 796 597 916
rect 602 913 605 1006
rect 610 973 613 1143
rect 618 1133 621 1153
rect 634 1133 637 1146
rect 626 1103 629 1126
rect 618 1003 621 1036
rect 610 893 613 926
rect 618 903 621 986
rect 626 933 629 1096
rect 634 1023 637 1036
rect 634 983 637 1016
rect 642 1013 645 1246
rect 650 1126 653 1263
rect 658 1133 661 1273
rect 666 1176 669 1266
rect 674 1203 677 1296
rect 690 1236 693 1303
rect 714 1293 717 1326
rect 722 1286 725 1326
rect 730 1313 733 1333
rect 714 1283 725 1286
rect 690 1233 701 1236
rect 682 1203 685 1216
rect 690 1186 693 1216
rect 682 1183 693 1186
rect 666 1173 677 1176
rect 650 1123 661 1126
rect 642 943 645 1006
rect 650 986 653 1116
rect 658 1053 661 1123
rect 658 996 661 1036
rect 666 1003 669 1166
rect 674 1083 677 1173
rect 682 1076 685 1183
rect 690 1083 693 1176
rect 698 1143 701 1233
rect 706 1213 709 1256
rect 706 1196 709 1206
rect 714 1203 717 1283
rect 722 1223 741 1226
rect 722 1213 725 1223
rect 722 1196 725 1206
rect 706 1193 725 1196
rect 706 1133 709 1186
rect 698 1103 701 1126
rect 682 1073 693 1076
rect 658 993 669 996
rect 650 983 661 986
rect 610 813 613 856
rect 602 803 613 806
rect 618 803 621 826
rect 626 803 629 896
rect 594 793 605 796
rect 594 733 597 786
rect 594 703 597 726
rect 602 723 605 793
rect 618 723 621 756
rect 626 716 629 796
rect 634 773 637 926
rect 642 863 645 936
rect 658 933 661 983
rect 666 933 669 993
rect 674 983 677 1046
rect 682 933 685 1006
rect 650 853 653 926
rect 650 796 653 846
rect 658 823 661 916
rect 666 893 669 916
rect 674 903 677 926
rect 682 913 685 926
rect 690 923 693 1073
rect 714 1066 717 1176
rect 722 1113 725 1136
rect 730 1116 733 1216
rect 738 1173 741 1223
rect 730 1113 741 1116
rect 706 1063 733 1066
rect 698 973 701 1006
rect 706 976 709 1063
rect 714 1013 725 1016
rect 730 1013 733 1063
rect 722 983 725 1006
rect 706 973 725 976
rect 682 823 685 866
rect 650 793 661 796
rect 562 673 581 676
rect 522 623 529 626
rect 522 603 525 623
rect 538 613 541 626
rect 530 603 541 606
rect 538 583 541 596
rect 546 576 549 616
rect 554 603 557 636
rect 562 613 565 673
rect 586 666 589 676
rect 570 663 589 666
rect 602 663 605 716
rect 570 603 573 663
rect 610 643 613 716
rect 618 713 629 716
rect 634 713 637 756
rect 578 583 581 616
rect 538 573 549 576
rect 538 566 541 573
rect 594 566 597 636
rect 618 586 621 713
rect 626 693 629 706
rect 522 563 541 566
rect 586 563 597 566
rect 614 583 621 586
rect 522 483 525 563
rect 530 523 533 556
rect 538 533 541 563
rect 554 533 565 536
rect 510 473 517 476
rect 510 416 513 473
rect 538 446 541 526
rect 562 513 565 526
rect 578 513 581 536
rect 522 443 541 446
rect 510 413 517 416
rect 522 413 525 443
rect 538 423 541 436
rect 546 423 549 506
rect 602 496 605 536
rect 594 493 605 496
rect 554 433 557 486
rect 578 423 581 466
rect 546 413 581 416
rect 514 396 517 413
rect 530 403 541 406
rect 586 403 589 426
rect 450 393 461 396
rect 514 393 533 396
rect 322 316 325 326
rect 346 323 349 336
rect 370 333 381 336
rect 378 316 381 333
rect 322 313 373 316
rect 378 313 385 316
rect 262 293 269 296
rect 242 283 253 286
rect 242 143 245 283
rect 266 246 269 293
rect 266 243 277 246
rect 274 196 277 243
rect 290 203 293 216
rect 266 193 277 196
rect 266 163 269 193
rect 346 173 349 306
rect 370 243 373 313
rect 382 246 385 313
rect 394 273 397 356
rect 418 296 421 316
rect 410 293 421 296
rect 378 243 385 246
rect 354 213 365 216
rect 354 203 365 206
rect 370 196 373 216
rect 378 206 381 243
rect 386 213 389 226
rect 378 203 389 206
rect 394 196 397 216
rect 402 206 405 236
rect 410 223 413 293
rect 442 236 445 326
rect 450 313 453 336
rect 458 333 461 393
rect 466 326 469 346
rect 458 323 469 326
rect 474 343 509 346
rect 474 323 477 343
rect 482 323 485 336
rect 442 233 461 236
rect 442 223 453 226
rect 410 213 421 216
rect 426 213 445 216
rect 426 206 429 213
rect 402 203 429 206
rect 370 193 397 196
rect 442 193 445 206
rect 394 183 397 193
rect 450 163 453 206
rect 458 193 461 233
rect 450 133 453 146
rect 490 143 493 326
rect 506 323 509 343
rect 498 303 501 316
rect 506 303 509 316
rect 522 313 525 336
rect 530 323 533 393
rect 538 296 541 326
rect 538 293 549 296
rect 546 233 549 293
rect 554 286 557 396
rect 594 343 597 493
rect 614 486 617 583
rect 626 533 629 666
rect 642 656 645 746
rect 650 733 653 786
rect 658 663 661 793
rect 666 773 669 806
rect 690 763 693 856
rect 698 836 701 966
rect 706 893 709 926
rect 714 873 717 936
rect 722 903 725 973
rect 730 943 733 1006
rect 698 833 717 836
rect 730 833 733 936
rect 738 923 741 1113
rect 698 816 701 826
rect 714 823 717 833
rect 698 813 709 816
rect 698 756 701 806
rect 706 776 709 813
rect 714 793 717 806
rect 722 803 733 806
rect 706 773 713 776
rect 666 753 701 756
rect 642 653 661 656
rect 634 566 637 626
rect 642 603 645 616
rect 634 563 645 566
rect 642 546 645 563
rect 642 543 649 546
rect 626 493 629 526
rect 646 486 649 543
rect 658 523 661 653
rect 666 596 669 753
rect 674 613 677 726
rect 690 723 701 726
rect 682 603 685 626
rect 690 613 693 723
rect 710 716 713 773
rect 722 733 725 803
rect 738 783 741 916
rect 746 793 749 1333
rect 754 1306 757 1326
rect 754 1303 773 1306
rect 754 1223 757 1256
rect 762 1213 765 1246
rect 754 1096 757 1206
rect 762 1183 765 1206
rect 762 1103 765 1116
rect 770 1113 773 1303
rect 778 1206 781 1326
rect 802 1313 805 1326
rect 786 1213 789 1256
rect 778 1203 789 1206
rect 754 1093 773 1096
rect 754 1006 757 1076
rect 762 1013 765 1026
rect 770 1013 773 1093
rect 754 1003 765 1006
rect 778 1003 781 1196
rect 786 1153 789 1203
rect 794 1166 797 1306
rect 810 1276 813 1376
rect 818 1293 821 1503
rect 826 1493 829 1556
rect 842 1533 845 1593
rect 866 1573 869 1606
rect 874 1603 885 1606
rect 874 1586 877 1603
rect 874 1583 881 1586
rect 842 1436 845 1516
rect 838 1433 845 1436
rect 838 1386 841 1433
rect 826 1306 829 1386
rect 838 1383 845 1386
rect 834 1353 837 1366
rect 842 1353 845 1383
rect 850 1346 853 1426
rect 834 1343 853 1346
rect 834 1333 837 1343
rect 858 1336 861 1456
rect 866 1446 869 1536
rect 878 1476 881 1583
rect 898 1566 901 1673
rect 910 1646 913 1723
rect 922 1713 925 1736
rect 930 1703 933 1726
rect 938 1713 941 1736
rect 946 1696 949 1836
rect 1034 1833 1037 1926
rect 1042 1886 1045 1926
rect 1050 1923 1061 1926
rect 1050 1903 1053 1923
rect 1066 1893 1069 1936
rect 1082 1913 1085 1943
rect 1042 1883 1049 1886
rect 978 1823 1029 1826
rect 962 1763 965 1816
rect 978 1803 981 1823
rect 986 1786 989 1816
rect 1002 1793 1005 1806
rect 986 1783 1005 1786
rect 962 1733 965 1746
rect 954 1703 957 1716
rect 946 1693 953 1696
rect 906 1643 913 1646
rect 906 1576 909 1643
rect 922 1603 925 1636
rect 950 1626 953 1693
rect 950 1623 957 1626
rect 906 1573 925 1576
rect 898 1563 909 1566
rect 890 1523 893 1536
rect 906 1486 909 1563
rect 874 1473 881 1476
rect 894 1483 909 1486
rect 874 1453 877 1473
rect 866 1443 885 1446
rect 850 1333 861 1336
rect 826 1303 833 1306
rect 810 1273 821 1276
rect 802 1213 805 1226
rect 810 1203 813 1246
rect 794 1163 813 1166
rect 786 1033 789 1146
rect 794 1133 797 1146
rect 802 1123 805 1156
rect 802 1066 805 1116
rect 810 1073 813 1163
rect 802 1063 813 1066
rect 802 1013 805 1036
rect 754 933 757 976
rect 762 953 765 1003
rect 794 993 797 1006
rect 810 973 813 1063
rect 778 936 781 946
rect 762 933 781 936
rect 786 943 813 946
rect 818 943 821 1273
rect 830 1226 833 1303
rect 842 1253 845 1326
rect 858 1273 861 1326
rect 866 1303 869 1436
rect 874 1403 877 1416
rect 882 1403 885 1443
rect 894 1396 897 1483
rect 906 1413 909 1426
rect 890 1393 897 1396
rect 874 1333 877 1366
rect 890 1333 893 1393
rect 914 1336 917 1566
rect 922 1486 925 1573
rect 930 1506 933 1526
rect 938 1523 941 1556
rect 946 1533 949 1606
rect 930 1503 941 1506
rect 922 1483 929 1486
rect 926 1366 929 1483
rect 906 1333 917 1336
rect 922 1363 929 1366
rect 874 1236 877 1326
rect 850 1233 877 1236
rect 830 1223 845 1226
rect 826 1156 829 1216
rect 842 1163 845 1223
rect 850 1203 853 1233
rect 866 1213 869 1226
rect 874 1206 877 1233
rect 882 1213 885 1256
rect 890 1213 893 1316
rect 898 1303 901 1326
rect 906 1226 909 1333
rect 914 1293 917 1326
rect 922 1263 925 1363
rect 930 1323 933 1336
rect 930 1256 933 1296
rect 898 1223 909 1226
rect 922 1253 933 1256
rect 858 1203 869 1206
rect 874 1203 893 1206
rect 826 1153 853 1156
rect 826 1113 829 1136
rect 826 996 829 1016
rect 834 1003 837 1146
rect 842 1103 845 1146
rect 850 1096 853 1153
rect 866 1123 869 1203
rect 874 1133 877 1146
rect 890 1133 893 1146
rect 898 1116 901 1223
rect 922 1216 925 1253
rect 906 1156 909 1216
rect 914 1213 925 1216
rect 914 1193 917 1213
rect 922 1166 925 1206
rect 930 1203 933 1246
rect 938 1223 941 1503
rect 954 1333 957 1623
rect 962 1453 965 1716
rect 970 1706 973 1736
rect 970 1703 981 1706
rect 986 1703 989 1736
rect 994 1716 997 1726
rect 1002 1723 1005 1783
rect 1010 1763 1013 1806
rect 1034 1793 1037 1806
rect 1046 1786 1049 1883
rect 1042 1783 1049 1786
rect 994 1713 1021 1716
rect 970 1613 973 1696
rect 978 1656 981 1703
rect 1026 1693 1029 1736
rect 1034 1713 1037 1736
rect 1042 1733 1045 1783
rect 1058 1773 1061 1816
rect 1074 1806 1077 1826
rect 1082 1816 1085 1856
rect 1122 1846 1125 1936
rect 1130 1916 1133 1976
rect 1234 1973 1237 2006
rect 1258 1983 1261 2043
rect 1282 2013 1285 2026
rect 1322 1993 1325 2016
rect 1338 2006 1341 2026
rect 1346 2023 1373 2026
rect 1346 2013 1349 2023
rect 1330 2003 1341 2006
rect 1138 1933 1141 1946
rect 1146 1923 1149 1936
rect 1154 1933 1165 1936
rect 1154 1916 1157 1926
rect 1130 1913 1157 1916
rect 1170 1906 1173 1936
rect 1178 1913 1181 1926
rect 1170 1903 1197 1906
rect 1122 1843 1149 1846
rect 1122 1826 1125 1836
rect 1090 1823 1125 1826
rect 1082 1813 1093 1816
rect 1066 1803 1085 1806
rect 1090 1803 1093 1813
rect 1082 1796 1085 1803
rect 1098 1796 1101 1806
rect 1106 1803 1109 1816
rect 1082 1793 1101 1796
rect 1058 1733 1061 1756
rect 1074 1733 1077 1746
rect 978 1653 1005 1656
rect 986 1566 989 1653
rect 978 1563 989 1566
rect 994 1553 997 1616
rect 1002 1613 1005 1653
rect 1018 1603 1021 1636
rect 1042 1603 1045 1726
rect 1058 1703 1061 1726
rect 1066 1723 1077 1726
rect 1058 1636 1061 1656
rect 1054 1633 1061 1636
rect 1054 1576 1057 1633
rect 1066 1576 1069 1616
rect 1082 1586 1085 1786
rect 1090 1733 1101 1736
rect 1090 1643 1093 1726
rect 1106 1673 1109 1776
rect 1114 1723 1117 1823
rect 1146 1816 1149 1843
rect 1154 1823 1157 1836
rect 1122 1803 1125 1816
rect 1130 1756 1133 1806
rect 1138 1786 1141 1816
rect 1146 1813 1157 1816
rect 1154 1803 1157 1813
rect 1162 1803 1165 1826
rect 1186 1823 1189 1836
rect 1138 1783 1165 1786
rect 1154 1756 1157 1776
rect 1130 1753 1157 1756
rect 1130 1723 1133 1753
rect 1146 1733 1149 1746
rect 1154 1733 1157 1753
rect 1162 1743 1165 1783
rect 1170 1736 1173 1816
rect 1178 1813 1189 1816
rect 1178 1803 1181 1813
rect 1186 1793 1189 1806
rect 1194 1796 1197 1903
rect 1202 1863 1205 1936
rect 1250 1913 1253 1926
rect 1282 1923 1285 1946
rect 1322 1906 1325 1926
rect 1314 1903 1325 1906
rect 1330 1903 1333 2003
rect 1346 1996 1349 2006
rect 1338 1993 1349 1996
rect 1338 1933 1341 1993
rect 1354 1926 1357 2016
rect 1370 2003 1373 2016
rect 1378 2013 1381 2106
rect 1434 2046 1437 2146
rect 1434 2043 1441 2046
rect 1314 1846 1317 1903
rect 1338 1893 1341 1926
rect 1346 1846 1349 1926
rect 1354 1923 1365 1926
rect 1314 1843 1325 1846
rect 1218 1833 1229 1836
rect 1226 1826 1229 1833
rect 1202 1823 1221 1826
rect 1226 1823 1261 1826
rect 1202 1803 1205 1823
rect 1218 1816 1221 1823
rect 1218 1813 1229 1816
rect 1242 1813 1261 1816
rect 1282 1813 1285 1836
rect 1226 1796 1229 1806
rect 1194 1793 1229 1796
rect 1162 1733 1173 1736
rect 1178 1733 1181 1756
rect 1202 1753 1213 1756
rect 1234 1753 1237 1806
rect 1146 1713 1149 1726
rect 1082 1583 1093 1586
rect 1054 1573 1061 1576
rect 1066 1573 1085 1576
rect 970 1533 981 1536
rect 978 1496 981 1516
rect 970 1493 981 1496
rect 994 1473 997 1536
rect 946 1316 949 1326
rect 962 1316 965 1336
rect 946 1313 965 1316
rect 970 1313 973 1326
rect 978 1276 981 1396
rect 1002 1363 1005 1406
rect 1018 1386 1021 1546
rect 1042 1523 1045 1536
rect 1058 1516 1061 1573
rect 1090 1556 1093 1583
rect 1082 1553 1093 1556
rect 1066 1523 1077 1526
rect 1058 1513 1069 1516
rect 1034 1403 1037 1476
rect 1018 1383 1029 1386
rect 1002 1333 1005 1346
rect 1018 1326 1021 1336
rect 1026 1333 1029 1383
rect 986 1303 989 1316
rect 954 1273 981 1276
rect 938 1183 941 1216
rect 946 1173 949 1246
rect 922 1163 933 1166
rect 954 1163 957 1273
rect 962 1203 965 1216
rect 906 1153 925 1156
rect 914 1123 917 1136
rect 922 1133 925 1153
rect 846 1093 853 1096
rect 866 1113 901 1116
rect 922 1113 925 1126
rect 846 1036 849 1093
rect 842 1033 849 1036
rect 826 993 837 996
rect 754 893 757 916
rect 762 913 765 933
rect 770 866 773 926
rect 786 923 789 943
rect 794 933 805 936
rect 778 903 781 916
rect 754 863 773 866
rect 754 853 757 863
rect 706 713 713 716
rect 706 626 709 713
rect 706 623 717 626
rect 690 603 701 606
rect 666 593 701 596
rect 666 533 669 546
rect 614 483 621 486
rect 602 323 605 386
rect 610 366 613 446
rect 618 376 621 483
rect 642 483 649 486
rect 642 436 645 483
rect 666 443 669 526
rect 626 413 629 436
rect 642 433 649 436
rect 626 383 629 406
rect 618 373 629 376
rect 610 363 621 366
rect 554 283 589 286
rect 514 223 549 226
rect 514 213 517 223
rect 530 213 557 216
rect 570 213 573 226
rect 554 206 557 213
rect 578 206 581 216
rect 506 173 509 206
rect 522 166 525 206
rect 530 203 541 206
rect 554 203 581 206
rect 498 163 525 166
rect 498 123 501 163
rect 530 123 533 146
rect 538 133 541 203
rect 578 193 581 203
rect 562 133 565 146
rect 586 143 589 283
rect 618 216 621 363
rect 626 263 629 373
rect 634 323 637 426
rect 646 366 649 433
rect 658 423 661 436
rect 658 393 661 406
rect 674 386 677 426
rect 682 413 685 526
rect 690 493 693 536
rect 698 533 701 593
rect 706 526 709 616
rect 714 613 717 623
rect 714 593 717 606
rect 722 583 725 626
rect 714 536 717 556
rect 714 533 725 536
rect 706 523 717 526
rect 714 446 717 516
rect 722 503 725 533
rect 658 383 677 386
rect 682 383 685 406
rect 646 363 653 366
rect 642 333 645 356
rect 642 223 645 326
rect 650 293 653 363
rect 658 313 661 383
rect 690 343 693 446
rect 714 443 725 446
rect 730 443 733 736
rect 738 733 741 746
rect 738 683 741 726
rect 754 723 757 816
rect 770 803 773 856
rect 778 776 781 836
rect 786 803 789 896
rect 794 853 797 926
rect 802 913 805 926
rect 810 816 813 943
rect 818 886 821 936
rect 826 893 829 976
rect 834 966 837 993
rect 842 966 845 1033
rect 850 1003 853 1016
rect 858 1013 861 1036
rect 850 973 853 996
rect 858 993 861 1006
rect 858 966 861 986
rect 866 973 869 1113
rect 874 1023 885 1026
rect 834 963 853 966
rect 858 963 869 966
rect 842 933 845 946
rect 850 933 853 963
rect 834 896 837 916
rect 842 913 845 926
rect 858 896 861 926
rect 834 893 861 896
rect 866 893 869 963
rect 818 883 853 886
rect 794 803 797 816
rect 810 813 829 816
rect 834 813 837 836
rect 810 803 813 813
rect 834 796 837 806
rect 842 803 845 826
rect 850 803 853 883
rect 858 796 861 806
rect 810 776 813 796
rect 834 793 861 796
rect 762 773 781 776
rect 786 773 837 776
rect 762 663 765 773
rect 770 723 773 746
rect 778 733 781 766
rect 786 733 789 773
rect 802 743 805 766
rect 810 733 821 736
rect 762 633 765 646
rect 754 623 765 626
rect 770 623 773 696
rect 802 693 805 726
rect 778 683 789 686
rect 762 616 765 623
rect 778 616 781 683
rect 738 603 749 606
rect 738 573 741 603
rect 754 563 757 616
rect 762 613 781 616
rect 770 603 781 606
rect 746 513 749 536
rect 786 533 789 666
rect 810 643 813 726
rect 818 693 821 733
rect 826 713 829 736
rect 834 723 837 773
rect 850 736 853 766
rect 842 733 853 736
rect 842 683 845 726
rect 850 643 853 733
rect 794 603 797 626
rect 802 563 805 616
rect 810 553 813 606
rect 826 603 829 636
rect 850 613 853 626
rect 858 576 861 726
rect 866 693 869 886
rect 874 833 877 1023
rect 882 946 885 1016
rect 890 1013 893 1076
rect 898 1013 901 1036
rect 914 1016 917 1026
rect 906 1013 917 1016
rect 890 1003 901 1006
rect 882 943 893 946
rect 882 906 885 936
rect 890 933 893 943
rect 898 933 901 956
rect 906 943 909 1006
rect 914 936 917 1013
rect 922 1003 925 1016
rect 930 1013 933 1163
rect 962 1156 965 1196
rect 970 1176 973 1216
rect 978 1183 981 1266
rect 986 1213 989 1226
rect 994 1203 997 1326
rect 1002 1263 1005 1326
rect 1018 1323 1029 1326
rect 1050 1323 1053 1346
rect 1058 1333 1061 1506
rect 1066 1333 1069 1513
rect 1082 1426 1085 1553
rect 1098 1546 1101 1616
rect 1090 1543 1101 1546
rect 1106 1613 1117 1616
rect 1090 1503 1093 1543
rect 1106 1536 1109 1613
rect 1122 1603 1125 1686
rect 1162 1663 1165 1733
rect 1178 1713 1181 1726
rect 1130 1623 1157 1626
rect 1130 1613 1133 1623
rect 1138 1556 1141 1616
rect 1146 1613 1157 1616
rect 1154 1573 1157 1606
rect 1162 1603 1165 1616
rect 1170 1613 1181 1616
rect 1098 1533 1109 1536
rect 1114 1553 1141 1556
rect 1098 1513 1101 1533
rect 1106 1516 1109 1526
rect 1114 1523 1117 1553
rect 1122 1533 1133 1536
rect 1106 1513 1133 1516
rect 1146 1496 1149 1536
rect 1138 1493 1149 1496
rect 1074 1423 1085 1426
rect 1074 1386 1077 1423
rect 1082 1393 1085 1416
rect 1114 1413 1117 1486
rect 1138 1473 1141 1493
rect 1170 1486 1173 1613
rect 1178 1583 1181 1606
rect 1186 1573 1189 1746
rect 1194 1743 1245 1746
rect 1194 1733 1197 1743
rect 1242 1733 1245 1743
rect 1194 1683 1197 1726
rect 1202 1723 1213 1726
rect 1194 1596 1197 1676
rect 1202 1613 1205 1723
rect 1218 1706 1221 1726
rect 1218 1703 1229 1706
rect 1226 1646 1229 1703
rect 1250 1683 1253 1806
rect 1258 1763 1261 1806
rect 1266 1796 1269 1806
rect 1282 1803 1293 1806
rect 1298 1796 1301 1806
rect 1266 1793 1301 1796
rect 1306 1773 1309 1816
rect 1314 1743 1317 1806
rect 1322 1773 1325 1843
rect 1330 1843 1349 1846
rect 1330 1803 1333 1843
rect 1338 1813 1341 1836
rect 1354 1826 1357 1846
rect 1346 1823 1357 1826
rect 1338 1736 1341 1766
rect 1274 1733 1285 1736
rect 1298 1733 1341 1736
rect 1258 1706 1261 1726
rect 1266 1713 1269 1726
rect 1282 1706 1285 1716
rect 1258 1703 1285 1706
rect 1218 1643 1229 1646
rect 1218 1626 1221 1643
rect 1218 1623 1285 1626
rect 1290 1616 1293 1726
rect 1298 1696 1301 1716
rect 1314 1713 1317 1726
rect 1298 1693 1317 1696
rect 1218 1603 1221 1616
rect 1234 1613 1293 1616
rect 1298 1606 1301 1666
rect 1314 1623 1317 1693
rect 1322 1613 1325 1726
rect 1346 1713 1349 1726
rect 1354 1703 1357 1806
rect 1362 1786 1365 1923
rect 1370 1913 1373 1936
rect 1378 1933 1381 2006
rect 1410 1973 1413 2006
rect 1438 1996 1441 2043
rect 1434 1993 1441 1996
rect 1418 1933 1421 1946
rect 1434 1926 1437 1993
rect 1450 1933 1453 2016
rect 1458 1966 1461 2166
rect 1466 2133 1469 2146
rect 1514 2133 1517 2156
rect 1514 2116 1517 2126
rect 1522 2123 1525 2136
rect 1530 2123 1533 2183
rect 1562 2143 1573 2146
rect 1554 2116 1557 2126
rect 1514 2113 1557 2116
rect 1570 2036 1573 2136
rect 1586 2123 1589 2156
rect 1594 2133 1597 2146
rect 1602 2123 1605 2156
rect 1642 2136 1645 2193
rect 1650 2153 1653 2326
rect 1666 2313 1669 2326
rect 1698 2303 1701 2326
rect 1658 2216 1661 2226
rect 1658 2213 1693 2216
rect 1682 2156 1685 2206
rect 1690 2203 1693 2213
rect 1706 2163 1709 2336
rect 1714 2323 1717 2336
rect 1730 2293 1733 2326
rect 1738 2313 1741 2416
rect 1722 2213 1725 2236
rect 1754 2223 1757 2326
rect 1786 2313 1789 2326
rect 1818 2303 1821 2316
rect 1786 2223 1789 2236
rect 1730 2176 1733 2216
rect 1730 2173 1741 2176
rect 1674 2153 1685 2156
rect 1618 2133 1637 2136
rect 1642 2133 1669 2136
rect 1610 2103 1613 2126
rect 1618 2066 1621 2133
rect 1626 2123 1637 2126
rect 1642 2103 1645 2126
rect 1666 2103 1669 2133
rect 1618 2063 1645 2066
rect 1586 2053 1629 2056
rect 1490 1993 1493 2016
rect 1498 2013 1501 2036
rect 1570 2033 1581 2036
rect 1522 2006 1525 2026
rect 1506 2003 1525 2006
rect 1458 1963 1469 1966
rect 1426 1916 1429 1926
rect 1434 1923 1445 1926
rect 1378 1893 1381 1916
rect 1418 1903 1421 1916
rect 1426 1913 1453 1916
rect 1466 1906 1469 1963
rect 1538 1956 1541 2026
rect 1546 2023 1573 2026
rect 1546 2013 1549 2023
rect 1578 2016 1581 2033
rect 1554 2013 1581 2016
rect 1546 1963 1549 2006
rect 1554 1956 1557 2013
rect 1586 2003 1589 2053
rect 1626 2013 1629 2053
rect 1642 2006 1645 2063
rect 1602 1973 1605 2006
rect 1634 2003 1645 2006
rect 1674 2003 1677 2153
rect 1722 2133 1725 2146
rect 1698 2123 1709 2126
rect 1738 2123 1741 2173
rect 1826 2166 1829 2453
rect 1874 2413 1877 2436
rect 1906 2413 1909 2426
rect 1914 2413 1917 2436
rect 1930 2413 1933 2436
rect 1914 2393 1917 2406
rect 1938 2343 1941 2533
rect 1946 2503 1949 2526
rect 1962 2523 1965 2543
rect 2162 2543 2181 2546
rect 1946 2393 1949 2416
rect 1962 2413 1965 2426
rect 1970 2406 1973 2536
rect 1986 2513 1989 2526
rect 1994 2423 1997 2526
rect 2018 2523 2061 2526
rect 2018 2513 2021 2523
rect 2050 2503 2053 2516
rect 2066 2513 2069 2536
rect 2138 2523 2141 2536
rect 2162 2523 2165 2543
rect 2074 2513 2093 2516
rect 2034 2423 2037 2436
rect 1954 2403 1973 2406
rect 1874 2203 1877 2216
rect 1770 2163 1829 2166
rect 1770 2133 1773 2163
rect 1810 2146 1813 2163
rect 1802 2143 1813 2146
rect 1898 2146 1901 2336
rect 1906 2213 1909 2226
rect 1914 2223 1949 2226
rect 1914 2203 1917 2223
rect 1922 2203 1925 2216
rect 1930 2213 1941 2216
rect 1946 2213 1949 2223
rect 1930 2146 1933 2206
rect 1954 2166 1957 2403
rect 1978 2226 1981 2416
rect 2018 2343 2037 2346
rect 2002 2313 2005 2326
rect 2018 2323 2021 2343
rect 2026 2323 2029 2336
rect 2034 2333 2037 2343
rect 2058 2326 2061 2336
rect 2042 2323 2061 2326
rect 2066 2256 2069 2326
rect 2074 2323 2077 2513
rect 2170 2493 2173 2536
rect 2178 2533 2181 2543
rect 2210 2533 2213 2546
rect 2178 2513 2181 2526
rect 2194 2486 2197 2526
rect 2234 2486 2237 2526
rect 2290 2513 2293 2526
rect 2194 2483 2237 2486
rect 2306 2426 2309 2546
rect 2378 2533 2397 2536
rect 2434 2533 2437 2546
rect 2098 2323 2141 2326
rect 2098 2313 2101 2323
rect 2122 2313 2133 2316
rect 2066 2253 2093 2256
rect 1962 2213 1965 2226
rect 1898 2143 1933 2146
rect 1938 2163 1957 2166
rect 1746 2103 1749 2116
rect 1802 2046 1805 2143
rect 1818 2086 1821 2126
rect 1850 2113 1853 2126
rect 1858 2086 1861 2126
rect 1874 2116 1877 2136
rect 1898 2133 1901 2143
rect 1890 2123 1901 2126
rect 1906 2116 1909 2126
rect 1874 2113 1909 2116
rect 1818 2083 1861 2086
rect 1914 2046 1917 2143
rect 1938 2136 1941 2163
rect 1930 2133 1941 2136
rect 1922 2113 1925 2126
rect 1946 2113 1949 2126
rect 1970 2113 1973 2226
rect 1978 2223 1997 2226
rect 2034 2213 2037 2226
rect 2090 2213 2093 2253
rect 2146 2213 2149 2326
rect 2154 2313 2157 2336
rect 2186 2313 2189 2406
rect 2202 2403 2205 2416
rect 2234 2403 2237 2426
rect 2306 2423 2325 2426
rect 2290 2356 2293 2406
rect 2298 2373 2301 2416
rect 2306 2413 2317 2416
rect 2322 2406 2325 2423
rect 2330 2413 2333 2526
rect 2378 2516 2381 2533
rect 2374 2513 2381 2516
rect 2374 2436 2377 2513
rect 2374 2433 2381 2436
rect 2362 2413 2365 2426
rect 2378 2413 2381 2433
rect 2386 2413 2389 2526
rect 2418 2513 2421 2526
rect 2458 2513 2461 2526
rect 2402 2413 2405 2506
rect 2514 2503 2517 2526
rect 2426 2423 2429 2456
rect 2466 2453 2477 2456
rect 2458 2423 2469 2426
rect 2290 2353 2297 2356
rect 2266 2343 2285 2346
rect 2234 2236 2237 2336
rect 2266 2323 2269 2343
rect 2230 2233 2237 2236
rect 1802 2043 1829 2046
rect 1914 2043 1941 2046
rect 1682 2013 1685 2026
rect 1826 2003 1829 2043
rect 1874 2013 1877 2036
rect 1906 2013 1909 2026
rect 1914 2013 1917 2036
rect 1930 2013 1933 2036
rect 1914 2003 1925 2006
rect 1530 1953 1541 1956
rect 1546 1953 1557 1956
rect 1498 1943 1509 1946
rect 1498 1926 1501 1943
rect 1434 1903 1469 1906
rect 1490 1923 1501 1926
rect 1506 1923 1517 1926
rect 1386 1813 1389 1826
rect 1370 1803 1381 1806
rect 1362 1783 1373 1786
rect 1362 1696 1365 1776
rect 1370 1743 1373 1783
rect 1378 1733 1381 1803
rect 1394 1793 1397 1816
rect 1418 1806 1421 1816
rect 1402 1793 1405 1806
rect 1410 1763 1413 1806
rect 1418 1803 1429 1806
rect 1434 1803 1437 1903
rect 1418 1743 1421 1796
rect 1426 1793 1429 1803
rect 1442 1776 1445 1866
rect 1490 1846 1493 1923
rect 1434 1773 1445 1776
rect 1354 1693 1365 1696
rect 1330 1606 1333 1666
rect 1346 1623 1349 1646
rect 1402 1643 1405 1716
rect 1418 1626 1421 1726
rect 1370 1623 1421 1626
rect 1226 1596 1229 1606
rect 1194 1593 1229 1596
rect 1250 1583 1253 1606
rect 1258 1573 1261 1606
rect 1282 1566 1285 1606
rect 1290 1603 1301 1606
rect 1146 1483 1173 1486
rect 1146 1403 1149 1483
rect 1154 1423 1181 1426
rect 1154 1413 1157 1423
rect 1186 1416 1189 1566
rect 1282 1563 1293 1566
rect 1194 1523 1197 1546
rect 1226 1513 1229 1526
rect 1250 1513 1253 1536
rect 1258 1533 1277 1536
rect 1282 1533 1285 1546
rect 1290 1533 1293 1563
rect 1314 1533 1317 1606
rect 1322 1603 1333 1606
rect 1346 1586 1349 1616
rect 1370 1603 1373 1623
rect 1330 1583 1349 1586
rect 1330 1533 1333 1583
rect 1274 1526 1277 1533
rect 1162 1413 1189 1416
rect 1178 1393 1181 1406
rect 1074 1383 1085 1386
rect 1002 1213 1005 1246
rect 1010 1206 1013 1316
rect 1018 1273 1021 1316
rect 1026 1266 1029 1323
rect 1002 1203 1013 1206
rect 1018 1263 1029 1266
rect 970 1173 997 1176
rect 962 1153 973 1156
rect 962 1133 965 1146
rect 970 1136 973 1153
rect 970 1133 981 1136
rect 978 1123 981 1133
rect 930 986 933 1006
rect 938 993 941 1036
rect 946 1003 949 1046
rect 962 986 965 1006
rect 906 933 917 936
rect 890 923 901 926
rect 906 916 909 933
rect 898 913 909 916
rect 882 903 893 906
rect 874 813 877 826
rect 882 806 885 896
rect 890 853 893 903
rect 890 816 893 836
rect 898 823 901 913
rect 914 866 917 926
rect 922 883 925 986
rect 930 983 965 986
rect 970 983 973 1116
rect 978 1036 981 1056
rect 986 1043 989 1136
rect 994 1036 997 1173
rect 1002 1123 1005 1203
rect 1018 1196 1021 1263
rect 1034 1213 1045 1216
rect 1050 1213 1053 1246
rect 1042 1206 1045 1213
rect 1026 1203 1037 1206
rect 1042 1203 1053 1206
rect 1018 1193 1045 1196
rect 1050 1193 1053 1203
rect 1010 1093 1013 1126
rect 1034 1123 1037 1146
rect 1042 1103 1045 1193
rect 1050 1123 1053 1156
rect 1058 1113 1061 1326
rect 1066 1313 1069 1326
rect 1074 1256 1077 1326
rect 1082 1293 1085 1383
rect 1226 1353 1229 1496
rect 1258 1476 1261 1526
rect 1266 1503 1269 1526
rect 1274 1523 1285 1526
rect 1282 1476 1285 1516
rect 1258 1473 1285 1476
rect 1290 1446 1293 1466
rect 1290 1443 1297 1446
rect 1274 1393 1277 1416
rect 1294 1376 1297 1443
rect 1306 1413 1309 1426
rect 1314 1413 1317 1456
rect 1322 1426 1325 1526
rect 1330 1523 1341 1526
rect 1330 1453 1333 1523
rect 1346 1516 1349 1583
rect 1354 1533 1357 1546
rect 1362 1533 1365 1596
rect 1378 1523 1381 1616
rect 1394 1593 1397 1606
rect 1402 1563 1405 1606
rect 1346 1513 1381 1516
rect 1394 1493 1397 1536
rect 1418 1523 1421 1546
rect 1426 1503 1429 1736
rect 1434 1686 1437 1773
rect 1450 1736 1453 1846
rect 1490 1843 1501 1846
rect 1498 1823 1501 1843
rect 1506 1816 1509 1923
rect 1530 1903 1533 1953
rect 1538 1923 1541 1946
rect 1546 1916 1549 1953
rect 1538 1913 1549 1916
rect 1554 1943 1565 1946
rect 1538 1856 1541 1913
rect 1538 1853 1549 1856
rect 1458 1813 1493 1816
rect 1498 1813 1509 1816
rect 1522 1833 1541 1836
rect 1458 1743 1461 1806
rect 1466 1793 1477 1796
rect 1482 1736 1485 1806
rect 1498 1803 1501 1813
rect 1514 1793 1517 1806
rect 1522 1803 1525 1833
rect 1450 1733 1461 1736
rect 1482 1733 1525 1736
rect 1530 1733 1533 1826
rect 1546 1823 1549 1853
rect 1554 1816 1557 1943
rect 1570 1916 1573 1936
rect 1566 1913 1573 1916
rect 1566 1846 1569 1913
rect 1578 1856 1581 1926
rect 1594 1923 1597 1966
rect 1634 1953 1637 2003
rect 1610 1943 1637 1946
rect 1610 1933 1613 1943
rect 1618 1933 1629 1936
rect 1682 1933 1685 1976
rect 1602 1903 1605 1926
rect 1666 1886 1669 1926
rect 1706 1886 1709 1926
rect 1762 1923 1765 1936
rect 1666 1883 1709 1886
rect 1578 1853 1597 1856
rect 1566 1843 1573 1846
rect 1546 1813 1557 1816
rect 1562 1756 1565 1826
rect 1570 1803 1573 1843
rect 1586 1823 1589 1846
rect 1578 1766 1581 1816
rect 1546 1753 1565 1756
rect 1570 1763 1581 1766
rect 1546 1733 1549 1753
rect 1570 1746 1573 1763
rect 1594 1756 1597 1853
rect 1618 1833 1645 1836
rect 1618 1813 1621 1833
rect 1634 1816 1637 1826
rect 1626 1813 1637 1816
rect 1634 1796 1637 1806
rect 1642 1803 1645 1826
rect 1650 1813 1653 1826
rect 1698 1823 1717 1826
rect 1554 1743 1573 1746
rect 1442 1693 1445 1726
rect 1498 1713 1501 1726
rect 1434 1683 1445 1686
rect 1442 1576 1445 1683
rect 1506 1626 1509 1726
rect 1530 1723 1549 1726
rect 1522 1703 1525 1716
rect 1506 1623 1533 1626
rect 1466 1593 1469 1616
rect 1438 1573 1445 1576
rect 1438 1506 1441 1573
rect 1438 1503 1445 1506
rect 1442 1483 1445 1503
rect 1322 1423 1373 1426
rect 1322 1403 1325 1423
rect 1346 1393 1349 1406
rect 1354 1403 1357 1416
rect 1442 1403 1445 1476
rect 1466 1413 1469 1546
rect 1474 1523 1477 1586
rect 1522 1563 1525 1616
rect 1530 1613 1533 1623
rect 1546 1616 1549 1723
rect 1554 1716 1557 1743
rect 1578 1733 1581 1756
rect 1586 1753 1597 1756
rect 1562 1723 1581 1726
rect 1554 1713 1565 1716
rect 1554 1623 1557 1646
rect 1546 1613 1557 1616
rect 1530 1573 1533 1606
rect 1554 1566 1557 1606
rect 1562 1573 1565 1713
rect 1578 1693 1581 1716
rect 1586 1683 1589 1753
rect 1618 1733 1621 1796
rect 1634 1793 1661 1796
rect 1674 1793 1677 1806
rect 1626 1733 1629 1746
rect 1634 1733 1645 1736
rect 1594 1723 1613 1726
rect 1594 1706 1597 1723
rect 1594 1703 1601 1706
rect 1586 1623 1589 1646
rect 1598 1636 1601 1703
rect 1610 1643 1613 1716
rect 1634 1663 1637 1733
rect 1594 1633 1601 1636
rect 1546 1563 1557 1566
rect 1490 1426 1493 1536
rect 1506 1513 1509 1536
rect 1514 1533 1533 1536
rect 1538 1533 1541 1546
rect 1546 1533 1549 1563
rect 1586 1556 1589 1606
rect 1594 1603 1597 1633
rect 1642 1623 1645 1726
rect 1554 1553 1589 1556
rect 1530 1526 1533 1533
rect 1554 1526 1557 1553
rect 1602 1546 1605 1616
rect 1650 1613 1653 1726
rect 1658 1606 1661 1793
rect 1666 1733 1669 1746
rect 1682 1736 1685 1816
rect 1698 1813 1701 1823
rect 1698 1783 1701 1806
rect 1714 1803 1717 1823
rect 1722 1823 1749 1826
rect 1722 1813 1725 1823
rect 1730 1746 1733 1816
rect 1754 1803 1757 1826
rect 1770 1756 1773 1976
rect 1938 1946 1941 2043
rect 1946 2003 1949 2016
rect 1962 2013 1965 2026
rect 1978 2013 1981 2046
rect 1994 2023 1997 2116
rect 2002 2113 2005 2126
rect 2034 2076 2037 2166
rect 2066 2163 2069 2206
rect 2162 2163 2165 2206
rect 2210 2203 2213 2216
rect 2230 2176 2233 2233
rect 2230 2173 2237 2176
rect 2082 2123 2085 2146
rect 2114 2113 2117 2126
rect 2122 2116 2125 2136
rect 2130 2123 2133 2146
rect 2138 2133 2141 2156
rect 2234 2153 2237 2173
rect 2242 2136 2245 2226
rect 2250 2203 2253 2236
rect 2258 2203 2261 2216
rect 2266 2213 2269 2246
rect 2274 2206 2277 2336
rect 2282 2333 2285 2343
rect 2282 2313 2285 2326
rect 2294 2306 2297 2353
rect 2306 2323 2309 2406
rect 2314 2373 2317 2406
rect 2322 2403 2333 2406
rect 2330 2333 2333 2403
rect 2338 2393 2341 2406
rect 2386 2383 2389 2406
rect 2410 2403 2413 2416
rect 2474 2413 2477 2453
rect 2482 2403 2485 2426
rect 2490 2423 2509 2426
rect 2490 2366 2493 2423
rect 2450 2363 2493 2366
rect 2290 2303 2297 2306
rect 2290 2236 2293 2303
rect 2314 2286 2317 2326
rect 2354 2286 2357 2326
rect 2410 2313 2413 2326
rect 2442 2313 2445 2336
rect 2450 2323 2453 2363
rect 2530 2316 2533 2396
rect 2554 2393 2557 2406
rect 2562 2376 2565 2546
rect 2570 2423 2589 2426
rect 2570 2383 2573 2423
rect 2578 2396 2581 2416
rect 2586 2403 2589 2423
rect 2594 2413 2597 2426
rect 2602 2413 2605 2526
rect 2642 2423 2645 2526
rect 2594 2396 2597 2406
rect 2578 2393 2597 2396
rect 2562 2373 2589 2376
rect 2538 2343 2557 2346
rect 2538 2323 2541 2343
rect 2314 2283 2357 2286
rect 2282 2213 2285 2236
rect 2290 2233 2309 2236
rect 2298 2213 2301 2226
rect 2306 2206 2309 2233
rect 2314 2213 2317 2246
rect 2322 2213 2333 2216
rect 2154 2133 2165 2136
rect 2242 2133 2253 2136
rect 2138 2123 2149 2126
rect 2154 2116 2157 2126
rect 2122 2113 2157 2116
rect 2010 2073 2037 2076
rect 1938 1943 1957 1946
rect 1962 1923 1965 2006
rect 2010 1976 2013 2073
rect 2034 2023 2037 2036
rect 2090 2013 2093 2036
rect 2106 2023 2109 2046
rect 2162 2026 2165 2133
rect 2170 2113 2173 2126
rect 2186 2103 2189 2126
rect 2234 2123 2245 2126
rect 2250 2123 2253 2133
rect 2202 2046 2205 2116
rect 2242 2113 2245 2123
rect 2266 2096 2269 2206
rect 2274 2203 2293 2206
rect 2306 2203 2325 2206
rect 2290 2166 2293 2203
rect 2282 2163 2293 2166
rect 1994 1973 2013 1976
rect 1794 1813 1797 1826
rect 1850 1783 1853 1816
rect 1770 1753 1805 1756
rect 1682 1733 1693 1736
rect 1666 1643 1669 1716
rect 1674 1693 1677 1726
rect 1690 1686 1693 1733
rect 1682 1683 1693 1686
rect 1682 1663 1685 1683
rect 1706 1646 1709 1736
rect 1714 1733 1717 1746
rect 1722 1743 1733 1746
rect 1722 1696 1725 1743
rect 1730 1733 1741 1736
rect 1730 1703 1733 1726
rect 1722 1693 1733 1696
rect 1682 1623 1685 1646
rect 1706 1643 1717 1646
rect 1690 1616 1693 1636
rect 1714 1623 1717 1643
rect 1690 1613 1717 1616
rect 1602 1543 1613 1546
rect 1514 1503 1517 1526
rect 1522 1513 1525 1526
rect 1530 1523 1541 1526
rect 1546 1523 1557 1526
rect 1538 1503 1541 1516
rect 1482 1423 1493 1426
rect 1290 1373 1297 1376
rect 1258 1346 1261 1366
rect 1254 1343 1261 1346
rect 1090 1263 1093 1336
rect 1074 1253 1085 1256
rect 1066 1196 1069 1216
rect 1074 1213 1077 1246
rect 1082 1203 1085 1253
rect 1090 1206 1093 1256
rect 1098 1223 1101 1286
rect 1106 1233 1109 1336
rect 1114 1273 1133 1276
rect 1114 1226 1117 1273
rect 1106 1223 1117 1226
rect 1106 1215 1109 1223
rect 1090 1203 1109 1206
rect 1114 1203 1117 1216
rect 1122 1206 1125 1266
rect 1130 1223 1133 1273
rect 1162 1226 1165 1336
rect 1170 1316 1173 1326
rect 1186 1316 1189 1336
rect 1170 1313 1189 1316
rect 1194 1303 1197 1326
rect 1218 1293 1221 1326
rect 1226 1303 1229 1326
rect 1138 1223 1165 1226
rect 1138 1213 1141 1223
rect 1146 1213 1157 1216
rect 1122 1203 1141 1206
rect 1066 1193 1073 1196
rect 1070 1126 1073 1193
rect 1066 1123 1073 1126
rect 1066 1106 1069 1123
rect 1050 1103 1069 1106
rect 978 1033 997 1036
rect 930 933 933 976
rect 978 973 981 1033
rect 986 986 989 1026
rect 1002 1006 1005 1056
rect 1010 1013 1013 1026
rect 1026 1013 1029 1036
rect 994 1003 1005 1006
rect 1018 993 1021 1006
rect 1034 1003 1037 1076
rect 986 983 1005 986
rect 938 953 949 956
rect 930 873 933 926
rect 938 883 941 953
rect 914 863 933 866
rect 890 813 901 816
rect 906 813 909 856
rect 878 803 885 806
rect 898 803 901 813
rect 878 746 881 803
rect 874 743 881 746
rect 874 686 877 743
rect 866 683 877 686
rect 866 603 869 683
rect 834 573 861 576
rect 834 533 837 573
rect 794 506 797 526
rect 842 506 845 566
rect 874 546 877 666
rect 882 653 885 726
rect 890 713 893 736
rect 898 633 901 726
rect 906 663 909 806
rect 914 673 917 806
rect 922 803 925 826
rect 930 813 933 863
rect 938 783 941 806
rect 946 803 949 926
rect 954 913 957 936
rect 962 923 965 946
rect 970 896 973 936
rect 978 933 997 936
rect 1002 933 1005 983
rect 1010 943 1013 956
rect 994 926 997 933
rect 986 913 989 926
rect 994 923 1005 926
rect 1018 916 1021 986
rect 1026 923 1029 966
rect 1042 943 1045 1046
rect 1050 963 1053 1103
rect 1058 993 1061 1006
rect 1066 986 1069 1016
rect 1074 1003 1077 1036
rect 1082 1016 1085 1136
rect 1106 1113 1109 1136
rect 1130 1073 1133 1196
rect 1138 1043 1141 1203
rect 1154 1173 1157 1206
rect 1162 1166 1165 1216
rect 1170 1203 1173 1226
rect 1082 1013 1109 1016
rect 1082 1003 1093 1006
rect 1098 986 1101 1006
rect 1106 996 1109 1013
rect 1114 1003 1117 1016
rect 1122 1013 1125 1026
rect 1146 1023 1149 1166
rect 1162 1163 1173 1166
rect 1154 1086 1157 1126
rect 1170 1096 1173 1163
rect 1178 1136 1181 1206
rect 1226 1203 1229 1236
rect 1234 1213 1237 1226
rect 1234 1193 1237 1206
rect 1242 1156 1245 1336
rect 1254 1246 1257 1343
rect 1274 1333 1285 1336
rect 1254 1243 1261 1246
rect 1250 1203 1253 1226
rect 1258 1196 1261 1243
rect 1266 1233 1269 1326
rect 1282 1313 1285 1326
rect 1194 1153 1245 1156
rect 1250 1193 1261 1196
rect 1194 1136 1197 1153
rect 1178 1133 1197 1136
rect 1250 1133 1253 1193
rect 1258 1133 1261 1146
rect 1186 1106 1189 1126
rect 1266 1116 1269 1216
rect 1282 1213 1285 1236
rect 1274 1203 1285 1206
rect 1290 1176 1293 1373
rect 1298 1323 1301 1336
rect 1346 1303 1349 1336
rect 1370 1333 1373 1346
rect 1354 1313 1357 1326
rect 1362 1316 1365 1326
rect 1378 1323 1381 1366
rect 1386 1343 1413 1346
rect 1386 1333 1389 1343
rect 1394 1333 1405 1336
rect 1394 1316 1397 1326
rect 1402 1323 1405 1333
rect 1362 1313 1397 1316
rect 1410 1313 1413 1343
rect 1458 1333 1461 1366
rect 1482 1356 1485 1423
rect 1522 1413 1525 1446
rect 1546 1403 1549 1523
rect 1586 1493 1589 1536
rect 1610 1486 1613 1543
rect 1618 1523 1621 1606
rect 1626 1596 1629 1606
rect 1658 1603 1669 1606
rect 1626 1593 1669 1596
rect 1682 1593 1685 1606
rect 1690 1603 1701 1606
rect 1586 1483 1613 1486
rect 1562 1433 1581 1436
rect 1562 1413 1565 1433
rect 1570 1413 1573 1426
rect 1578 1423 1581 1433
rect 1586 1413 1589 1483
rect 1602 1423 1613 1426
rect 1562 1393 1565 1406
rect 1626 1376 1629 1406
rect 1642 1403 1645 1476
rect 1666 1426 1669 1593
rect 1714 1586 1717 1606
rect 1722 1603 1725 1666
rect 1682 1583 1717 1586
rect 1682 1533 1685 1583
rect 1690 1543 1717 1546
rect 1690 1523 1693 1543
rect 1698 1456 1701 1536
rect 1714 1513 1717 1543
rect 1722 1516 1725 1526
rect 1730 1523 1733 1693
rect 1738 1623 1741 1733
rect 1746 1703 1749 1736
rect 1754 1716 1757 1726
rect 1762 1723 1765 1736
rect 1754 1713 1781 1716
rect 1786 1713 1789 1736
rect 1746 1623 1749 1646
rect 1802 1626 1805 1753
rect 1826 1713 1829 1726
rect 1810 1633 1813 1656
rect 1802 1623 1813 1626
rect 1786 1613 1797 1616
rect 1786 1593 1789 1606
rect 1802 1593 1805 1616
rect 1746 1563 1789 1566
rect 1746 1533 1749 1563
rect 1722 1513 1749 1516
rect 1690 1453 1701 1456
rect 1666 1423 1677 1426
rect 1666 1376 1669 1416
rect 1626 1373 1669 1376
rect 1674 1373 1677 1423
rect 1690 1403 1693 1453
rect 1466 1353 1485 1356
rect 1282 1173 1293 1176
rect 1274 1123 1277 1136
rect 1282 1123 1285 1173
rect 1290 1133 1293 1156
rect 1298 1116 1301 1206
rect 1346 1203 1349 1226
rect 1362 1213 1365 1246
rect 1410 1233 1445 1236
rect 1410 1186 1413 1233
rect 1418 1203 1421 1216
rect 1434 1213 1437 1226
rect 1410 1183 1421 1186
rect 1354 1133 1357 1146
rect 1410 1133 1413 1176
rect 1186 1103 1197 1106
rect 1170 1093 1181 1096
rect 1154 1083 1169 1086
rect 1166 1026 1169 1083
rect 1178 1053 1181 1093
rect 1194 1046 1197 1103
rect 1186 1043 1197 1046
rect 1166 1023 1173 1026
rect 1122 1003 1133 1006
rect 1138 996 1141 1006
rect 1106 993 1141 996
rect 1066 983 1101 986
rect 1034 933 1045 936
rect 1002 913 1021 916
rect 1034 903 1037 926
rect 970 893 989 896
rect 930 733 933 746
rect 922 686 925 716
rect 930 693 933 726
rect 938 686 941 736
rect 946 713 949 726
rect 922 683 941 686
rect 898 606 901 616
rect 906 613 909 646
rect 874 543 885 546
rect 858 513 861 536
rect 786 503 797 506
rect 826 503 845 506
rect 786 456 789 503
rect 786 453 797 456
rect 698 413 701 426
rect 706 413 709 436
rect 722 413 725 443
rect 794 436 797 453
rect 794 433 805 436
rect 786 416 789 426
rect 762 413 805 416
rect 706 403 717 406
rect 722 383 725 406
rect 746 403 757 406
rect 666 333 685 336
rect 706 333 709 356
rect 730 346 733 396
rect 714 343 733 346
rect 762 343 765 396
rect 778 393 781 406
rect 786 343 789 396
rect 794 336 797 396
rect 738 333 757 336
rect 778 333 797 336
rect 650 216 653 246
rect 674 223 677 326
rect 682 313 685 326
rect 714 323 733 326
rect 730 283 733 323
rect 754 313 757 326
rect 618 213 637 216
rect 650 213 677 216
rect 706 213 709 226
rect 722 213 725 236
rect 594 153 597 206
rect 610 203 637 206
rect 650 203 653 213
rect 610 123 613 203
rect 674 166 677 206
rect 682 203 693 206
rect 674 163 693 166
rect 698 163 701 206
rect 730 203 733 276
rect 762 273 765 326
rect 778 283 781 333
rect 786 323 805 326
rect 802 283 805 323
rect 738 196 741 216
rect 746 203 749 266
rect 762 216 765 246
rect 770 223 773 236
rect 738 193 749 196
rect 754 193 757 216
rect 762 213 773 216
rect 770 203 773 213
rect 778 203 781 226
rect 810 213 813 456
rect 826 326 829 503
rect 842 446 845 496
rect 882 483 885 543
rect 838 443 845 446
rect 838 396 841 443
rect 850 403 853 436
rect 866 433 869 476
rect 874 413 877 426
rect 858 403 877 406
rect 838 393 845 396
rect 834 333 837 346
rect 842 333 845 393
rect 882 373 885 396
rect 818 223 821 326
rect 826 323 845 326
rect 826 313 837 316
rect 826 223 829 276
rect 834 233 837 256
rect 642 123 645 156
rect 666 133 669 146
rect 690 123 693 163
rect 746 123 749 193
rect 794 183 797 206
rect 826 166 829 206
rect 834 193 837 226
rect 842 213 845 323
rect 850 306 853 326
rect 858 313 861 326
rect 866 323 869 356
rect 890 336 893 606
rect 898 603 909 606
rect 898 523 901 546
rect 898 393 901 416
rect 906 396 909 603
rect 922 583 925 626
rect 938 473 941 556
rect 946 533 949 636
rect 930 406 933 416
rect 922 403 933 406
rect 954 403 957 836
rect 962 813 965 876
rect 970 733 973 816
rect 962 663 965 726
rect 970 673 973 726
rect 978 696 981 886
rect 986 813 989 893
rect 1002 806 1005 866
rect 1010 813 1013 856
rect 986 796 989 806
rect 1002 803 1013 806
rect 1018 796 1021 846
rect 1026 823 1029 836
rect 1034 823 1037 896
rect 1042 866 1045 933
rect 1050 913 1053 936
rect 1058 923 1061 946
rect 1066 873 1069 936
rect 1042 863 1053 866
rect 1042 833 1045 856
rect 1050 833 1053 863
rect 1074 853 1077 936
rect 1082 923 1085 966
rect 1106 936 1109 976
rect 1098 933 1109 936
rect 1090 896 1093 926
rect 1098 903 1101 926
rect 1106 916 1109 933
rect 1114 923 1117 946
rect 1122 923 1125 936
rect 1138 926 1141 993
rect 1146 933 1149 986
rect 1138 923 1149 926
rect 1154 923 1157 1016
rect 1170 1003 1173 1023
rect 1146 916 1149 923
rect 1106 913 1117 916
rect 1122 913 1141 916
rect 1146 913 1153 916
rect 1090 893 1109 896
rect 1090 856 1093 893
rect 1082 853 1093 856
rect 1082 846 1085 853
rect 1066 843 1085 846
rect 1050 823 1061 826
rect 1066 816 1069 843
rect 1090 816 1093 846
rect 986 793 1021 796
rect 1026 813 1069 816
rect 1026 786 1029 813
rect 1010 783 1029 786
rect 1042 776 1045 786
rect 1026 773 1045 776
rect 1074 773 1077 816
rect 1082 813 1093 816
rect 986 723 989 746
rect 978 693 989 696
rect 962 573 965 646
rect 970 593 973 616
rect 986 603 989 693
rect 994 683 997 736
rect 1002 733 1005 766
rect 1010 733 1021 736
rect 1002 723 1012 726
rect 994 576 997 636
rect 978 573 997 576
rect 962 513 965 526
rect 970 453 973 556
rect 978 436 981 573
rect 986 533 989 546
rect 994 533 997 566
rect 1002 523 1005 723
rect 1018 706 1021 733
rect 1010 703 1021 706
rect 1026 703 1029 773
rect 1034 723 1037 746
rect 1058 743 1061 766
rect 1074 733 1077 746
rect 1074 716 1077 726
rect 1082 723 1085 813
rect 1090 716 1093 806
rect 1098 763 1101 836
rect 1106 806 1109 893
rect 1114 813 1117 913
rect 1138 833 1141 913
rect 1150 846 1153 913
rect 1150 843 1157 846
rect 1162 843 1165 996
rect 1178 973 1181 1026
rect 1186 993 1189 1043
rect 1122 823 1149 826
rect 1122 813 1125 823
rect 1106 803 1125 806
rect 1130 803 1133 816
rect 1098 723 1101 756
rect 1114 723 1117 736
rect 1034 713 1045 716
rect 1050 713 1077 716
rect 1082 713 1101 716
rect 1082 706 1085 713
rect 1074 703 1085 706
rect 1010 613 1013 703
rect 1018 613 1021 626
rect 1026 613 1029 686
rect 1034 623 1037 656
rect 1042 633 1045 696
rect 1074 646 1077 703
rect 1138 686 1141 816
rect 1146 693 1149 766
rect 1106 683 1141 686
rect 1050 643 1077 646
rect 1010 603 1021 606
rect 1042 603 1045 616
rect 1050 603 1053 643
rect 1058 596 1061 636
rect 1010 533 1013 596
rect 1042 593 1061 596
rect 1026 533 1029 576
rect 1066 563 1069 616
rect 1074 603 1077 643
rect 1066 543 1069 556
rect 1050 533 1069 536
rect 1018 523 1045 526
rect 986 446 989 516
rect 1018 513 1021 523
rect 986 443 997 446
rect 978 433 989 436
rect 978 403 981 416
rect 906 393 917 396
rect 890 333 901 336
rect 914 333 917 393
rect 922 333 925 403
rect 930 393 933 403
rect 962 383 965 396
rect 930 353 949 356
rect 866 313 885 316
rect 866 306 869 313
rect 850 303 869 306
rect 874 293 877 306
rect 890 273 893 326
rect 898 323 909 326
rect 810 163 829 166
rect 762 133 765 146
rect 810 123 813 163
rect 850 123 853 216
rect 866 213 869 236
rect 882 146 885 226
rect 906 223 917 226
rect 922 223 925 326
rect 930 306 933 326
rect 946 323 949 353
rect 954 333 957 346
rect 978 336 981 356
rect 970 333 981 336
rect 986 333 989 433
rect 994 413 997 443
rect 1002 413 1005 426
rect 930 303 941 306
rect 938 226 941 303
rect 962 253 965 326
rect 938 223 949 226
rect 890 213 917 216
rect 890 203 893 213
rect 866 133 869 146
rect 882 143 893 146
rect 890 73 893 143
rect 914 123 917 206
rect 922 203 941 206
rect 946 203 949 223
rect 954 213 957 226
rect 970 213 973 326
rect 978 313 981 326
rect 986 293 989 326
rect 994 296 997 406
rect 1002 393 1005 406
rect 1002 303 1005 326
rect 1010 313 1013 336
rect 1018 333 1021 346
rect 994 293 1001 296
rect 978 213 981 266
rect 998 236 1001 293
rect 998 233 1005 236
rect 986 213 997 216
rect 938 196 941 203
rect 938 193 949 196
rect 946 123 949 193
rect 954 173 957 206
rect 962 123 965 146
rect 986 123 989 206
rect 1002 123 1005 233
rect 1010 213 1013 266
rect 1018 233 1021 326
rect 1026 303 1029 326
rect 1034 323 1037 506
rect 1050 503 1053 533
rect 1058 513 1061 526
rect 1074 486 1077 576
rect 1082 533 1085 626
rect 1090 623 1093 636
rect 1082 503 1085 526
rect 1058 483 1077 486
rect 1058 476 1061 483
rect 1050 473 1061 476
rect 1058 403 1061 473
rect 1066 403 1069 476
rect 1042 323 1045 396
rect 1074 393 1077 426
rect 1082 393 1085 446
rect 1090 363 1093 616
rect 1098 603 1101 676
rect 1098 573 1101 596
rect 1098 523 1101 546
rect 1106 516 1109 683
rect 1114 596 1117 666
rect 1122 603 1125 646
rect 1114 593 1125 596
rect 1114 533 1117 546
rect 1122 533 1125 593
rect 1130 523 1133 616
rect 1138 603 1141 676
rect 1154 633 1157 843
rect 1170 836 1173 936
rect 1194 913 1197 1026
rect 1226 976 1229 1116
rect 1266 1113 1301 1116
rect 1362 1113 1365 1126
rect 1266 1063 1269 1113
rect 1410 1096 1413 1126
rect 1386 1066 1389 1086
rect 1382 1063 1389 1066
rect 1210 973 1229 976
rect 1210 933 1213 973
rect 1250 966 1253 1046
rect 1274 1013 1277 1026
rect 1306 1013 1309 1046
rect 1314 1006 1317 1016
rect 1242 963 1253 966
rect 1306 1003 1317 1006
rect 1242 916 1245 963
rect 1258 923 1261 956
rect 1282 933 1301 936
rect 1282 916 1285 933
rect 1242 913 1249 916
rect 1162 833 1173 836
rect 1162 723 1165 833
rect 1170 813 1173 826
rect 1178 813 1181 836
rect 1186 806 1189 856
rect 1194 813 1197 826
rect 1202 806 1205 906
rect 1246 856 1249 913
rect 1278 913 1285 916
rect 1246 853 1253 856
rect 1250 836 1253 853
rect 1170 803 1189 806
rect 1194 803 1205 806
rect 1210 803 1213 816
rect 1194 796 1197 803
rect 1186 793 1197 796
rect 1186 736 1189 793
rect 1182 733 1189 736
rect 1182 676 1185 733
rect 1194 713 1197 726
rect 1182 673 1189 676
rect 1186 653 1189 673
rect 1138 533 1141 576
rect 1146 523 1149 626
rect 1154 583 1157 606
rect 1170 593 1173 646
rect 1194 613 1197 676
rect 1202 586 1205 796
rect 1218 773 1221 826
rect 1226 813 1229 836
rect 1234 833 1253 836
rect 1242 746 1245 826
rect 1258 823 1261 866
rect 1278 856 1281 913
rect 1278 853 1285 856
rect 1290 853 1293 926
rect 1306 923 1309 1003
rect 1322 986 1325 1056
rect 1346 1003 1349 1026
rect 1314 916 1317 986
rect 1322 983 1337 986
rect 1322 933 1325 956
rect 1298 913 1317 916
rect 1282 836 1285 853
rect 1266 833 1293 836
rect 1266 813 1269 833
rect 1258 803 1269 806
rect 1226 743 1245 746
rect 1162 583 1173 586
rect 1194 583 1205 586
rect 1210 583 1213 726
rect 1218 713 1221 726
rect 1226 656 1229 743
rect 1218 653 1229 656
rect 1102 513 1109 516
rect 1102 446 1105 513
rect 1098 443 1105 446
rect 1098 413 1101 443
rect 1114 413 1117 516
rect 1162 496 1165 583
rect 1194 566 1197 583
rect 1218 566 1221 653
rect 1234 643 1237 736
rect 1242 713 1245 726
rect 1250 676 1253 756
rect 1258 723 1261 736
rect 1266 706 1269 803
rect 1282 746 1285 826
rect 1290 813 1293 826
rect 1242 673 1253 676
rect 1262 703 1269 706
rect 1186 556 1189 566
rect 1194 563 1205 566
rect 1218 563 1229 566
rect 1186 553 1197 556
rect 1186 523 1189 546
rect 1154 493 1165 496
rect 1122 413 1125 426
rect 1130 413 1133 486
rect 1138 366 1141 436
rect 1154 376 1157 493
rect 1194 456 1197 553
rect 1202 523 1205 563
rect 1154 373 1165 376
rect 1138 363 1145 366
rect 1050 333 1053 356
rect 1074 333 1077 356
rect 1058 306 1061 326
rect 1122 313 1125 326
rect 1142 316 1145 363
rect 1162 353 1165 373
rect 1138 313 1145 316
rect 1042 303 1061 306
rect 1018 206 1021 226
rect 1010 203 1021 206
rect 1026 203 1029 296
rect 1034 216 1037 256
rect 1042 223 1045 303
rect 1034 213 1045 216
rect 1026 153 1029 196
rect 1042 123 1045 206
rect 1050 203 1053 236
rect 1050 183 1053 196
rect 1058 193 1061 296
rect 1074 276 1077 306
rect 1138 293 1141 313
rect 1066 163 1069 276
rect 1074 273 1081 276
rect 1078 176 1081 273
rect 1154 246 1157 326
rect 1138 243 1157 246
rect 1138 223 1141 243
rect 1162 236 1165 336
rect 1170 323 1173 456
rect 1194 453 1201 456
rect 1178 283 1181 416
rect 1186 403 1189 446
rect 1198 396 1201 453
rect 1194 393 1201 396
rect 1194 373 1197 393
rect 1210 353 1213 556
rect 1226 516 1229 563
rect 1234 526 1237 576
rect 1242 533 1245 673
rect 1250 613 1253 666
rect 1262 626 1265 703
rect 1262 623 1269 626
rect 1250 603 1261 606
rect 1234 523 1245 526
rect 1250 523 1253 603
rect 1266 596 1269 623
rect 1258 593 1269 596
rect 1274 593 1277 746
rect 1282 743 1293 746
rect 1282 703 1285 736
rect 1282 613 1285 626
rect 1290 613 1293 743
rect 1298 713 1301 913
rect 1334 906 1337 983
rect 1370 966 1373 1026
rect 1346 963 1373 966
rect 1346 913 1349 963
rect 1382 956 1385 1063
rect 1362 933 1365 956
rect 1382 953 1389 956
rect 1334 903 1341 906
rect 1306 773 1309 886
rect 1314 726 1317 826
rect 1322 823 1325 846
rect 1330 813 1333 836
rect 1338 813 1341 903
rect 1346 756 1349 826
rect 1362 783 1365 926
rect 1386 863 1389 953
rect 1394 923 1397 1096
rect 1406 1093 1413 1096
rect 1406 1026 1409 1093
rect 1418 1033 1421 1183
rect 1426 1176 1429 1206
rect 1442 1203 1445 1233
rect 1450 1213 1453 1246
rect 1450 1193 1453 1206
rect 1458 1186 1461 1326
rect 1466 1233 1469 1353
rect 1474 1303 1477 1326
rect 1482 1313 1485 1336
rect 1530 1333 1533 1346
rect 1538 1333 1557 1336
rect 1490 1213 1493 1246
rect 1514 1243 1517 1326
rect 1530 1313 1533 1326
rect 1554 1323 1557 1333
rect 1554 1303 1557 1316
rect 1586 1306 1589 1326
rect 1582 1303 1589 1306
rect 1582 1246 1585 1303
rect 1594 1293 1597 1326
rect 1610 1303 1613 1336
rect 1514 1233 1549 1236
rect 1506 1203 1509 1226
rect 1458 1183 1469 1186
rect 1426 1173 1445 1176
rect 1426 1106 1429 1136
rect 1434 1123 1437 1146
rect 1442 1133 1445 1173
rect 1450 1113 1453 1126
rect 1458 1123 1461 1136
rect 1466 1116 1469 1183
rect 1514 1153 1517 1233
rect 1514 1133 1517 1146
rect 1522 1126 1525 1226
rect 1546 1213 1549 1233
rect 1554 1213 1557 1246
rect 1570 1243 1585 1246
rect 1458 1113 1469 1116
rect 1514 1123 1525 1126
rect 1458 1106 1461 1113
rect 1426 1103 1461 1106
rect 1406 1023 1413 1026
rect 1410 1003 1413 1023
rect 1458 1003 1461 1103
rect 1514 1096 1517 1123
rect 1506 1093 1517 1096
rect 1482 1013 1485 1026
rect 1490 1006 1493 1036
rect 1506 1026 1509 1093
rect 1506 1023 1517 1026
rect 1514 1006 1517 1023
rect 1522 1013 1525 1086
rect 1530 1056 1533 1136
rect 1538 1123 1541 1146
rect 1546 1133 1549 1156
rect 1570 1133 1573 1243
rect 1594 1213 1597 1226
rect 1626 1213 1629 1326
rect 1658 1286 1661 1326
rect 1666 1293 1669 1326
rect 1658 1283 1677 1286
rect 1658 1226 1661 1283
rect 1578 1173 1581 1206
rect 1586 1203 1597 1206
rect 1642 1203 1645 1226
rect 1658 1223 1665 1226
rect 1650 1203 1653 1216
rect 1662 1176 1665 1223
rect 1658 1173 1665 1176
rect 1658 1156 1661 1173
rect 1626 1153 1661 1156
rect 1530 1053 1549 1056
rect 1482 973 1485 1006
rect 1490 1003 1501 1006
rect 1514 1003 1533 1006
rect 1490 966 1493 996
rect 1482 963 1493 966
rect 1410 923 1413 956
rect 1442 883 1445 926
rect 1450 853 1453 936
rect 1458 923 1461 946
rect 1474 933 1477 956
rect 1458 896 1461 916
rect 1458 893 1469 896
rect 1370 793 1373 806
rect 1386 793 1389 816
rect 1394 803 1397 836
rect 1402 833 1421 836
rect 1402 803 1405 833
rect 1426 826 1429 846
rect 1466 836 1469 893
rect 1482 883 1485 963
rect 1498 926 1501 996
rect 1490 923 1501 926
rect 1506 933 1525 936
rect 1458 833 1469 836
rect 1418 823 1429 826
rect 1394 783 1397 796
rect 1410 793 1413 816
rect 1418 776 1421 823
rect 1426 813 1437 816
rect 1442 793 1445 826
rect 1450 783 1453 806
rect 1322 743 1325 756
rect 1330 753 1349 756
rect 1306 723 1317 726
rect 1322 723 1325 736
rect 1330 726 1333 753
rect 1338 743 1365 746
rect 1338 733 1341 743
rect 1330 723 1341 726
rect 1258 553 1293 556
rect 1226 513 1241 516
rect 1218 376 1221 416
rect 1226 393 1229 486
rect 1238 446 1241 513
rect 1238 443 1245 446
rect 1234 403 1237 426
rect 1242 396 1245 443
rect 1250 413 1253 466
rect 1258 453 1261 553
rect 1266 436 1269 536
rect 1274 513 1277 526
rect 1258 433 1269 436
rect 1258 413 1261 433
rect 1266 413 1269 426
rect 1282 413 1285 546
rect 1290 533 1293 553
rect 1290 506 1293 526
rect 1298 523 1301 666
rect 1306 656 1309 723
rect 1314 683 1317 716
rect 1338 676 1341 723
rect 1346 703 1349 736
rect 1362 733 1365 743
rect 1394 733 1397 776
rect 1410 773 1421 776
rect 1458 773 1461 833
rect 1466 776 1469 806
rect 1482 803 1485 826
rect 1490 793 1493 923
rect 1498 903 1501 916
rect 1506 913 1509 933
rect 1514 913 1517 926
rect 1498 826 1501 896
rect 1506 833 1509 906
rect 1522 893 1525 933
rect 1530 913 1533 976
rect 1538 943 1541 1016
rect 1546 1013 1549 1053
rect 1554 1033 1557 1126
rect 1578 1103 1581 1126
rect 1586 1046 1589 1136
rect 1594 1113 1597 1126
rect 1586 1043 1597 1046
rect 1546 993 1549 1006
rect 1570 993 1573 1006
rect 1594 976 1597 1043
rect 1602 1023 1605 1136
rect 1626 1133 1629 1153
rect 1674 1133 1677 1276
rect 1682 1213 1685 1336
rect 1690 1306 1693 1396
rect 1722 1393 1725 1416
rect 1738 1406 1741 1486
rect 1762 1473 1765 1536
rect 1786 1523 1789 1563
rect 1802 1426 1805 1496
rect 1810 1486 1813 1623
rect 1818 1613 1821 1636
rect 1826 1566 1829 1626
rect 1858 1623 1861 1636
rect 1866 1616 1869 1816
rect 1874 1793 1877 1806
rect 1890 1756 1893 1806
rect 1898 1796 1901 1906
rect 1994 1896 1997 1973
rect 1978 1893 1997 1896
rect 1906 1813 1933 1816
rect 1914 1803 1933 1806
rect 1898 1793 1925 1796
rect 1882 1753 1893 1756
rect 1882 1733 1885 1753
rect 1874 1723 1885 1726
rect 1898 1706 1901 1786
rect 1834 1603 1837 1616
rect 1842 1613 1869 1616
rect 1882 1703 1901 1706
rect 1826 1563 1833 1566
rect 1810 1483 1821 1486
rect 1802 1423 1813 1426
rect 1746 1413 1805 1416
rect 1738 1403 1765 1406
rect 1698 1326 1701 1376
rect 1794 1366 1797 1406
rect 1802 1373 1805 1413
rect 1810 1366 1813 1423
rect 1818 1403 1821 1483
rect 1830 1396 1833 1563
rect 1850 1533 1853 1596
rect 1842 1513 1845 1526
rect 1858 1523 1861 1613
rect 1866 1583 1869 1606
rect 1882 1593 1885 1703
rect 1922 1686 1925 1793
rect 1930 1786 1933 1803
rect 1946 1793 1949 1806
rect 1930 1783 1937 1786
rect 1918 1683 1925 1686
rect 1906 1583 1909 1616
rect 1918 1566 1921 1683
rect 1934 1676 1937 1783
rect 1978 1746 1981 1893
rect 2042 1886 2045 1926
rect 2074 1913 2077 1996
rect 2146 1976 2149 2026
rect 2106 1973 2149 1976
rect 2154 2023 2165 2026
rect 2178 2043 2205 2046
rect 2258 2093 2269 2096
rect 2082 1886 2085 1926
rect 2090 1916 2093 1936
rect 2106 1923 2109 1973
rect 2114 1943 2141 1946
rect 2114 1933 2117 1943
rect 2122 1916 2125 1926
rect 2090 1913 2125 1916
rect 2042 1883 2085 1886
rect 2130 1906 2133 1936
rect 2138 1933 2141 1943
rect 2138 1913 2141 1926
rect 2154 1906 2157 2023
rect 2162 1923 2165 2016
rect 2178 2013 2181 2043
rect 2194 2023 2197 2036
rect 2258 2026 2261 2093
rect 2274 2076 2277 2136
rect 2282 2133 2285 2163
rect 2338 2136 2341 2216
rect 2370 2213 2373 2256
rect 2466 2253 2469 2316
rect 2522 2313 2533 2316
rect 2394 2223 2397 2236
rect 2426 2213 2429 2226
rect 2442 2213 2445 2236
rect 2522 2226 2525 2313
rect 2450 2206 2453 2226
rect 2346 2193 2349 2206
rect 2338 2133 2349 2136
rect 2362 2133 2365 2206
rect 2442 2203 2453 2206
rect 2418 2133 2421 2186
rect 2474 2176 2477 2226
rect 2522 2223 2533 2226
rect 2450 2173 2477 2176
rect 2450 2136 2453 2173
rect 2450 2133 2461 2136
rect 2298 2103 2301 2116
rect 2274 2073 2309 2076
rect 2234 2013 2237 2026
rect 2258 2023 2269 2026
rect 2170 1976 2173 2006
rect 2170 1973 2205 1976
rect 2178 1943 2197 1946
rect 2178 1923 2181 1943
rect 2186 1923 2189 1936
rect 2194 1933 2197 1943
rect 2130 1903 2157 1906
rect 2202 1903 2205 1973
rect 2250 1933 2253 1956
rect 2266 1946 2269 2023
rect 2274 2013 2277 2066
rect 2282 2023 2301 2026
rect 2282 1966 2285 2023
rect 2290 1996 2293 2016
rect 2298 2003 2301 2023
rect 2306 2013 2309 2073
rect 2338 2063 2341 2116
rect 2402 2086 2405 2126
rect 2442 2086 2445 2126
rect 2402 2083 2445 2086
rect 2458 2076 2461 2133
rect 2498 2123 2501 2136
rect 2450 2073 2461 2076
rect 2330 2053 2373 2056
rect 2330 2013 2333 2053
rect 2370 2013 2373 2053
rect 2450 2033 2453 2073
rect 2426 2013 2429 2026
rect 2434 2023 2469 2026
rect 2306 1996 2309 2006
rect 2290 1993 2309 1996
rect 2282 1963 2293 1966
rect 2346 1963 2349 2006
rect 2266 1943 2277 1946
rect 2234 1913 2237 1926
rect 2026 1853 2069 1856
rect 2002 1763 2005 1806
rect 2010 1756 2013 1816
rect 2026 1813 2029 1853
rect 2066 1813 2069 1853
rect 2130 1833 2133 1903
rect 2178 1816 2181 1836
rect 2042 1783 2045 1806
rect 1970 1743 1981 1746
rect 2002 1753 2013 1756
rect 1946 1703 1949 1726
rect 1930 1673 1937 1676
rect 1918 1563 1925 1566
rect 1850 1403 1853 1476
rect 1874 1413 1877 1536
rect 1882 1523 1885 1536
rect 1794 1363 1813 1366
rect 1826 1393 1833 1396
rect 1714 1343 1733 1346
rect 1714 1336 1717 1343
rect 1706 1333 1717 1336
rect 1698 1323 1709 1326
rect 1690 1303 1697 1306
rect 1694 1236 1697 1303
rect 1694 1233 1701 1236
rect 1690 1083 1693 1226
rect 1698 1116 1701 1233
rect 1706 1133 1709 1323
rect 1714 1283 1717 1326
rect 1722 1273 1725 1336
rect 1730 1333 1733 1343
rect 1778 1333 1781 1346
rect 1786 1333 1821 1336
rect 1826 1333 1829 1393
rect 1842 1333 1845 1376
rect 1882 1366 1885 1516
rect 1890 1496 1893 1556
rect 1898 1513 1901 1546
rect 1890 1493 1897 1496
rect 1874 1363 1885 1366
rect 1762 1236 1765 1326
rect 1714 1233 1765 1236
rect 1714 1193 1717 1233
rect 1786 1226 1789 1333
rect 1802 1323 1853 1326
rect 1730 1213 1733 1226
rect 1722 1116 1725 1136
rect 1730 1133 1733 1146
rect 1746 1123 1749 1216
rect 1770 1206 1773 1226
rect 1762 1203 1773 1206
rect 1778 1223 1789 1226
rect 1762 1156 1765 1203
rect 1762 1153 1773 1156
rect 1754 1116 1757 1136
rect 1698 1113 1705 1116
rect 1702 1046 1705 1113
rect 1714 1103 1717 1116
rect 1722 1113 1757 1116
rect 1770 1096 1773 1153
rect 1698 1043 1705 1046
rect 1762 1093 1773 1096
rect 1762 1046 1765 1093
rect 1762 1043 1773 1046
rect 1578 973 1597 976
rect 1538 923 1541 936
rect 1554 933 1557 956
rect 1570 936 1573 946
rect 1562 933 1573 936
rect 1498 823 1509 826
rect 1514 823 1517 846
rect 1522 823 1525 836
rect 1538 823 1541 886
rect 1546 873 1549 926
rect 1562 866 1565 933
rect 1570 913 1573 926
rect 1578 886 1581 973
rect 1586 923 1589 956
rect 1594 916 1597 926
rect 1546 863 1565 866
rect 1570 883 1581 886
rect 1586 913 1597 916
rect 1506 786 1509 823
rect 1514 813 1525 816
rect 1546 806 1549 863
rect 1466 773 1473 776
rect 1338 673 1349 676
rect 1362 673 1365 726
rect 1370 713 1389 716
rect 1386 696 1389 713
rect 1394 706 1397 726
rect 1402 723 1405 736
rect 1394 703 1405 706
rect 1386 693 1397 696
rect 1306 653 1317 656
rect 1306 613 1309 646
rect 1314 596 1317 653
rect 1322 623 1325 666
rect 1330 613 1333 636
rect 1310 593 1317 596
rect 1322 593 1333 596
rect 1310 526 1313 593
rect 1322 543 1325 593
rect 1330 536 1333 586
rect 1322 533 1333 536
rect 1310 523 1317 526
rect 1290 503 1297 506
rect 1294 416 1297 503
rect 1306 423 1309 506
rect 1314 416 1317 523
rect 1322 503 1325 533
rect 1338 426 1341 616
rect 1346 613 1349 673
rect 1378 633 1381 646
rect 1362 623 1381 626
rect 1394 623 1397 693
rect 1354 603 1357 616
rect 1362 603 1365 623
rect 1370 603 1373 616
rect 1378 606 1381 623
rect 1402 613 1405 666
rect 1378 603 1397 606
rect 1354 563 1357 596
rect 1346 493 1349 556
rect 1362 526 1365 536
rect 1370 533 1373 546
rect 1354 523 1365 526
rect 1370 523 1381 526
rect 1386 523 1389 576
rect 1394 533 1397 596
rect 1410 546 1413 773
rect 1418 763 1461 766
rect 1418 733 1421 763
rect 1418 673 1421 716
rect 1434 646 1437 736
rect 1458 723 1461 763
rect 1470 716 1473 773
rect 1466 713 1473 716
rect 1466 656 1469 713
rect 1482 693 1485 786
rect 1498 783 1509 786
rect 1514 803 1549 806
rect 1498 673 1501 783
rect 1466 653 1501 656
rect 1418 583 1421 646
rect 1434 643 1469 646
rect 1426 623 1445 626
rect 1450 623 1453 636
rect 1426 613 1429 623
rect 1426 576 1429 606
rect 1418 573 1429 576
rect 1434 573 1437 616
rect 1442 613 1445 623
rect 1450 583 1453 606
rect 1402 543 1413 546
rect 1418 563 1461 566
rect 1418 533 1421 563
rect 1434 533 1437 556
rect 1354 436 1357 523
rect 1362 503 1365 516
rect 1394 463 1397 526
rect 1418 513 1421 526
rect 1354 433 1373 436
rect 1290 413 1297 416
rect 1306 413 1317 416
rect 1322 423 1349 426
rect 1234 393 1245 396
rect 1218 373 1229 376
rect 1218 343 1221 366
rect 1226 336 1229 373
rect 1186 313 1189 336
rect 1194 333 1213 336
rect 1218 333 1229 336
rect 1218 323 1221 333
rect 1234 263 1237 393
rect 1250 386 1253 406
rect 1242 383 1253 386
rect 1242 333 1245 383
rect 1146 233 1165 236
rect 1146 216 1149 233
rect 1114 213 1149 216
rect 1154 223 1189 226
rect 1154 213 1157 223
rect 1170 213 1181 216
rect 1186 213 1189 223
rect 1194 213 1205 216
rect 1074 173 1081 176
rect 1090 173 1093 206
rect 1074 153 1077 173
rect 1058 133 1061 146
rect 1106 123 1109 206
rect 1122 133 1125 206
rect 1130 183 1133 206
rect 1138 203 1141 213
rect 1210 206 1213 256
rect 1146 173 1149 206
rect 1162 166 1165 206
rect 1138 123 1141 166
rect 1162 163 1173 166
rect 1170 146 1173 163
rect 1178 156 1181 206
rect 1186 203 1229 206
rect 1242 203 1245 326
rect 1178 153 1189 156
rect 1202 153 1205 196
rect 1154 133 1157 146
rect 1170 143 1181 146
rect 1178 123 1181 143
rect 1186 123 1189 153
rect 1226 146 1229 203
rect 1242 176 1245 196
rect 1250 193 1253 356
rect 1258 336 1261 406
rect 1290 393 1293 413
rect 1306 346 1309 413
rect 1322 393 1325 423
rect 1330 413 1341 416
rect 1330 376 1333 413
rect 1338 383 1341 406
rect 1346 393 1349 423
rect 1330 373 1349 376
rect 1290 336 1293 346
rect 1298 343 1309 346
rect 1330 343 1333 366
rect 1298 336 1301 343
rect 1258 333 1269 336
rect 1290 333 1301 336
rect 1258 263 1261 326
rect 1266 323 1269 333
rect 1282 303 1285 316
rect 1258 233 1277 236
rect 1282 233 1285 256
rect 1290 233 1293 326
rect 1298 313 1301 333
rect 1306 323 1309 336
rect 1314 333 1325 336
rect 1330 316 1333 326
rect 1338 323 1341 336
rect 1346 316 1349 373
rect 1354 333 1357 366
rect 1362 326 1365 416
rect 1378 413 1381 426
rect 1386 413 1389 436
rect 1402 423 1405 496
rect 1426 423 1429 506
rect 1434 486 1437 526
rect 1458 523 1461 563
rect 1466 536 1469 643
rect 1490 586 1493 616
rect 1482 583 1493 586
rect 1466 533 1473 536
rect 1434 483 1445 486
rect 1434 423 1437 476
rect 1370 403 1413 406
rect 1418 393 1421 416
rect 1442 406 1445 483
rect 1458 453 1461 506
rect 1470 456 1473 533
rect 1482 486 1485 556
rect 1498 493 1501 653
rect 1506 593 1509 776
rect 1514 523 1517 803
rect 1522 733 1525 796
rect 1554 773 1557 836
rect 1562 796 1565 816
rect 1570 803 1573 883
rect 1578 813 1581 826
rect 1586 803 1589 913
rect 1602 896 1605 946
rect 1610 906 1613 1016
rect 1650 953 1653 1016
rect 1674 993 1677 1006
rect 1698 976 1701 1043
rect 1682 973 1701 976
rect 1682 956 1685 973
rect 1674 953 1685 956
rect 1618 943 1653 946
rect 1618 923 1621 936
rect 1626 933 1637 936
rect 1626 913 1629 926
rect 1642 906 1645 936
rect 1650 933 1653 943
rect 1674 936 1677 953
rect 1706 943 1709 1026
rect 1770 1023 1773 1043
rect 1722 973 1725 1016
rect 1754 1013 1773 1016
rect 1754 946 1757 1013
rect 1778 996 1781 1223
rect 1786 1126 1789 1216
rect 1802 1203 1805 1226
rect 1810 1216 1813 1316
rect 1874 1266 1877 1363
rect 1894 1356 1897 1493
rect 1914 1456 1917 1546
rect 1922 1533 1925 1563
rect 1922 1516 1925 1526
rect 1930 1523 1933 1673
rect 1962 1663 1965 1736
rect 1922 1513 1933 1516
rect 1914 1453 1921 1456
rect 1918 1376 1921 1453
rect 1930 1413 1933 1513
rect 1946 1493 1949 1596
rect 1962 1553 1965 1656
rect 1970 1616 1973 1743
rect 1978 1636 1981 1726
rect 1986 1713 1989 1736
rect 2002 1726 2005 1753
rect 2042 1736 2045 1776
rect 2018 1733 2029 1736
rect 2034 1733 2045 1736
rect 2114 1733 2117 1806
rect 2122 1773 2125 1816
rect 2170 1813 2181 1816
rect 2138 1783 2141 1806
rect 2170 1766 2173 1813
rect 2186 1776 2189 1816
rect 2218 1803 2221 1816
rect 2186 1773 2221 1776
rect 2026 1726 2029 1733
rect 1994 1723 2005 1726
rect 2010 1703 2013 1726
rect 2018 1713 2021 1726
rect 2026 1723 2037 1726
rect 2034 1693 2037 1723
rect 2042 1716 2045 1733
rect 2066 1723 2109 1726
rect 2042 1713 2061 1716
rect 2066 1713 2069 1723
rect 2122 1713 2125 1766
rect 2170 1763 2181 1766
rect 1978 1633 1989 1636
rect 1970 1613 1977 1616
rect 1974 1516 1977 1613
rect 1986 1603 1989 1633
rect 1970 1513 1977 1516
rect 1986 1513 1989 1526
rect 1970 1496 1973 1513
rect 1962 1493 1973 1496
rect 1890 1353 1897 1356
rect 1914 1373 1921 1376
rect 1962 1373 1965 1493
rect 1994 1453 1997 1666
rect 2002 1566 2005 1686
rect 2034 1613 2037 1636
rect 2058 1603 2061 1713
rect 2138 1646 2141 1716
rect 2114 1643 2141 1646
rect 2114 1613 2117 1643
rect 2130 1633 2141 1636
rect 2130 1613 2133 1633
rect 2146 1613 2149 1636
rect 2154 1623 2157 1636
rect 2002 1563 2021 1566
rect 2018 1496 2021 1563
rect 2058 1536 2061 1556
rect 2026 1503 2029 1526
rect 2034 1513 2037 1536
rect 2042 1523 2045 1536
rect 2058 1533 2069 1536
rect 2050 1523 2061 1526
rect 2090 1513 2093 1526
rect 2114 1503 2117 1536
rect 2122 1506 2125 1536
rect 2130 1523 2133 1606
rect 2154 1513 2157 1556
rect 2122 1503 2133 1506
rect 2018 1493 2045 1496
rect 2042 1426 2045 1493
rect 2034 1423 2045 1426
rect 2066 1426 2069 1456
rect 2066 1423 2077 1426
rect 1874 1263 1885 1266
rect 1818 1226 1821 1246
rect 1818 1223 1829 1226
rect 1810 1213 1829 1216
rect 1866 1213 1869 1226
rect 1810 1203 1821 1206
rect 1826 1186 1829 1213
rect 1822 1183 1829 1186
rect 1842 1183 1845 1206
rect 1874 1196 1877 1246
rect 1870 1193 1877 1196
rect 1786 1123 1813 1126
rect 1786 1003 1789 1076
rect 1802 1013 1805 1046
rect 1810 1013 1813 1123
rect 1822 1096 1825 1183
rect 1834 1133 1837 1156
rect 1870 1136 1873 1193
rect 1882 1163 1885 1263
rect 1890 1193 1893 1353
rect 1914 1336 1917 1373
rect 1906 1333 1917 1336
rect 1930 1333 1941 1336
rect 1906 1256 1909 1333
rect 1914 1316 1917 1326
rect 1938 1323 1941 1333
rect 1962 1316 1965 1326
rect 1978 1316 1981 1336
rect 1914 1313 1965 1316
rect 1974 1313 1981 1316
rect 1906 1253 1913 1256
rect 1910 1196 1913 1253
rect 1922 1203 1925 1216
rect 1910 1193 1925 1196
rect 1870 1133 1877 1136
rect 1890 1133 1893 1186
rect 1834 1113 1837 1126
rect 1842 1106 1845 1126
rect 1874 1116 1877 1133
rect 1834 1103 1845 1106
rect 1850 1113 1877 1116
rect 1914 1113 1917 1126
rect 1822 1093 1829 1096
rect 1826 1046 1829 1093
rect 1826 1043 1833 1046
rect 1818 1023 1821 1036
rect 1770 993 1781 996
rect 1802 993 1805 1006
rect 1770 983 1773 993
rect 1818 986 1821 1006
rect 1810 983 1821 986
rect 1786 973 1805 976
rect 1786 946 1789 973
rect 1754 943 1789 946
rect 1610 903 1645 906
rect 1602 893 1633 896
rect 1594 803 1597 816
rect 1602 803 1605 866
rect 1618 813 1621 856
rect 1630 836 1633 893
rect 1650 846 1653 926
rect 1642 843 1653 846
rect 1658 843 1661 936
rect 1666 903 1669 936
rect 1674 933 1685 936
rect 1690 933 1709 936
rect 1714 933 1741 936
rect 1674 923 1677 933
rect 1674 896 1677 916
rect 1682 903 1685 926
rect 1690 913 1693 926
rect 1674 893 1685 896
rect 1630 833 1637 836
rect 1618 796 1621 806
rect 1626 803 1629 816
rect 1634 806 1637 833
rect 1642 813 1645 843
rect 1654 833 1677 836
rect 1634 803 1645 806
rect 1562 793 1645 796
rect 1546 763 1589 766
rect 1522 693 1525 726
rect 1530 696 1533 736
rect 1546 733 1549 763
rect 1562 723 1565 736
rect 1586 723 1589 763
rect 1642 723 1645 793
rect 1654 766 1657 833
rect 1666 813 1669 826
rect 1674 813 1677 833
rect 1682 813 1685 893
rect 1698 846 1701 926
rect 1714 916 1717 933
rect 1722 923 1733 926
rect 1706 913 1717 916
rect 1706 903 1717 906
rect 1722 903 1725 916
rect 1714 893 1717 903
rect 1730 866 1733 923
rect 1738 913 1741 933
rect 1746 873 1749 936
rect 1754 923 1757 943
rect 1730 863 1749 866
rect 1694 843 1701 846
rect 1674 803 1685 806
rect 1694 796 1697 843
rect 1706 823 1709 836
rect 1714 813 1733 816
rect 1738 813 1741 826
rect 1714 803 1717 813
rect 1650 763 1657 766
rect 1682 793 1697 796
rect 1546 703 1549 716
rect 1650 706 1653 763
rect 1658 713 1661 746
rect 1650 703 1661 706
rect 1530 693 1549 696
rect 1530 593 1533 686
rect 1522 513 1525 576
rect 1538 526 1541 656
rect 1546 533 1549 693
rect 1554 543 1557 696
rect 1562 563 1565 676
rect 1578 653 1645 656
rect 1578 603 1581 653
rect 1610 623 1613 636
rect 1594 603 1605 606
rect 1570 583 1573 596
rect 1562 543 1597 546
rect 1554 526 1557 536
rect 1538 523 1557 526
rect 1562 523 1565 543
rect 1570 523 1573 536
rect 1482 483 1493 486
rect 1466 453 1473 456
rect 1466 436 1469 453
rect 1450 423 1453 436
rect 1458 433 1469 436
rect 1426 383 1429 406
rect 1438 403 1445 406
rect 1370 333 1373 346
rect 1378 333 1381 366
rect 1330 313 1349 316
rect 1354 313 1357 326
rect 1362 323 1381 326
rect 1386 306 1389 326
rect 1378 303 1389 306
rect 1378 246 1381 303
rect 1378 243 1389 246
rect 1258 213 1261 233
rect 1274 226 1277 233
rect 1266 213 1269 226
rect 1274 223 1293 226
rect 1322 216 1325 226
rect 1330 223 1333 236
rect 1386 223 1389 243
rect 1394 216 1397 356
rect 1438 346 1441 403
rect 1450 353 1453 416
rect 1458 403 1461 433
rect 1402 323 1405 336
rect 1426 333 1429 346
rect 1434 343 1441 346
rect 1402 296 1405 316
rect 1418 303 1421 326
rect 1426 296 1429 326
rect 1402 293 1429 296
rect 1274 203 1277 216
rect 1298 203 1301 216
rect 1314 213 1333 216
rect 1362 213 1397 216
rect 1314 203 1333 206
rect 1362 203 1365 213
rect 1378 203 1381 213
rect 1242 173 1249 176
rect 1226 143 1237 146
rect 1234 123 1237 143
rect 1246 96 1249 173
rect 1266 123 1269 136
rect 1314 123 1317 203
rect 1346 123 1349 156
rect 1362 123 1365 186
rect 1386 123 1389 206
rect 1394 193 1397 206
rect 1410 203 1413 256
rect 1434 243 1437 343
rect 1442 333 1453 336
rect 1466 326 1469 426
rect 1474 403 1477 426
rect 1482 333 1485 416
rect 1450 313 1453 326
rect 1418 213 1421 226
rect 1450 223 1453 306
rect 1458 296 1461 326
rect 1466 323 1477 326
rect 1474 313 1477 323
rect 1458 293 1469 296
rect 1482 263 1485 326
rect 1490 223 1493 483
rect 1554 476 1557 523
rect 1578 513 1581 536
rect 1594 533 1597 543
rect 1554 473 1565 476
rect 1498 423 1525 426
rect 1498 403 1501 416
rect 1506 383 1509 416
rect 1522 413 1525 423
rect 1514 373 1517 406
rect 1498 333 1509 336
rect 1506 293 1509 316
rect 1522 256 1525 406
rect 1530 403 1533 446
rect 1554 413 1557 466
rect 1546 323 1549 336
rect 1514 253 1525 256
rect 1434 193 1445 196
rect 1442 123 1445 193
rect 1450 176 1453 206
rect 1466 183 1469 206
rect 1490 176 1493 216
rect 1514 193 1517 253
rect 1554 213 1557 406
rect 1562 373 1565 473
rect 1586 453 1589 526
rect 1602 506 1605 526
rect 1598 503 1605 506
rect 1610 503 1613 546
rect 1618 536 1621 586
rect 1626 543 1629 636
rect 1634 623 1637 646
rect 1642 633 1645 653
rect 1642 603 1645 626
rect 1650 613 1653 636
rect 1658 603 1661 703
rect 1666 693 1669 726
rect 1682 713 1685 793
rect 1714 783 1717 796
rect 1722 753 1725 806
rect 1738 773 1741 806
rect 1746 793 1749 863
rect 1690 743 1741 746
rect 1690 706 1693 736
rect 1698 723 1709 726
rect 1714 716 1717 736
rect 1674 703 1693 706
rect 1706 713 1717 716
rect 1706 656 1709 713
rect 1722 693 1725 716
rect 1738 713 1741 743
rect 1754 726 1757 866
rect 1762 783 1765 936
rect 1770 903 1773 926
rect 1778 893 1781 936
rect 1786 933 1789 943
rect 1786 913 1789 926
rect 1794 906 1797 966
rect 1802 923 1805 973
rect 1810 963 1813 983
rect 1810 933 1813 956
rect 1818 936 1821 976
rect 1830 966 1833 1043
rect 1842 1013 1845 1036
rect 1850 1016 1853 1113
rect 1922 1063 1925 1193
rect 1850 1013 1869 1016
rect 1850 1006 1853 1013
rect 1882 1006 1885 1036
rect 1890 1013 1917 1016
rect 1842 1003 1853 1006
rect 1826 963 1833 966
rect 1826 943 1829 963
rect 1818 933 1829 936
rect 1842 933 1845 966
rect 1850 933 1853 956
rect 1826 922 1837 925
rect 1826 916 1829 922
rect 1786 903 1797 906
rect 1802 913 1829 916
rect 1770 843 1773 876
rect 1750 723 1757 726
rect 1770 723 1773 816
rect 1786 813 1789 903
rect 1802 883 1805 913
rect 1794 813 1797 826
rect 1810 813 1813 846
rect 1818 813 1821 886
rect 1826 813 1829 826
rect 1834 806 1837 916
rect 1786 786 1789 806
rect 1778 783 1789 786
rect 1778 763 1781 783
rect 1730 656 1733 706
rect 1750 676 1753 723
rect 1778 716 1781 746
rect 1750 673 1757 676
rect 1666 583 1669 626
rect 1674 553 1677 626
rect 1682 603 1685 616
rect 1690 546 1693 636
rect 1698 623 1701 656
rect 1706 653 1717 656
rect 1634 536 1637 546
rect 1666 543 1693 546
rect 1698 536 1701 596
rect 1706 593 1709 646
rect 1714 603 1717 653
rect 1722 613 1725 656
rect 1730 653 1749 656
rect 1754 653 1757 673
rect 1746 636 1749 653
rect 1762 643 1765 716
rect 1770 713 1781 716
rect 1786 713 1789 776
rect 1770 696 1773 713
rect 1794 706 1797 786
rect 1802 743 1805 806
rect 1818 783 1821 806
rect 1826 803 1837 806
rect 1842 796 1845 926
rect 1850 903 1853 926
rect 1858 923 1861 1006
rect 1882 1003 1909 1006
rect 1914 996 1917 1006
rect 1890 993 1917 996
rect 1890 946 1893 993
rect 1882 943 1893 946
rect 1866 913 1869 936
rect 1874 883 1877 926
rect 1882 873 1885 943
rect 1890 933 1901 936
rect 1914 933 1917 986
rect 1922 966 1925 1046
rect 1930 1016 1933 1256
rect 1938 1023 1941 1226
rect 1954 1086 1957 1226
rect 1962 1213 1965 1306
rect 1974 1246 1977 1313
rect 1974 1243 1981 1246
rect 1970 1213 1973 1226
rect 1962 1183 1965 1206
rect 1978 1173 1981 1243
rect 1986 1203 1989 1416
rect 2034 1366 2037 1423
rect 1994 1203 1997 1366
rect 2034 1363 2045 1366
rect 2050 1363 2053 1416
rect 2026 1336 2029 1346
rect 2002 1333 2029 1336
rect 1962 1153 1973 1156
rect 1970 1123 1973 1153
rect 1946 1083 1957 1086
rect 1930 1013 1941 1016
rect 1922 963 1933 966
rect 1938 963 1941 1013
rect 1930 943 1933 963
rect 1890 903 1893 926
rect 1938 913 1941 926
rect 1850 803 1853 826
rect 1866 816 1869 856
rect 1874 823 1877 836
rect 1842 793 1853 796
rect 1858 793 1861 816
rect 1866 813 1877 816
rect 1834 733 1845 736
rect 1850 726 1853 793
rect 1778 703 1797 706
rect 1802 706 1805 726
rect 1834 723 1853 726
rect 1802 703 1813 706
rect 1770 693 1801 696
rect 1770 636 1773 686
rect 1746 633 1757 636
rect 1738 623 1749 626
rect 1754 616 1757 633
rect 1722 593 1725 606
rect 1730 573 1733 616
rect 1746 613 1757 616
rect 1762 633 1773 636
rect 1762 613 1765 633
rect 1778 613 1781 626
rect 1786 613 1789 676
rect 1798 626 1801 693
rect 1810 683 1813 703
rect 1818 663 1821 716
rect 1834 703 1837 723
rect 1798 623 1805 626
rect 1618 533 1629 536
rect 1618 523 1621 533
rect 1626 523 1629 533
rect 1634 533 1677 536
rect 1682 533 1701 536
rect 1714 536 1717 556
rect 1738 543 1741 586
rect 1714 533 1725 536
rect 1570 413 1573 436
rect 1578 403 1581 446
rect 1598 426 1601 503
rect 1598 423 1605 426
rect 1586 353 1589 416
rect 1602 403 1605 423
rect 1594 346 1597 396
rect 1594 343 1605 346
rect 1562 213 1565 336
rect 1602 323 1605 343
rect 1610 293 1613 466
rect 1618 403 1621 446
rect 1634 423 1637 533
rect 1682 526 1685 533
rect 1746 526 1749 613
rect 1802 606 1805 623
rect 1810 613 1813 636
rect 1754 603 1765 606
rect 1786 593 1789 606
rect 1794 586 1797 606
rect 1802 603 1813 606
rect 1810 593 1813 603
rect 1818 586 1821 616
rect 1826 603 1829 646
rect 1842 603 1845 716
rect 1858 653 1861 776
rect 1874 736 1877 813
rect 1882 803 1885 846
rect 1922 826 1925 846
rect 1890 823 1925 826
rect 1930 823 1933 896
rect 1946 863 1949 1083
rect 1954 963 1957 1066
rect 1986 1036 1989 1196
rect 2002 1123 2005 1333
rect 2034 1303 2037 1336
rect 2010 1176 2013 1246
rect 2026 1213 2029 1236
rect 2042 1213 2045 1363
rect 2058 1343 2061 1416
rect 2074 1366 2077 1423
rect 2066 1363 2077 1366
rect 2050 1323 2053 1336
rect 2058 1303 2061 1336
rect 2066 1296 2069 1363
rect 2058 1293 2069 1296
rect 2058 1226 2061 1293
rect 2074 1253 2077 1346
rect 2066 1233 2085 1236
rect 2018 1196 2021 1206
rect 2050 1196 2053 1226
rect 2058 1223 2077 1226
rect 2018 1193 2053 1196
rect 2010 1173 2021 1176
rect 2018 1116 2021 1173
rect 2058 1143 2061 1216
rect 2082 1183 2085 1233
rect 2090 1213 2093 1226
rect 2098 1213 2101 1436
rect 2114 1426 2117 1496
rect 2110 1423 2117 1426
rect 2110 1356 2113 1423
rect 2130 1416 2133 1503
rect 2162 1496 2165 1626
rect 2170 1503 2173 1606
rect 2178 1576 2181 1763
rect 2202 1636 2205 1726
rect 2218 1723 2221 1773
rect 2202 1633 2229 1636
rect 2178 1573 2189 1576
rect 2186 1516 2189 1573
rect 2226 1523 2229 1633
rect 2234 1583 2237 1806
rect 2258 1746 2261 1806
rect 2258 1743 2265 1746
rect 2262 1696 2265 1743
rect 2258 1693 2265 1696
rect 2242 1603 2245 1626
rect 2258 1603 2261 1693
rect 2266 1613 2269 1626
rect 2178 1513 2189 1516
rect 2154 1493 2165 1496
rect 2178 1493 2181 1513
rect 2154 1436 2157 1493
rect 2154 1433 2165 1436
rect 2130 1413 2157 1416
rect 2122 1373 2125 1406
rect 2110 1353 2117 1356
rect 2114 1333 2117 1353
rect 2154 1333 2157 1413
rect 2162 1376 2165 1433
rect 2178 1403 2181 1486
rect 2242 1456 2245 1526
rect 2266 1506 2269 1526
rect 2262 1503 2269 1506
rect 2226 1453 2245 1456
rect 2226 1413 2229 1453
rect 2162 1373 2169 1376
rect 2166 1326 2169 1373
rect 2162 1323 2169 1326
rect 2106 1213 2109 1236
rect 2098 1203 2109 1206
rect 2114 1203 2117 1246
rect 2122 1203 2125 1226
rect 2146 1223 2149 1236
rect 2162 1216 2165 1323
rect 2178 1313 2181 1326
rect 2170 1223 2173 1246
rect 2210 1223 2213 1326
rect 2234 1313 2237 1336
rect 2250 1293 2253 1466
rect 2262 1436 2265 1503
rect 2274 1463 2277 1943
rect 2282 1913 2285 1926
rect 2290 1923 2293 1963
rect 2330 1903 2333 1926
rect 2282 1813 2285 1836
rect 2314 1813 2317 1826
rect 2322 1813 2325 1836
rect 2330 1823 2357 1826
rect 2330 1806 2333 1823
rect 2338 1813 2349 1816
rect 2354 1813 2357 1823
rect 2322 1803 2333 1806
rect 2322 1733 2333 1736
rect 2346 1733 2349 1806
rect 2362 1733 2365 1926
rect 2426 1923 2429 1936
rect 2434 1923 2437 2023
rect 2442 2003 2445 2016
rect 2370 1813 2373 1826
rect 2386 1813 2389 1836
rect 2410 1776 2413 1826
rect 2442 1813 2445 1826
rect 2458 1813 2461 1916
rect 2514 1896 2517 2006
rect 2530 2003 2533 2223
rect 2538 2203 2541 2216
rect 2546 2193 2549 2336
rect 2554 2333 2557 2343
rect 2554 2313 2557 2326
rect 2562 2236 2565 2373
rect 2586 2333 2589 2373
rect 2570 2286 2573 2326
rect 2610 2286 2613 2326
rect 2666 2313 2669 2326
rect 2570 2283 2613 2286
rect 2618 2253 2661 2256
rect 2562 2233 2573 2236
rect 2554 2213 2557 2226
rect 2570 2126 2573 2233
rect 2618 2213 2621 2253
rect 2650 2213 2653 2226
rect 2658 2213 2661 2253
rect 2650 2203 2661 2206
rect 2570 2123 2589 2126
rect 2538 1993 2541 2016
rect 2546 2013 2557 2016
rect 2570 2013 2573 2026
rect 2546 1936 2549 2006
rect 2554 1993 2557 2006
rect 2586 1986 2589 2123
rect 2610 2013 2613 2026
rect 2658 2013 2669 2016
rect 2522 1933 2549 1936
rect 2570 1983 2589 1986
rect 2522 1903 2525 1926
rect 2530 1923 2541 1926
rect 2546 1903 2549 1926
rect 2554 1913 2557 1926
rect 2514 1893 2533 1896
rect 2482 1823 2485 1836
rect 2458 1803 2469 1806
rect 2386 1773 2413 1776
rect 2282 1703 2285 1726
rect 2314 1713 2317 1726
rect 2322 1703 2325 1726
rect 2330 1686 2333 1733
rect 2338 1723 2349 1726
rect 2354 1686 2357 1726
rect 2370 1713 2373 1726
rect 2386 1723 2389 1773
rect 2410 1703 2413 1716
rect 2442 1713 2445 1726
rect 2450 1703 2453 1726
rect 2458 1713 2461 1736
rect 2330 1683 2357 1686
rect 2290 1623 2301 1626
rect 2298 1613 2301 1623
rect 2282 1533 2285 1586
rect 2482 1583 2485 1716
rect 2530 1606 2533 1893
rect 2554 1813 2557 1876
rect 2570 1856 2573 1983
rect 2658 1933 2669 1936
rect 2594 1913 2597 1926
rect 2642 1923 2653 1926
rect 2658 1856 2661 1926
rect 2666 1873 2669 1933
rect 2570 1853 2589 1856
rect 2554 1613 2557 1726
rect 2562 1696 2565 1806
rect 2570 1803 2573 1816
rect 2586 1733 2589 1853
rect 2634 1853 2661 1856
rect 2634 1813 2637 1853
rect 2666 1803 2669 1816
rect 2570 1713 2573 1726
rect 2562 1693 2573 1696
rect 2514 1603 2533 1606
rect 2306 1543 2325 1546
rect 2290 1503 2293 1526
rect 2298 1463 2301 1536
rect 2306 1523 2309 1543
rect 2262 1433 2269 1436
rect 2258 1403 2261 1416
rect 2266 1343 2269 1433
rect 2314 1406 2317 1536
rect 2322 1533 2325 1543
rect 2482 1536 2485 1556
rect 2322 1513 2325 1526
rect 2330 1413 2333 1526
rect 2346 1516 2349 1536
rect 2426 1533 2437 1536
rect 2474 1533 2485 1536
rect 2338 1513 2349 1516
rect 2354 1513 2357 1526
rect 2346 1416 2349 1513
rect 2370 1426 2373 1516
rect 2410 1503 2413 1516
rect 2434 1503 2437 1526
rect 2442 1513 2453 1516
rect 2474 1466 2477 1533
rect 2474 1463 2485 1466
rect 2482 1446 2485 1463
rect 2482 1443 2489 1446
rect 2370 1423 2377 1426
rect 2346 1413 2365 1416
rect 2282 1356 2285 1406
rect 2314 1403 2333 1406
rect 2274 1353 2285 1356
rect 2266 1313 2269 1336
rect 2274 1296 2277 1353
rect 2282 1343 2317 1346
rect 2282 1323 2285 1343
rect 2290 1306 2293 1326
rect 2298 1316 2301 1336
rect 2314 1333 2317 1343
rect 2330 1336 2333 1403
rect 2374 1376 2377 1423
rect 2466 1413 2469 1426
rect 2418 1393 2421 1406
rect 2486 1376 2489 1443
rect 2498 1413 2501 1536
rect 2506 1413 2509 1426
rect 2506 1393 2509 1406
rect 2374 1373 2381 1376
rect 2330 1333 2341 1336
rect 2314 1323 2325 1326
rect 2330 1316 2333 1326
rect 2298 1313 2333 1316
rect 2290 1303 2317 1306
rect 2274 1293 2293 1296
rect 2218 1223 2221 1236
rect 2130 1213 2149 1216
rect 2162 1213 2173 1216
rect 2010 1113 2021 1116
rect 1986 1033 1993 1036
rect 1970 1003 1973 1016
rect 1978 1013 1981 1026
rect 1954 893 1957 946
rect 1890 813 1893 823
rect 1882 743 1893 746
rect 1866 693 1869 736
rect 1874 733 1885 736
rect 1866 593 1869 616
rect 1794 583 1821 586
rect 1754 533 1765 536
rect 1674 523 1685 526
rect 1690 516 1693 526
rect 1698 523 1717 526
rect 1690 513 1709 516
rect 1714 503 1717 523
rect 1722 523 1749 526
rect 1642 423 1645 436
rect 1650 433 1653 446
rect 1682 433 1685 456
rect 1650 416 1653 426
rect 1626 413 1653 416
rect 1586 243 1613 246
rect 1618 243 1621 346
rect 1586 213 1589 243
rect 1602 213 1605 236
rect 1610 226 1613 243
rect 1610 223 1621 226
rect 1578 183 1581 206
rect 1450 173 1493 176
rect 1562 133 1565 146
rect 1594 123 1597 206
rect 1610 173 1613 216
rect 1618 213 1621 223
rect 1626 216 1629 413
rect 1642 373 1645 406
rect 1658 363 1661 416
rect 1690 366 1693 416
rect 1706 406 1709 426
rect 1706 403 1717 406
rect 1722 403 1725 523
rect 1754 516 1757 526
rect 1730 513 1757 516
rect 1762 503 1765 533
rect 1770 523 1781 526
rect 1770 476 1773 516
rect 1778 483 1781 523
rect 1786 513 1789 576
rect 1874 573 1877 726
rect 1794 543 1805 546
rect 1794 476 1797 536
rect 1802 503 1805 543
rect 1826 543 1869 546
rect 1826 533 1829 543
rect 1826 503 1829 526
rect 1834 523 1837 536
rect 1842 533 1861 536
rect 1866 533 1869 543
rect 1858 526 1861 533
rect 1882 526 1885 733
rect 1898 723 1901 806
rect 1906 803 1909 816
rect 1914 803 1917 816
rect 1930 783 1933 816
rect 1938 776 1941 836
rect 1906 773 1941 776
rect 1906 676 1909 773
rect 1946 756 1949 826
rect 1954 813 1957 846
rect 1938 753 1949 756
rect 1930 733 1933 746
rect 1914 723 1933 726
rect 1898 673 1909 676
rect 1890 583 1893 666
rect 1770 473 1797 476
rect 1754 433 1789 436
rect 1714 393 1717 403
rect 1738 373 1741 416
rect 1754 403 1757 433
rect 1778 416 1781 426
rect 1786 423 1789 433
rect 1794 423 1805 426
rect 1810 423 1813 496
rect 1690 363 1709 366
rect 1634 323 1637 336
rect 1658 333 1669 336
rect 1642 323 1661 326
rect 1642 316 1645 323
rect 1634 313 1645 316
rect 1634 283 1637 306
rect 1650 303 1653 316
rect 1626 213 1637 216
rect 1642 206 1645 296
rect 1658 293 1661 323
rect 1666 206 1669 333
rect 1674 313 1677 336
rect 1682 323 1685 336
rect 1618 203 1645 206
rect 1642 123 1645 203
rect 1650 203 1669 206
rect 1650 183 1653 203
rect 1674 173 1677 206
rect 1682 203 1685 216
rect 1690 153 1693 336
rect 1698 333 1701 356
rect 1698 293 1701 326
rect 1706 303 1709 363
rect 1698 213 1701 236
rect 1698 203 1709 206
rect 1674 133 1677 146
rect 1698 123 1701 176
rect 1722 143 1725 336
rect 1746 313 1749 326
rect 1762 213 1765 416
rect 1770 413 1781 416
rect 1786 413 1797 416
rect 1770 403 1773 413
rect 1778 363 1781 406
rect 1794 396 1797 413
rect 1802 406 1805 423
rect 1802 403 1813 406
rect 1790 393 1797 396
rect 1790 336 1793 393
rect 1790 333 1797 336
rect 1794 316 1797 333
rect 1802 323 1805 356
rect 1810 333 1813 403
rect 1794 313 1805 316
rect 1810 313 1813 326
rect 1786 223 1789 266
rect 1778 213 1789 216
rect 1754 123 1757 206
rect 1762 203 1773 206
rect 1770 133 1773 196
rect 1778 163 1781 213
rect 1786 183 1789 206
rect 1802 203 1805 313
rect 1818 296 1821 426
rect 1826 316 1829 476
rect 1842 413 1845 526
rect 1858 523 1885 526
rect 1850 406 1853 416
rect 1834 403 1853 406
rect 1858 403 1861 466
rect 1866 413 1869 516
rect 1882 513 1885 523
rect 1890 493 1893 526
rect 1898 503 1901 536
rect 1906 533 1909 673
rect 1914 613 1925 616
rect 1930 613 1933 723
rect 1938 713 1941 753
rect 1946 733 1949 746
rect 1954 723 1957 786
rect 1962 773 1965 956
rect 1978 836 1981 1006
rect 1990 956 1993 1033
rect 2010 1013 2013 1113
rect 2010 996 2013 1006
rect 2018 1003 2021 1026
rect 2050 1013 2053 1036
rect 2002 973 2005 996
rect 2010 993 2037 996
rect 1970 833 1981 836
rect 1986 953 1993 956
rect 1986 833 1989 953
rect 1994 923 1997 936
rect 2002 933 2005 956
rect 1970 753 1973 833
rect 1978 803 1981 826
rect 1986 783 1989 816
rect 1994 746 1997 876
rect 2002 813 2005 846
rect 2010 813 2013 936
rect 2018 933 2021 946
rect 2002 803 2013 806
rect 2018 786 2021 846
rect 2026 793 2029 926
rect 2034 843 2037 976
rect 2042 913 2045 936
rect 2050 923 2053 936
rect 2066 906 2069 1136
rect 2090 1013 2093 1036
rect 2090 923 2093 946
rect 2098 916 2101 1196
rect 2106 1153 2109 1203
rect 2146 1176 2149 1206
rect 2154 1193 2157 1206
rect 2170 1203 2173 1213
rect 2178 1193 2181 1206
rect 2202 1193 2205 1216
rect 2218 1183 2221 1216
rect 2234 1203 2237 1226
rect 2242 1203 2245 1226
rect 2266 1216 2269 1246
rect 2266 1213 2277 1216
rect 2146 1173 2181 1176
rect 2138 1146 2141 1166
rect 2130 1143 2141 1146
rect 2130 1066 2133 1143
rect 2154 1066 2157 1136
rect 2178 1123 2181 1173
rect 2234 1123 2237 1186
rect 2130 1063 2137 1066
rect 2154 1063 2165 1066
rect 2042 903 2069 906
rect 2090 913 2101 916
rect 2014 783 2021 786
rect 1994 743 2005 746
rect 1970 713 1973 736
rect 1994 723 1997 736
rect 2002 696 2005 743
rect 1986 693 2005 696
rect 1946 623 1949 646
rect 1954 616 1957 636
rect 1938 613 1957 616
rect 1938 606 1941 613
rect 1962 606 1965 656
rect 1978 613 1981 646
rect 1930 603 1941 606
rect 1954 603 1965 606
rect 1970 603 1981 606
rect 1930 536 1933 596
rect 1914 526 1917 536
rect 1922 533 1933 536
rect 1954 536 1957 603
rect 1986 583 1989 693
rect 2014 686 2017 783
rect 2042 776 2045 903
rect 2090 856 2093 913
rect 2134 906 2137 1063
rect 2146 933 2149 1026
rect 2162 1003 2165 1063
rect 2242 1026 2245 1196
rect 2266 1183 2269 1206
rect 2250 1116 2253 1146
rect 2274 1126 2277 1213
rect 2258 1123 2277 1126
rect 2250 1113 2261 1116
rect 2186 996 2189 1016
rect 2146 913 2149 926
rect 2134 903 2141 906
rect 2082 853 2093 856
rect 2066 813 2069 826
rect 2038 773 2045 776
rect 2082 776 2085 853
rect 2122 803 2125 816
rect 2082 773 2093 776
rect 2038 706 2041 773
rect 2090 746 2093 773
rect 2130 746 2133 806
rect 2050 723 2053 746
rect 2082 743 2093 746
rect 2114 743 2133 746
rect 2038 703 2045 706
rect 2042 686 2045 703
rect 2014 683 2021 686
rect 2042 683 2053 686
rect 2018 646 2021 683
rect 2002 643 2021 646
rect 1994 613 1997 636
rect 1994 563 1997 606
rect 2002 566 2005 643
rect 2018 576 2021 606
rect 2042 603 2045 616
rect 2050 576 2053 683
rect 2082 666 2085 743
rect 2082 663 2093 666
rect 2090 593 2093 663
rect 2018 573 2053 576
rect 2002 563 2021 566
rect 1954 533 1989 536
rect 1906 496 1909 526
rect 1914 523 1925 526
rect 1930 516 1933 533
rect 1954 523 1965 526
rect 1970 523 1989 526
rect 1926 513 1933 516
rect 1906 493 1917 496
rect 1874 403 1877 416
rect 1834 383 1837 403
rect 1882 373 1885 416
rect 1890 403 1893 466
rect 1898 393 1901 416
rect 1906 403 1909 486
rect 1834 323 1837 336
rect 1826 313 1837 316
rect 1818 293 1829 296
rect 1826 226 1829 293
rect 1850 286 1853 336
rect 1874 323 1877 366
rect 1906 363 1909 396
rect 1914 353 1917 493
rect 1926 446 1929 513
rect 1938 493 1941 516
rect 1946 503 1949 516
rect 1954 473 1957 523
rect 1970 516 1973 523
rect 1962 513 1973 516
rect 1978 513 1997 516
rect 2002 513 2005 536
rect 1922 443 1929 446
rect 1922 403 1925 443
rect 1930 413 1933 426
rect 1962 423 1965 436
rect 1938 413 1965 416
rect 1954 396 1957 406
rect 1922 393 1957 396
rect 1922 363 1925 393
rect 1850 283 1861 286
rect 1818 223 1829 226
rect 1818 203 1821 223
rect 1858 193 1861 283
rect 1882 213 1885 326
rect 1922 256 1925 336
rect 1930 323 1933 386
rect 1922 253 1929 256
rect 1926 196 1929 253
rect 1938 213 1941 376
rect 1946 316 1949 346
rect 1954 333 1957 356
rect 1962 323 1965 413
rect 1970 393 1973 406
rect 1978 346 1981 416
rect 1970 343 1981 346
rect 1970 326 1973 343
rect 1986 336 1989 506
rect 1994 423 1997 513
rect 2010 473 2013 526
rect 2018 453 2021 563
rect 2026 533 2029 546
rect 2026 493 2029 526
rect 1994 403 1997 416
rect 2002 403 2005 426
rect 2010 413 2013 446
rect 2018 393 2021 436
rect 2026 423 2029 436
rect 2050 416 2053 573
rect 2074 513 2077 526
rect 2074 436 2077 456
rect 2042 413 2053 416
rect 2066 433 2077 436
rect 1978 333 1989 336
rect 1994 333 1997 346
rect 1970 323 1981 326
rect 1946 313 1973 316
rect 1978 226 1981 323
rect 1986 303 1989 326
rect 2002 313 2005 326
rect 2010 273 2013 386
rect 2018 313 2021 336
rect 2026 303 2029 366
rect 1962 223 1997 226
rect 1962 213 1965 223
rect 1922 193 1929 196
rect 1802 123 1805 186
rect 1922 173 1925 193
rect 1946 173 1949 206
rect 1842 163 1853 166
rect 1850 123 1853 163
rect 1970 146 1973 206
rect 1978 203 1981 216
rect 1986 203 1989 216
rect 1994 213 1997 223
rect 1994 166 1997 206
rect 1994 163 2037 166
rect 1954 133 1957 146
rect 1970 143 1981 146
rect 1978 123 1981 143
rect 2034 123 2037 163
rect 2042 143 2045 413
rect 2066 366 2069 433
rect 2082 383 2085 586
rect 2098 563 2101 616
rect 2106 613 2109 736
rect 2114 613 2117 626
rect 2106 593 2109 606
rect 2122 533 2125 743
rect 2130 633 2133 646
rect 2130 613 2133 626
rect 2130 523 2133 546
rect 2138 463 2141 903
rect 2146 723 2149 826
rect 2154 813 2157 946
rect 2162 933 2165 996
rect 2186 993 2197 996
rect 2170 823 2173 966
rect 2194 946 2197 993
rect 2234 966 2237 1026
rect 2242 1023 2253 1026
rect 2186 943 2197 946
rect 2218 963 2237 966
rect 2178 816 2181 846
rect 2162 803 2165 816
rect 2170 813 2181 816
rect 2186 803 2189 943
rect 2194 906 2197 926
rect 2194 903 2205 906
rect 2202 846 2205 903
rect 2194 843 2205 846
rect 2218 846 2221 963
rect 2242 926 2245 1016
rect 2234 923 2245 926
rect 2234 866 2237 923
rect 2234 863 2245 866
rect 2218 843 2237 846
rect 2194 803 2197 843
rect 2210 796 2213 826
rect 2178 793 2213 796
rect 2162 693 2165 736
rect 2170 716 2173 726
rect 2178 723 2181 793
rect 2186 733 2197 736
rect 2210 733 2213 746
rect 2186 716 2189 726
rect 2170 713 2189 716
rect 2146 633 2165 636
rect 2154 583 2157 626
rect 2162 456 2165 633
rect 2178 613 2181 626
rect 2186 613 2189 646
rect 2194 633 2197 733
rect 2218 713 2221 736
rect 2226 706 2229 816
rect 2234 806 2237 843
rect 2242 823 2245 863
rect 2250 813 2253 1023
rect 2258 926 2261 1113
rect 2266 1103 2269 1116
rect 2290 1106 2293 1293
rect 2314 1213 2317 1303
rect 2370 1213 2373 1326
rect 2378 1323 2381 1373
rect 2482 1373 2489 1376
rect 2442 1333 2445 1346
rect 2394 1246 2397 1316
rect 2434 1313 2437 1326
rect 2386 1243 2397 1246
rect 2378 1203 2381 1226
rect 2386 1213 2389 1243
rect 2410 1223 2413 1236
rect 2450 1206 2453 1296
rect 2450 1203 2461 1206
rect 2474 1196 2477 1216
rect 2306 1113 2309 1196
rect 2450 1193 2477 1196
rect 2482 1193 2485 1373
rect 2514 1333 2517 1603
rect 2570 1586 2573 1693
rect 2610 1613 2613 1726
rect 2666 1713 2669 1726
rect 2530 1533 2533 1556
rect 2522 1506 2525 1526
rect 2538 1523 2541 1536
rect 2546 1513 2549 1536
rect 2554 1523 2557 1586
rect 2562 1583 2573 1586
rect 2562 1563 2565 1583
rect 2618 1533 2621 1546
rect 2650 1533 2653 1556
rect 2522 1503 2533 1506
rect 2570 1503 2573 1516
rect 2530 1446 2533 1503
rect 2522 1443 2533 1446
rect 2522 1393 2525 1443
rect 2586 1413 2589 1426
rect 2618 1413 2621 1516
rect 2626 1413 2629 1426
rect 2642 1406 2645 1526
rect 2658 1513 2661 1526
rect 2538 1383 2541 1406
rect 2626 1403 2645 1406
rect 2522 1343 2541 1346
rect 2506 1243 2509 1326
rect 2522 1323 2525 1343
rect 2530 1323 2533 1336
rect 2538 1333 2541 1343
rect 2586 1333 2589 1386
rect 2538 1236 2541 1326
rect 2570 1286 2573 1326
rect 2610 1286 2613 1326
rect 2666 1313 2669 1326
rect 2570 1283 2613 1286
rect 2490 1213 2493 1226
rect 2498 1213 2501 1236
rect 2506 1233 2541 1236
rect 2506 1206 2509 1233
rect 2530 1213 2533 1226
rect 2498 1203 2509 1206
rect 2290 1103 2297 1106
rect 2282 1013 2285 1096
rect 2294 1056 2297 1103
rect 2314 1076 2317 1186
rect 2322 1086 2325 1126
rect 2338 1093 2341 1136
rect 2450 1133 2453 1193
rect 2474 1133 2477 1176
rect 2362 1086 2365 1126
rect 2322 1083 2365 1086
rect 2314 1073 2325 1076
rect 2294 1053 2301 1056
rect 2298 1006 2301 1053
rect 2290 1003 2301 1006
rect 2266 943 2285 946
rect 2258 923 2265 926
rect 2234 803 2253 806
rect 2234 713 2237 796
rect 2226 703 2245 706
rect 2210 633 2229 636
rect 2210 626 2213 633
rect 2194 623 2213 626
rect 2178 546 2181 606
rect 2194 603 2197 623
rect 2202 613 2213 616
rect 2218 613 2221 626
rect 2234 623 2237 646
rect 2234 583 2237 616
rect 2242 606 2245 703
rect 2250 653 2253 803
rect 2262 786 2265 923
rect 2274 813 2277 926
rect 2282 833 2285 936
rect 2290 916 2293 1003
rect 2322 963 2325 1073
rect 2418 1066 2421 1126
rect 2458 1086 2461 1126
rect 2498 1086 2501 1126
rect 2554 1123 2557 1226
rect 2562 1223 2565 1246
rect 2610 1233 2653 1236
rect 2578 1213 2581 1226
rect 2562 1203 2573 1206
rect 2594 1183 2597 1216
rect 2602 1193 2605 1206
rect 2610 1186 2613 1233
rect 2618 1203 2621 1216
rect 2642 1213 2645 1226
rect 2650 1213 2653 1233
rect 2610 1183 2653 1186
rect 2570 1133 2573 1176
rect 2458 1083 2501 1086
rect 2618 1086 2621 1126
rect 2650 1123 2653 1183
rect 2658 1133 2661 1186
rect 2658 1086 2661 1126
rect 2618 1083 2661 1086
rect 2418 1063 2429 1066
rect 2426 1033 2429 1063
rect 2442 983 2445 1026
rect 2298 933 2301 946
rect 2314 916 2317 926
rect 2322 923 2325 946
rect 2362 943 2365 966
rect 2394 943 2397 956
rect 2330 923 2333 936
rect 2338 933 2357 936
rect 2338 916 2341 933
rect 2290 913 2301 916
rect 2314 913 2341 916
rect 2298 826 2301 913
rect 2354 906 2357 926
rect 2370 913 2373 926
rect 2322 903 2357 906
rect 2290 823 2301 826
rect 2314 823 2317 836
rect 2258 783 2265 786
rect 2258 763 2261 783
rect 2290 766 2293 823
rect 2322 813 2325 903
rect 2346 806 2349 816
rect 2322 793 2325 806
rect 2338 803 2349 806
rect 2290 763 2301 766
rect 2290 723 2293 746
rect 2250 623 2253 636
rect 2242 603 2249 606
rect 2178 543 2197 546
rect 2162 453 2169 456
rect 2098 366 2101 406
rect 2138 366 2141 396
rect 2066 363 2077 366
rect 2066 323 2069 346
rect 2074 316 2077 363
rect 2066 313 2077 316
rect 2086 363 2141 366
rect 2146 366 2149 416
rect 2166 376 2169 453
rect 2178 413 2181 536
rect 2194 466 2197 543
rect 2246 536 2249 603
rect 2258 543 2261 626
rect 2266 623 2269 636
rect 2274 616 2277 646
rect 2290 636 2293 696
rect 2282 633 2293 636
rect 2282 623 2285 633
rect 2266 613 2277 616
rect 2290 546 2293 586
rect 2298 576 2301 763
rect 2322 583 2325 766
rect 2330 713 2333 726
rect 2338 613 2341 803
rect 2354 796 2357 836
rect 2362 813 2365 846
rect 2378 803 2381 816
rect 2394 806 2397 926
rect 2402 923 2405 936
rect 2410 933 2413 946
rect 2418 836 2421 926
rect 2426 923 2429 936
rect 2450 926 2453 1016
rect 2466 1006 2469 1026
rect 2474 1013 2485 1016
rect 2466 1003 2477 1006
rect 2498 963 2501 1016
rect 2466 933 2485 936
rect 2490 933 2493 956
rect 2482 926 2485 933
rect 2434 913 2437 926
rect 2450 923 2461 926
rect 2390 803 2397 806
rect 2402 833 2421 836
rect 2346 743 2349 796
rect 2354 793 2381 796
rect 2362 656 2365 736
rect 2378 733 2381 793
rect 2390 746 2393 803
rect 2402 776 2405 833
rect 2410 813 2413 826
rect 2418 813 2421 826
rect 2426 816 2429 836
rect 2434 823 2437 846
rect 2426 813 2445 816
rect 2458 813 2461 923
rect 2474 913 2477 926
rect 2482 923 2501 926
rect 2490 843 2493 916
rect 2442 803 2453 806
rect 2402 773 2437 776
rect 2386 743 2393 746
rect 2402 743 2405 766
rect 2386 723 2389 743
rect 2402 723 2405 736
rect 2362 653 2369 656
rect 2366 576 2369 653
rect 2298 573 2341 576
rect 2266 536 2269 546
rect 2290 543 2301 546
rect 2246 533 2277 536
rect 2186 463 2197 466
rect 2274 466 2277 533
rect 2274 463 2285 466
rect 2166 373 2173 376
rect 2146 363 2165 366
rect 2066 213 2069 313
rect 2086 306 2089 363
rect 2138 333 2141 363
rect 2122 313 2125 326
rect 2082 303 2089 306
rect 2082 203 2085 303
rect 2162 273 2165 363
rect 2130 213 2133 236
rect 2170 213 2173 373
rect 2186 366 2189 463
rect 2202 393 2205 406
rect 2250 393 2253 416
rect 2186 363 2221 366
rect 2186 323 2189 346
rect 2218 323 2221 363
rect 2274 333 2277 416
rect 2282 413 2285 463
rect 2298 436 2301 543
rect 2338 533 2341 573
rect 2362 573 2369 576
rect 2290 433 2301 436
rect 2290 403 2293 433
rect 2314 373 2317 416
rect 2298 333 2301 346
rect 2202 213 2205 226
rect 2210 193 2213 206
rect 2234 203 2237 236
rect 2242 203 2245 306
rect 2250 296 2253 326
rect 2258 303 2261 316
rect 2266 313 2269 326
rect 2250 293 2269 296
rect 2258 226 2261 236
rect 2250 223 2261 226
rect 2258 213 2261 223
rect 2266 216 2269 293
rect 2266 213 2277 216
rect 2282 193 2285 326
rect 2290 323 2301 326
rect 2298 313 2301 323
rect 2322 296 2325 526
rect 2362 523 2365 573
rect 2378 446 2381 616
rect 2426 613 2429 736
rect 2434 723 2437 773
rect 2450 703 2453 726
rect 2458 713 2461 736
rect 2466 723 2469 816
rect 2482 793 2485 806
rect 2490 786 2493 816
rect 2498 793 2501 923
rect 2506 916 2509 946
rect 2522 923 2525 996
rect 2530 923 2533 986
rect 2562 943 2565 1026
rect 2578 1003 2581 1016
rect 2618 1013 2621 1026
rect 2546 916 2549 936
rect 2506 913 2533 916
rect 2538 913 2557 916
rect 2562 913 2565 926
rect 2538 906 2541 913
rect 2554 906 2557 913
rect 2514 903 2541 906
rect 2514 813 2517 903
rect 2522 833 2533 836
rect 2530 803 2533 826
rect 2538 803 2541 816
rect 2546 813 2549 906
rect 2554 903 2561 906
rect 2558 836 2561 903
rect 2558 833 2565 836
rect 2562 813 2565 833
rect 2482 783 2493 786
rect 2474 743 2477 766
rect 2482 733 2485 783
rect 2530 733 2533 746
rect 2546 733 2549 746
rect 2554 736 2557 806
rect 2562 743 2565 796
rect 2570 756 2573 936
rect 2586 933 2589 996
rect 2594 953 2597 1006
rect 2602 963 2621 966
rect 2594 933 2597 946
rect 2578 916 2581 926
rect 2602 923 2605 963
rect 2610 933 2613 956
rect 2618 933 2621 963
rect 2618 916 2621 926
rect 2626 923 2629 936
rect 2578 913 2621 916
rect 2578 896 2581 913
rect 2578 893 2585 896
rect 2582 816 2585 893
rect 2578 813 2585 816
rect 2594 833 2613 836
rect 2578 766 2581 813
rect 2594 803 2597 833
rect 2586 793 2597 796
rect 2578 763 2589 766
rect 2570 753 2581 756
rect 2554 733 2565 736
rect 2570 733 2573 746
rect 2474 656 2477 726
rect 2482 713 2485 726
rect 2522 723 2533 726
rect 2546 703 2549 726
rect 2562 716 2565 733
rect 2578 723 2581 753
rect 2586 726 2589 763
rect 2594 733 2597 746
rect 2602 726 2605 816
rect 2610 743 2613 826
rect 2618 736 2621 816
rect 2634 813 2637 826
rect 2642 803 2645 836
rect 2650 796 2653 946
rect 2618 733 2629 736
rect 2586 723 2605 726
rect 2610 723 2621 726
rect 2586 716 2589 723
rect 2626 716 2629 726
rect 2562 713 2589 716
rect 2594 713 2629 716
rect 2438 653 2477 656
rect 2438 606 2441 653
rect 2394 573 2397 606
rect 2434 603 2441 606
rect 2434 553 2437 603
rect 2442 533 2445 576
rect 2474 566 2477 626
rect 2474 563 2481 566
rect 2354 443 2381 446
rect 2354 413 2357 443
rect 2362 426 2365 436
rect 2370 433 2389 436
rect 2362 423 2381 426
rect 2386 416 2389 433
rect 2330 393 2333 406
rect 2362 386 2365 416
rect 2346 383 2365 386
rect 2378 413 2389 416
rect 2426 416 2429 526
rect 2466 523 2469 556
rect 2478 496 2481 563
rect 2474 493 2481 496
rect 2474 476 2477 493
rect 2466 473 2477 476
rect 2426 413 2453 416
rect 2330 323 2333 336
rect 2322 293 2333 296
rect 2306 213 2309 236
rect 2346 223 2349 383
rect 2362 333 2365 376
rect 2370 343 2373 356
rect 2362 303 2365 316
rect 2370 313 2373 336
rect 2378 326 2381 413
rect 2386 403 2389 413
rect 2434 386 2437 396
rect 2466 386 2469 473
rect 2434 383 2469 386
rect 2378 323 2389 326
rect 2394 323 2397 336
rect 2290 183 2293 206
rect 2314 203 2317 216
rect 2322 193 2325 216
rect 2354 203 2357 276
rect 2378 203 2381 246
rect 2426 233 2429 356
rect 2442 303 2445 326
rect 2394 213 2397 226
rect 2338 183 2341 196
rect 2410 183 2413 226
rect 2434 206 2437 226
rect 2450 213 2453 346
rect 2458 303 2461 383
rect 2466 313 2469 336
rect 2474 313 2477 416
rect 2434 203 2445 206
rect 2458 203 2461 216
rect 2466 183 2469 216
rect 2474 203 2477 306
rect 2482 276 2485 406
rect 2490 383 2493 656
rect 2562 646 2565 713
rect 2634 656 2637 796
rect 2642 793 2653 796
rect 2642 743 2645 793
rect 2658 726 2661 816
rect 2650 723 2661 726
rect 2650 666 2653 723
rect 2650 663 2661 666
rect 2626 653 2637 656
rect 2562 643 2573 646
rect 2514 603 2517 616
rect 2570 613 2573 643
rect 2610 613 2613 626
rect 2538 533 2541 546
rect 2586 543 2589 606
rect 2626 576 2629 653
rect 2658 606 2661 663
rect 2666 613 2669 746
rect 2658 603 2669 606
rect 2626 573 2637 576
rect 2522 406 2525 526
rect 2570 453 2573 526
rect 2634 523 2637 573
rect 2666 566 2669 603
rect 2658 563 2669 566
rect 2658 466 2661 563
rect 2658 463 2669 466
rect 2506 403 2525 406
rect 2498 333 2501 346
rect 2490 283 2493 316
rect 2482 273 2493 276
rect 2482 213 2485 226
rect 2490 213 2493 273
rect 2506 246 2509 356
rect 2514 323 2517 403
rect 2538 346 2541 416
rect 2610 413 2613 426
rect 2666 413 2669 463
rect 2586 366 2589 406
rect 2522 343 2541 346
rect 2522 333 2525 343
rect 2530 323 2533 336
rect 2538 333 2541 343
rect 2582 363 2589 366
rect 2498 243 2509 246
rect 2498 216 2501 243
rect 2506 223 2517 226
rect 2522 223 2525 236
rect 2498 213 2509 216
rect 2530 203 2533 316
rect 2538 213 2541 306
rect 2546 216 2549 326
rect 2562 303 2565 336
rect 2570 323 2573 336
rect 2570 293 2573 316
rect 2582 306 2585 363
rect 2618 313 2621 326
rect 2634 323 2637 336
rect 2582 303 2589 306
rect 2554 223 2557 236
rect 2546 213 2557 216
rect 2570 213 2573 226
rect 2554 193 2557 206
rect 2586 203 2589 303
rect 2610 193 2613 216
rect 2666 213 2669 296
rect 1242 93 1249 96
rect 1242 73 1245 93
rect 2686 37 2706 2603
rect 2710 13 2730 2627
<< metal3 >>
rect 1161 2562 1262 2567
rect 1161 2557 1166 2562
rect 889 2552 982 2557
rect 1137 2552 1166 2557
rect 1257 2557 1262 2562
rect 1353 2562 1478 2567
rect 1353 2557 1358 2562
rect 1257 2552 1310 2557
rect 1329 2552 1358 2557
rect 1473 2557 1478 2562
rect 1473 2552 1590 2557
rect 1921 2552 2158 2557
rect 1921 2547 1926 2552
rect 265 2542 358 2547
rect 393 2542 486 2547
rect 569 2542 662 2547
rect 697 2542 790 2547
rect 1169 2542 1230 2547
rect 1369 2542 1462 2547
rect 1689 2542 1782 2547
rect 1841 2542 1926 2547
rect 2153 2547 2158 2552
rect 2153 2542 2214 2547
rect 2305 2542 2566 2547
rect 273 2532 430 2537
rect 561 2527 566 2537
rect 577 2532 734 2537
rect 993 2532 1246 2537
rect 1313 2532 1358 2537
rect 1377 2532 1534 2537
rect 2049 2532 2118 2537
rect 993 2527 998 2532
rect 1961 2527 2054 2532
rect 2113 2527 2118 2532
rect 265 2522 358 2527
rect 353 2517 358 2522
rect 433 2522 550 2527
rect 561 2522 678 2527
rect 689 2522 830 2527
rect 897 2522 998 2527
rect 1017 2522 1118 2527
rect 1353 2522 1478 2527
rect 1489 2522 1630 2527
rect 1937 2522 1966 2527
rect 2113 2522 2142 2527
rect 433 2517 438 2522
rect 121 2512 206 2517
rect 353 2512 438 2517
rect 545 2507 550 2522
rect 673 2517 678 2522
rect 1473 2517 1478 2522
rect 673 2512 766 2517
rect 1025 2512 1142 2517
rect 1473 2512 1566 2517
rect 1665 2512 1710 2517
rect 1921 2512 1990 2517
rect 2065 2512 2294 2517
rect 2417 2512 2462 2517
rect 73 2502 182 2507
rect 545 2502 574 2507
rect 1009 2502 1070 2507
rect 1065 2497 1070 2502
rect 1153 2502 1294 2507
rect 1681 2502 1758 2507
rect 1945 2502 2054 2507
rect 2401 2502 2518 2507
rect 1153 2497 1158 2502
rect 897 2492 1046 2497
rect 1065 2492 1158 2497
rect 1969 2492 1998 2497
rect 1993 2487 1998 2492
rect 2145 2492 2174 2497
rect 2145 2487 2150 2492
rect 1993 2482 2150 2487
rect 857 2462 1022 2467
rect 1065 2452 1222 2457
rect 2425 2452 2470 2457
rect 929 2442 1022 2447
rect 1017 2437 1022 2442
rect 1137 2442 1166 2447
rect 1137 2437 1142 2442
rect 785 2432 950 2437
rect 1017 2432 1142 2437
rect 1425 2432 1526 2437
rect 1625 2432 1694 2437
rect 1873 2432 1918 2437
rect 1929 2432 2038 2437
rect 129 2422 222 2427
rect 289 2422 398 2427
rect 497 2422 566 2427
rect 761 2422 822 2427
rect 881 2422 998 2427
rect 1777 2422 1814 2427
rect 1905 2422 1966 2427
rect 2361 2422 2462 2427
rect 2481 2422 2646 2427
rect 1777 2417 1782 2422
rect 73 2412 150 2417
rect 385 2412 494 2417
rect 625 2412 774 2417
rect 1705 2412 1782 2417
rect 2201 2412 2390 2417
rect 1601 2402 1694 2407
rect 2233 2402 2414 2407
rect 129 2392 198 2397
rect 401 2392 486 2397
rect 585 2392 646 2397
rect 681 2392 854 2397
rect 1073 2392 1166 2397
rect 1201 2392 1446 2397
rect 1913 2392 1950 2397
rect 2289 2392 2558 2397
rect 417 2382 518 2387
rect 1137 2382 1222 2387
rect 2305 2382 2414 2387
rect 2409 2377 2414 2382
rect 2545 2382 2574 2387
rect 2545 2377 2550 2382
rect 2297 2372 2318 2377
rect 2409 2372 2550 2377
rect 121 2352 278 2357
rect 289 2352 366 2357
rect 473 2352 590 2357
rect 777 2352 910 2357
rect 1249 2352 1438 2357
rect 145 2342 230 2347
rect 1385 2342 1566 2347
rect 201 2332 382 2337
rect 569 2332 654 2337
rect 801 2332 1102 2337
rect 1337 2332 1494 2337
rect 1593 2332 1670 2337
rect 497 2322 790 2327
rect 785 2317 790 2322
rect 873 2322 902 2327
rect 1713 2322 1790 2327
rect 1953 2322 2030 2327
rect 2057 2322 2150 2327
rect 2273 2322 2310 2327
rect 873 2317 878 2322
rect 529 2312 702 2317
rect 785 2312 878 2317
rect 1009 2312 1038 2317
rect 1033 2307 1038 2312
rect 1113 2312 1262 2317
rect 1545 2312 1630 2317
rect 1665 2312 1742 2317
rect 2001 2312 2030 2317
rect 1113 2307 1118 2312
rect 2025 2307 2030 2312
rect 2097 2312 2126 2317
rect 2153 2312 2414 2317
rect 2441 2312 2670 2317
rect 2097 2307 2102 2312
rect 1033 2302 1118 2307
rect 1697 2302 1822 2307
rect 2025 2302 2102 2307
rect 1449 2292 1542 2297
rect 1649 2292 1734 2297
rect 2369 2252 2470 2257
rect 809 2242 942 2247
rect 993 2242 1086 2247
rect 1161 2242 1350 2247
rect 2265 2242 2318 2247
rect 809 2237 814 2242
rect 785 2232 814 2237
rect 937 2237 942 2242
rect 937 2232 966 2237
rect 1145 2232 1222 2237
rect 129 2222 198 2227
rect 281 2222 366 2227
rect 393 2222 462 2227
rect 985 2222 1014 2227
rect 745 2217 886 2222
rect 1009 2217 1014 2222
rect 1161 2222 1206 2227
rect 1161 2217 1166 2222
rect 185 2212 254 2217
rect 305 2212 406 2217
rect 529 2212 638 2217
rect 721 2212 750 2217
rect 881 2212 974 2217
rect 1009 2212 1166 2217
rect 193 2202 302 2207
rect 409 2202 518 2207
rect 545 2202 870 2207
rect 865 2197 870 2202
rect 1217 2197 1222 2232
rect 1441 2232 1558 2237
rect 1721 2232 1790 2237
rect 2249 2232 2286 2237
rect 2393 2232 2446 2237
rect 1441 2227 1446 2232
rect 1417 2222 1446 2227
rect 1553 2227 1558 2232
rect 1553 2222 1582 2227
rect 1641 2222 1662 2227
rect 1905 2222 1966 2227
rect 2241 2222 2302 2227
rect 2449 2222 2654 2227
rect 1393 2212 1598 2217
rect 1937 2212 2038 2217
rect 2329 2212 2430 2217
rect 1489 2202 1526 2207
rect 1873 2202 1926 2207
rect 2209 2202 2262 2207
rect 2537 2202 2654 2207
rect 1489 2197 1494 2202
rect 73 2192 134 2197
rect 529 2192 846 2197
rect 865 2192 966 2197
rect 1185 2192 1222 2197
rect 1345 2192 1494 2197
rect 2289 2192 2550 2197
rect 393 2182 422 2187
rect 417 2177 422 2182
rect 513 2182 646 2187
rect 745 2182 886 2187
rect 985 2182 1062 2187
rect 1465 2182 1550 2187
rect 2417 2182 2446 2187
rect 513 2177 518 2182
rect 985 2177 990 2182
rect 417 2172 518 2177
rect 537 2172 630 2177
rect 865 2172 990 2177
rect 1057 2177 1062 2182
rect 2441 2177 2446 2182
rect 2545 2182 2574 2187
rect 2545 2177 2550 2182
rect 1057 2172 1086 2177
rect 1569 2172 1686 2177
rect 1481 2167 1574 2172
rect 1681 2167 1686 2172
rect 1913 2172 2014 2177
rect 2441 2172 2550 2177
rect 1913 2167 1918 2172
rect 849 2162 878 2167
rect 873 2157 878 2162
rect 1001 2162 1046 2167
rect 1457 2162 1486 2167
rect 1681 2162 1710 2167
rect 1825 2162 1918 2167
rect 2009 2167 2014 2172
rect 2009 2162 2166 2167
rect 1001 2157 1006 2162
rect 873 2152 1006 2157
rect 1121 2152 1198 2157
rect 1433 2152 1590 2157
rect 1601 2152 1654 2157
rect 1929 2152 1998 2157
rect 2057 2152 2270 2157
rect 1993 2147 2062 2152
rect 145 2142 182 2147
rect 377 2142 638 2147
rect 1417 2142 1438 2147
rect 1465 2142 1566 2147
rect 1593 2142 1726 2147
rect 2081 2142 2134 2147
rect 177 2137 182 2142
rect 1073 2137 1190 2142
rect 177 2132 214 2137
rect 729 2132 1078 2137
rect 1185 2132 1270 2137
rect 1385 2132 1414 2137
rect 273 2122 358 2127
rect 1097 2122 1158 2127
rect 273 2117 278 2122
rect 249 2112 278 2117
rect 353 2117 358 2122
rect 1265 2117 1270 2132
rect 1409 2127 1414 2132
rect 1497 2132 1606 2137
rect 1937 2132 2286 2137
rect 2361 2132 2502 2137
rect 1497 2127 1502 2132
rect 1289 2122 1374 2127
rect 1409 2122 1502 2127
rect 1625 2122 1702 2127
rect 1897 2122 2006 2127
rect 2145 2122 2238 2127
rect 353 2112 494 2117
rect 529 2112 718 2117
rect 713 2107 718 2112
rect 865 2112 894 2117
rect 945 2112 974 2117
rect 865 2107 870 2112
rect 121 2102 238 2107
rect 233 2097 238 2102
rect 321 2102 350 2107
rect 657 2102 686 2107
rect 713 2102 870 2107
rect 969 2107 974 2112
rect 1057 2112 1086 2117
rect 1265 2112 1286 2117
rect 1849 2112 1926 2117
rect 1945 2112 1998 2117
rect 2113 2112 2174 2117
rect 1057 2107 1062 2112
rect 969 2102 1062 2107
rect 1281 2107 1286 2112
rect 1281 2102 1382 2107
rect 1609 2102 1646 2107
rect 1665 2102 1750 2107
rect 2185 2102 2302 2107
rect 321 2097 326 2102
rect 233 2092 326 2097
rect 505 2072 654 2077
rect 505 2067 510 2072
rect 433 2062 510 2067
rect 649 2067 654 2072
rect 649 2062 678 2067
rect 2273 2062 2342 2067
rect 545 2052 774 2057
rect 865 2052 926 2057
rect 961 2052 1070 2057
rect 961 2047 966 2052
rect 329 2042 414 2047
rect 521 2042 718 2047
rect 737 2042 814 2047
rect 849 2042 966 2047
rect 1065 2047 1070 2052
rect 2001 2052 2086 2057
rect 2001 2047 2006 2052
rect 1065 2042 1094 2047
rect 1217 2042 1390 2047
rect 1977 2042 2006 2047
rect 2081 2047 2086 2052
rect 2081 2042 2110 2047
rect 329 2037 334 2042
rect 305 2032 334 2037
rect 409 2037 414 2042
rect 409 2032 454 2037
rect 537 2032 646 2037
rect 777 2032 910 2037
rect 1041 2032 1158 2037
rect 1041 2027 1046 2032
rect 1217 2027 1222 2042
rect 1385 2037 1390 2042
rect 1385 2032 1502 2037
rect 1545 2032 1662 2037
rect 1873 2032 1918 2037
rect 1929 2032 2038 2037
rect 2089 2032 2198 2037
rect 1545 2027 1550 2032
rect 321 2022 398 2027
rect 465 2022 654 2027
rect 665 2022 854 2027
rect 897 2022 1046 2027
rect 1065 2022 1134 2027
rect 1153 2022 1222 2027
rect 1281 2022 1318 2027
rect 1521 2022 1550 2027
rect 1657 2027 1662 2032
rect 1657 2022 1686 2027
rect 1905 2022 1966 2027
rect 2305 2022 2430 2027
rect 2569 2022 2614 2027
rect 393 2017 470 2022
rect 529 2012 886 2017
rect 993 2007 1118 2012
rect 1153 2007 1158 2022
rect 1313 2017 1318 2022
rect 1313 2012 1374 2017
rect 1393 2012 1502 2017
rect 2161 2012 2238 2017
rect 2441 2012 2662 2017
rect 1393 2007 1398 2012
rect 265 2002 398 2007
rect 433 2002 494 2007
rect 513 2002 670 2007
rect 681 2002 830 2007
rect 897 2002 998 2007
rect 1113 2002 1182 2007
rect 1201 2002 1278 2007
rect 1353 2002 1398 2007
rect 1497 2007 1502 2012
rect 1497 2002 1678 2007
rect 1921 2002 1950 2007
rect 265 1997 270 2002
rect 241 1992 270 1997
rect 393 1997 398 2002
rect 825 1997 902 2002
rect 1201 1997 1206 2002
rect 393 1992 422 1997
rect 537 1992 662 1997
rect 1009 1992 1206 1997
rect 1273 1997 1278 2002
rect 1273 1992 1326 1997
rect 1377 1992 1494 1997
rect 2537 1992 2558 1997
rect 681 1987 806 1992
rect 217 1982 294 1987
rect 313 1982 414 1987
rect 505 1982 686 1987
rect 801 1982 934 1987
rect 945 1982 1262 1987
rect 1513 1982 1582 1987
rect 289 1977 294 1982
rect 929 1977 934 1982
rect 1513 1977 1518 1982
rect 289 1972 878 1977
rect 929 1972 1134 1977
rect 1233 1972 1518 1977
rect 1577 1977 1582 1982
rect 1577 1972 1774 1977
rect 113 1962 246 1967
rect 273 1962 718 1967
rect 273 1957 278 1962
rect 713 1957 718 1962
rect 809 1962 998 1967
rect 1505 1962 1598 1967
rect 2017 1962 2134 1967
rect 809 1957 814 1962
rect 249 1952 278 1957
rect 289 1952 526 1957
rect 585 1952 694 1957
rect 713 1952 814 1957
rect 1161 1952 1262 1957
rect 1161 1947 1166 1952
rect 305 1942 478 1947
rect 905 1942 1118 1947
rect 1137 1942 1166 1947
rect 1257 1947 1262 1952
rect 1505 1947 1510 1962
rect 2017 1957 2022 1962
rect 1633 1947 1638 1957
rect 1993 1952 2022 1957
rect 2129 1957 2134 1962
rect 2321 1962 2350 1967
rect 2321 1957 2326 1962
rect 2129 1952 2326 1957
rect 1257 1942 1286 1947
rect 1337 1942 1510 1947
rect 1537 1942 1638 1947
rect 1953 1942 2118 1947
rect 2401 1942 2502 1947
rect 905 1937 910 1942
rect 153 1932 230 1937
rect 265 1932 510 1937
rect 153 1927 158 1932
rect 129 1922 158 1927
rect 225 1927 230 1932
rect 505 1927 510 1932
rect 641 1932 758 1937
rect 881 1932 910 1937
rect 1113 1937 1118 1942
rect 1113 1932 1150 1937
rect 1161 1932 1534 1937
rect 641 1927 646 1932
rect 1529 1927 1534 1932
rect 1601 1932 1766 1937
rect 1601 1927 1606 1932
rect 2073 1927 2166 1932
rect 2401 1927 2406 1942
rect 2497 1937 2502 1942
rect 2497 1932 2526 1937
rect 225 1922 278 1927
rect 505 1922 646 1927
rect 865 1922 1062 1927
rect 1321 1922 1510 1927
rect 1529 1922 1606 1927
rect 1961 1922 1990 1927
rect 1057 1917 1062 1922
rect 1985 1917 1990 1922
rect 2049 1922 2078 1927
rect 2161 1922 2406 1927
rect 2425 1922 2646 1927
rect 2049 1917 2054 1922
rect 137 1912 254 1917
rect 321 1912 430 1917
rect 665 1912 686 1917
rect 1057 1912 1094 1917
rect 1089 1907 1094 1912
rect 1153 1912 1182 1917
rect 1249 1912 1374 1917
rect 1985 1912 2054 1917
rect 2073 1912 2142 1917
rect 2233 1912 2286 1917
rect 2553 1912 2598 1917
rect 1153 1907 1158 1912
rect 313 1902 342 1907
rect 425 1902 454 1907
rect 993 1902 1054 1907
rect 1089 1902 1158 1907
rect 1329 1902 1446 1907
rect 337 1897 430 1902
rect 1441 1897 1446 1902
rect 1505 1902 1902 1907
rect 2201 1902 2230 1907
rect 1505 1897 1510 1902
rect 825 1892 886 1897
rect 1033 1892 1070 1897
rect 1337 1892 1382 1897
rect 1441 1892 1510 1897
rect 2225 1897 2230 1902
rect 2305 1902 2334 1907
rect 2521 1902 2550 1907
rect 2305 1897 2310 1902
rect 2225 1892 2310 1897
rect 145 1882 302 1887
rect 297 1877 302 1882
rect 393 1882 422 1887
rect 545 1882 622 1887
rect 697 1882 806 1887
rect 393 1877 398 1882
rect 697 1877 702 1882
rect 297 1872 398 1877
rect 673 1872 702 1877
rect 801 1877 806 1882
rect 801 1872 878 1877
rect 961 1872 1102 1877
rect 2553 1872 2670 1877
rect 961 1867 966 1872
rect 689 1862 966 1867
rect 1097 1867 1102 1872
rect 1097 1862 1446 1867
rect 689 1857 694 1862
rect 473 1852 694 1857
rect 705 1852 1086 1857
rect 729 1842 902 1847
rect 1353 1842 1454 1847
rect 1545 1842 1590 1847
rect 617 1837 694 1842
rect 537 1832 622 1837
rect 689 1832 718 1837
rect 793 1832 1038 1837
rect 1121 1832 1222 1837
rect 1233 1832 1286 1837
rect 1337 1832 1366 1837
rect 2129 1832 2182 1837
rect 2281 1832 2326 1837
rect 2385 1832 2486 1837
rect 713 1827 798 1832
rect 1233 1827 1238 1832
rect 1361 1827 1366 1832
rect 633 1822 678 1827
rect 817 1822 838 1827
rect 1073 1822 1238 1827
rect 1249 1822 1350 1827
rect 1361 1822 1390 1827
rect 1497 1822 1534 1827
rect 1553 1822 1654 1827
rect 1753 1822 1798 1827
rect 2313 1822 2374 1827
rect 657 1812 1126 1817
rect 1329 1812 1438 1817
rect 1569 1812 1630 1817
rect 1817 1812 1894 1817
rect 2345 1812 2446 1817
rect 1817 1807 1822 1812
rect 545 1802 614 1807
rect 1105 1802 1142 1807
rect 1177 1802 1254 1807
rect 1289 1802 1518 1807
rect 1641 1802 1822 1807
rect 1889 1807 1894 1812
rect 1889 1802 1918 1807
rect 2113 1802 2262 1807
rect 2465 1802 2670 1807
rect 545 1797 550 1802
rect 521 1792 550 1797
rect 609 1797 614 1802
rect 609 1792 654 1797
rect 673 1792 830 1797
rect 849 1792 918 1797
rect 929 1792 1006 1797
rect 1033 1792 1190 1797
rect 1297 1792 1406 1797
rect 1425 1792 1470 1797
rect 1617 1792 1678 1797
rect 1873 1792 2014 1797
rect 2361 1792 2454 1797
rect 673 1787 678 1792
rect 257 1782 382 1787
rect 489 1782 678 1787
rect 825 1787 830 1792
rect 2449 1787 2454 1792
rect 2537 1792 2566 1797
rect 2537 1787 2542 1792
rect 825 1782 1726 1787
rect 257 1777 262 1782
rect 121 1772 262 1777
rect 377 1777 382 1782
rect 1721 1777 1726 1782
rect 1825 1782 1854 1787
rect 1897 1782 2142 1787
rect 2449 1782 2542 1787
rect 1825 1777 1830 1782
rect 377 1772 734 1777
rect 745 1772 846 1777
rect 913 1772 1030 1777
rect 1057 1772 1110 1777
rect 1153 1772 1310 1777
rect 1321 1772 1366 1777
rect 1721 1772 1830 1777
rect 2041 1772 2126 1777
rect 1025 1767 1030 1772
rect 313 1762 790 1767
rect 857 1762 1014 1767
rect 1025 1762 1262 1767
rect 1337 1762 1414 1767
rect 1609 1762 1686 1767
rect 2001 1762 2030 1767
rect 785 1757 862 1762
rect 1609 1757 1614 1762
rect 273 1752 374 1757
rect 481 1752 558 1757
rect 625 1752 766 1757
rect 1057 1752 1182 1757
rect 369 1747 374 1752
rect 1201 1747 1206 1757
rect 1233 1752 1550 1757
rect 1577 1752 1614 1757
rect 1681 1747 1686 1762
rect 2025 1757 2030 1762
rect 2097 1762 2126 1767
rect 2369 1762 2510 1767
rect 2097 1757 2102 1762
rect 2369 1757 2374 1762
rect 2025 1752 2102 1757
rect 2345 1752 2374 1757
rect 2505 1757 2510 1762
rect 2505 1752 2534 1757
rect 185 1742 302 1747
rect 369 1742 462 1747
rect 521 1742 598 1747
rect 649 1742 718 1747
rect 865 1742 966 1747
rect 1073 1742 1150 1747
rect 1161 1742 1206 1747
rect 217 1732 326 1737
rect 377 1732 902 1737
rect 937 1732 1046 1737
rect 1097 1732 1278 1737
rect 1313 1727 1318 1747
rect 1369 1742 1462 1747
rect 1625 1742 1670 1747
rect 1681 1742 1718 1747
rect 1785 1742 1862 1747
rect 2233 1742 2494 1747
rect 2561 1742 2590 1747
rect 1785 1737 1790 1742
rect 1425 1732 1614 1737
rect 1713 1732 1790 1737
rect 1857 1737 1862 1742
rect 2489 1737 2566 1742
rect 1857 1732 1966 1737
rect 1609 1727 1718 1732
rect 137 1722 174 1727
rect 169 1717 174 1722
rect 257 1722 390 1727
rect 473 1722 542 1727
rect 585 1722 710 1727
rect 921 1722 1070 1727
rect 1113 1722 1222 1727
rect 1313 1722 1502 1727
rect 1737 1722 1878 1727
rect 2345 1722 2446 1727
rect 257 1717 262 1722
rect 385 1717 390 1722
rect 169 1712 262 1717
rect 281 1712 374 1717
rect 385 1712 550 1717
rect 849 1712 966 1717
rect 1033 1712 1078 1717
rect 1265 1712 1350 1717
rect 1361 1712 1398 1717
rect 1505 1712 1654 1717
rect 1785 1712 1830 1717
rect 1985 1712 2022 1717
rect 2313 1712 2374 1717
rect 2457 1712 2670 1717
rect 1073 1707 1078 1712
rect 1393 1707 1486 1712
rect 425 1702 470 1707
rect 569 1702 646 1707
rect 489 1697 574 1702
rect 641 1697 646 1702
rect 689 1702 774 1707
rect 929 1702 958 1707
rect 985 1702 1062 1707
rect 1073 1702 1358 1707
rect 1481 1702 1526 1707
rect 1729 1702 1750 1707
rect 1945 1702 2014 1707
rect 2281 1702 2326 1707
rect 2409 1702 2454 1707
rect 689 1697 694 1702
rect 337 1692 382 1697
rect 433 1692 494 1697
rect 641 1692 694 1697
rect 769 1697 774 1702
rect 769 1692 798 1697
rect 969 1692 1030 1697
rect 1441 1692 1750 1697
rect 1273 1687 1422 1692
rect 1745 1687 1750 1692
rect 1841 1692 1958 1697
rect 1977 1692 2038 1697
rect 1841 1687 1846 1692
rect 345 1682 750 1687
rect 745 1677 750 1682
rect 809 1682 982 1687
rect 1121 1682 1198 1687
rect 1249 1682 1278 1687
rect 1417 1682 1590 1687
rect 1745 1682 1846 1687
rect 1953 1687 1958 1692
rect 1953 1682 2006 1687
rect 809 1677 814 1682
rect 313 1672 438 1677
rect 513 1672 630 1677
rect 745 1672 814 1677
rect 1105 1672 1662 1677
rect 177 1662 294 1667
rect 377 1662 694 1667
rect 873 1662 1038 1667
rect 1161 1662 1726 1667
rect 1961 1662 1998 1667
rect 177 1657 182 1662
rect 153 1652 182 1657
rect 289 1657 294 1662
rect 873 1657 878 1662
rect 289 1652 878 1657
rect 1033 1657 1038 1662
rect 1033 1652 1966 1657
rect 913 1647 1014 1652
rect 65 1642 142 1647
rect 137 1637 142 1642
rect 257 1642 638 1647
rect 649 1642 678 1647
rect 889 1642 918 1647
rect 1009 1642 1094 1647
rect 1313 1642 1430 1647
rect 1521 1642 1750 1647
rect 257 1637 262 1642
rect 1425 1637 1526 1642
rect 137 1632 262 1637
rect 297 1632 326 1637
rect 409 1632 446 1637
rect 537 1632 662 1637
rect 753 1632 1022 1637
rect 1201 1632 1326 1637
rect 1545 1632 1694 1637
rect 1817 1632 1862 1637
rect 2033 1632 2150 1637
rect 1097 1627 1182 1632
rect 433 1622 486 1627
rect 497 1622 1102 1627
rect 1177 1622 1246 1627
rect 481 1617 486 1622
rect 1241 1617 1246 1622
rect 1337 1622 1494 1627
rect 1337 1617 1342 1622
rect 281 1612 470 1617
rect 481 1612 998 1617
rect 1113 1612 1150 1617
rect 1161 1612 1222 1617
rect 1241 1612 1342 1617
rect 1489 1617 1494 1622
rect 1641 1622 1830 1627
rect 2153 1622 2246 1627
rect 2265 1622 2294 1627
rect 1641 1617 1646 1622
rect 1489 1612 1646 1617
rect 1793 1612 1838 1617
rect 2113 1607 2118 1617
rect 593 1602 886 1607
rect 945 1602 1046 1607
rect 1665 1602 1702 1607
rect 2113 1602 2134 1607
rect 1161 1597 1270 1602
rect 289 1592 366 1597
rect 529 1592 678 1597
rect 689 1592 798 1597
rect 1057 1592 1166 1597
rect 1265 1592 1382 1597
rect 1393 1592 1470 1597
rect 1681 1592 1790 1597
rect 1801 1592 1854 1597
rect 1881 1592 1950 1597
rect 793 1587 894 1592
rect 1057 1587 1062 1592
rect 1377 1587 1382 1592
rect 233 1582 262 1587
rect 377 1582 422 1587
rect 449 1582 494 1587
rect 545 1582 574 1587
rect 585 1582 702 1587
rect 889 1582 1062 1587
rect 1177 1582 1254 1587
rect 1377 1582 1478 1587
rect 1865 1582 1910 1587
rect 2233 1582 2286 1587
rect 257 1577 382 1582
rect 401 1572 598 1577
rect 617 1572 726 1577
rect 801 1572 870 1577
rect 1081 1572 1158 1577
rect 1185 1572 1566 1577
rect 249 1562 350 1567
rect 449 1562 494 1567
rect 529 1562 614 1567
rect 625 1562 758 1567
rect 913 1562 982 1567
rect 1137 1562 1190 1567
rect 1377 1562 1526 1567
rect 1201 1557 1382 1562
rect 2561 1557 2566 1567
rect 177 1552 806 1557
rect 825 1552 942 1557
rect 993 1552 1206 1557
rect 1889 1552 1966 1557
rect 2057 1552 2158 1557
rect 2481 1552 2654 1557
rect 145 1542 246 1547
rect 329 1542 1022 1547
rect 1193 1542 1286 1547
rect 1353 1542 1422 1547
rect 1465 1542 1542 1547
rect 1753 1542 1830 1547
rect 1849 1542 1902 1547
rect 2513 1542 2622 1547
rect 1753 1537 1758 1542
rect 225 1532 302 1537
rect 417 1532 566 1537
rect 625 1532 726 1537
rect 793 1532 870 1537
rect 889 1532 974 1537
rect 1041 1532 1126 1537
rect 1609 1532 1758 1537
rect 1825 1537 1830 1542
rect 1825 1532 1862 1537
rect 1929 1532 2230 1537
rect 2433 1532 2542 1537
rect 561 1527 566 1532
rect 281 1522 470 1527
rect 481 1522 550 1527
rect 561 1522 1070 1527
rect 1337 1522 1382 1527
rect 1881 1522 1926 1527
rect 1985 1522 2054 1527
rect 1377 1517 1382 1522
rect 145 1512 166 1517
rect 337 1512 382 1517
rect 489 1512 1230 1517
rect 1377 1512 1614 1517
rect 1697 1512 1886 1517
rect 1985 1512 1990 1522
rect 2033 1512 2094 1517
rect 2321 1512 2342 1517
rect 2353 1512 2446 1517
rect 2545 1512 2662 1517
rect 289 1502 414 1507
rect 545 1502 1094 1507
rect 1185 1502 1430 1507
rect 1513 1502 1542 1507
rect 2025 1502 2174 1507
rect 2289 1502 2318 1507
rect 1609 1497 1782 1502
rect 2313 1497 2318 1502
rect 2385 1502 2414 1507
rect 2433 1502 2574 1507
rect 2385 1497 2390 1502
rect 553 1492 614 1497
rect 705 1492 790 1497
rect 825 1492 974 1497
rect 1225 1492 1614 1497
rect 1777 1492 1974 1497
rect 2113 1492 2182 1497
rect 2313 1492 2390 1497
rect 465 1487 534 1492
rect 1969 1487 1974 1492
rect 393 1482 470 1487
rect 529 1482 1118 1487
rect 1441 1482 1494 1487
rect 1593 1482 1742 1487
rect 1969 1482 2182 1487
rect 1161 1477 1310 1482
rect 1489 1477 1598 1482
rect 481 1472 670 1477
rect 689 1472 958 1477
rect 993 1472 1166 1477
rect 1305 1472 1470 1477
rect 1465 1467 1470 1472
rect 1617 1472 1670 1477
rect 1617 1467 1622 1472
rect 169 1462 1294 1467
rect 1465 1462 1622 1467
rect 1665 1467 1670 1472
rect 1737 1472 1854 1477
rect 1737 1467 1742 1472
rect 1665 1462 1742 1467
rect 2249 1462 2302 1467
rect 409 1452 430 1457
rect 521 1452 662 1457
rect 961 1452 1334 1457
rect 1993 1452 2070 1457
rect 745 1447 886 1452
rect 385 1442 430 1447
rect 441 1442 750 1447
rect 881 1442 1526 1447
rect 1553 1442 1622 1447
rect 1553 1437 1558 1442
rect 185 1432 238 1437
rect 353 1432 422 1437
rect 513 1432 630 1437
rect 761 1432 870 1437
rect 993 1432 1382 1437
rect 993 1427 998 1432
rect 1377 1427 1382 1432
rect 1537 1432 1558 1437
rect 1617 1437 1622 1442
rect 1617 1432 1982 1437
rect 1537 1427 1542 1432
rect 1977 1427 1982 1432
rect 2073 1432 2102 1437
rect 2073 1427 2078 1432
rect 225 1422 254 1427
rect 361 1422 998 1427
rect 1017 1422 1334 1427
rect 1377 1422 1542 1427
rect 1569 1422 1606 1427
rect 1977 1422 2078 1427
rect 2465 1422 2510 1427
rect 2585 1422 2630 1427
rect 225 1417 230 1422
rect 1329 1417 1334 1422
rect 185 1412 230 1417
rect 249 1412 310 1417
rect 337 1412 406 1417
rect 489 1412 598 1417
rect 697 1412 718 1417
rect 873 1412 910 1417
rect 1329 1412 1358 1417
rect 785 1407 854 1412
rect 1065 1407 1198 1412
rect 1545 1407 1670 1412
rect 193 1402 278 1407
rect 385 1402 790 1407
rect 849 1402 1070 1407
rect 1193 1402 1550 1407
rect 1665 1402 1694 1407
rect 2153 1402 2262 1407
rect 289 1392 382 1397
rect 441 1392 494 1397
rect 561 1392 590 1397
rect 649 1392 734 1397
rect 801 1392 854 1397
rect 849 1387 854 1392
rect 953 1392 982 1397
rect 1081 1392 1182 1397
rect 1273 1392 1350 1397
rect 1561 1392 1590 1397
rect 953 1387 958 1392
rect 297 1382 830 1387
rect 849 1382 958 1387
rect 1585 1387 1590 1392
rect 1649 1392 1726 1397
rect 2281 1392 2486 1397
rect 2505 1392 2526 1397
rect 1649 1387 1654 1392
rect 2481 1387 2486 1392
rect 1585 1382 1654 1387
rect 1985 1382 2070 1387
rect 2481 1382 2590 1387
rect 1985 1377 1990 1382
rect 281 1372 350 1377
rect 441 1372 470 1377
rect 569 1372 598 1377
rect 657 1372 814 1377
rect 1673 1372 1702 1377
rect 1801 1372 1846 1377
rect 1961 1372 1990 1377
rect 2065 1377 2070 1382
rect 2065 1372 2126 1377
rect 345 1367 446 1372
rect 657 1367 662 1372
rect 81 1362 326 1367
rect 529 1362 566 1367
rect 577 1362 662 1367
rect 673 1362 806 1367
rect 833 1362 878 1367
rect 1001 1362 1462 1367
rect 1993 1362 2054 1367
rect 81 1302 86 1362
rect 97 1352 222 1357
rect 97 1312 102 1352
rect 113 1342 158 1347
rect 217 1342 254 1347
rect 113 1297 118 1342
rect 177 1332 246 1337
rect 305 1332 310 1357
rect 321 1347 326 1362
rect 577 1357 582 1362
rect 353 1352 582 1357
rect 593 1352 630 1357
rect 673 1347 678 1362
rect 321 1342 342 1347
rect 337 1337 342 1342
rect 497 1342 678 1347
rect 497 1337 502 1342
rect 689 1337 694 1357
rect 337 1332 502 1337
rect 521 1332 694 1337
rect 721 1352 750 1357
rect 817 1352 846 1357
rect 1201 1352 1230 1357
rect 1553 1352 1646 1357
rect 177 1327 182 1332
rect 137 1322 182 1327
rect 217 1322 302 1327
rect 617 1322 646 1327
rect 721 1322 726 1352
rect 737 1342 806 1347
rect 817 1327 822 1352
rect 1201 1347 1206 1352
rect 1393 1347 1510 1352
rect 1001 1342 1054 1347
rect 1089 1342 1206 1347
rect 1369 1342 1398 1347
rect 1505 1342 1534 1347
rect 777 1322 822 1327
rect 833 1317 838 1337
rect 929 1332 1022 1337
rect 1041 1332 1070 1337
rect 1041 1327 1046 1332
rect 1089 1327 1094 1342
rect 1553 1337 1558 1352
rect 1641 1347 1646 1352
rect 2145 1352 2246 1357
rect 2145 1347 2150 1352
rect 1641 1342 1782 1347
rect 2025 1342 2150 1347
rect 2241 1347 2246 1352
rect 2337 1352 2422 1357
rect 2337 1347 2342 1352
rect 2241 1342 2270 1347
rect 2313 1342 2342 1347
rect 2417 1347 2422 1352
rect 2417 1342 2446 1347
rect 1281 1332 1558 1337
rect 1809 1332 1830 1337
rect 2049 1332 2078 1337
rect 945 1322 1046 1327
rect 1057 1322 1094 1327
rect 1297 1322 1462 1327
rect 1553 1322 1630 1327
rect 945 1317 950 1322
rect 129 1312 166 1317
rect 249 1312 342 1317
rect 441 1312 478 1317
rect 657 1312 734 1317
rect 801 1312 838 1317
rect 889 1312 950 1317
rect 969 1312 1070 1317
rect 1185 1312 1286 1317
rect 1353 1312 1414 1317
rect 1481 1312 1534 1317
rect 1809 1312 1814 1332
rect 2073 1327 2078 1332
rect 2153 1332 2230 1337
rect 2297 1332 2454 1337
rect 2153 1327 2158 1332
rect 2225 1327 2302 1332
rect 2449 1327 2454 1332
rect 2073 1322 2158 1327
rect 2321 1322 2350 1327
rect 2345 1317 2350 1322
rect 2409 1322 2438 1327
rect 2449 1322 2534 1327
rect 2409 1317 2414 1322
rect 2177 1312 2270 1317
rect 2345 1312 2414 1317
rect 2537 1312 2670 1317
rect 137 1302 238 1307
rect 297 1302 590 1307
rect 609 1302 630 1307
rect 793 1302 870 1307
rect 897 1302 990 1307
rect 1193 1302 1350 1307
rect 1473 1302 1614 1307
rect 1961 1302 2062 1307
rect 233 1297 302 1302
rect 89 1292 118 1297
rect 321 1292 350 1297
rect 409 1292 678 1297
rect 713 1292 822 1297
rect 873 1292 918 1297
rect 929 1292 1086 1297
rect 1217 1292 1246 1297
rect 73 1282 102 1287
rect 97 1277 102 1282
rect 241 1282 750 1287
rect 769 1282 1102 1287
rect 241 1277 246 1282
rect 769 1277 774 1282
rect 1241 1277 1246 1292
rect 1569 1292 1670 1297
rect 2249 1292 2454 1297
rect 1569 1277 1574 1292
rect 1673 1282 1718 1287
rect 97 1272 246 1277
rect 265 1272 606 1277
rect 641 1272 774 1277
rect 857 1272 1022 1277
rect 1241 1272 1574 1277
rect 1673 1272 1726 1277
rect 641 1267 646 1272
rect 273 1262 406 1267
rect 457 1262 510 1267
rect 521 1262 646 1267
rect 665 1262 926 1267
rect 977 1262 1006 1267
rect 1089 1262 1126 1267
rect 1953 1262 2054 1267
rect 1953 1257 1958 1262
rect 417 1252 630 1257
rect 705 1252 758 1257
rect 785 1252 870 1257
rect 881 1252 1094 1257
rect 1929 1252 1958 1257
rect 2049 1257 2054 1262
rect 2049 1252 2078 1257
rect 865 1247 870 1252
rect 297 1242 366 1247
rect 401 1242 438 1247
rect 473 1242 646 1247
rect 761 1242 814 1247
rect 865 1242 934 1247
rect 945 1242 1006 1247
rect 1049 1242 1078 1247
rect 1361 1242 1454 1247
rect 1489 1242 1558 1247
rect 1817 1242 1902 1247
rect 1985 1242 2014 1247
rect 2113 1242 2270 1247
rect 2505 1242 2566 1247
rect 1897 1237 1990 1242
rect 249 1232 1286 1237
rect 1465 1232 1526 1237
rect 2025 1232 2150 1237
rect 2409 1232 2502 1237
rect 209 1222 230 1227
rect 289 1222 534 1227
rect 569 1222 718 1227
rect 801 1222 870 1227
rect 897 1222 942 1227
rect 985 1222 1174 1227
rect 1233 1222 1350 1227
rect 1433 1222 1510 1227
rect 1521 1222 1526 1232
rect 1593 1222 1678 1227
rect 1689 1222 1734 1227
rect 1801 1222 1870 1227
rect 1937 1222 1974 1227
rect 2089 1222 2126 1227
rect 2217 1222 2246 1227
rect 2377 1222 2558 1227
rect 2577 1222 2646 1227
rect 121 1212 198 1217
rect 369 1212 470 1217
rect 545 1212 566 1217
rect 593 1212 830 1217
rect 561 1207 566 1212
rect 897 1207 902 1222
rect 1089 1212 1158 1217
rect 1441 1212 1654 1217
rect 2097 1212 2134 1217
rect 2529 1212 2622 1217
rect 185 1202 286 1207
rect 329 1202 350 1207
rect 377 1202 414 1207
rect 433 1202 478 1207
rect 537 1202 566 1207
rect 593 1202 630 1207
rect 681 1202 710 1207
rect 897 1202 926 1207
rect 961 1202 1030 1207
rect 1081 1202 1166 1207
rect 1281 1202 1398 1207
rect 1417 1202 1478 1207
rect 729 1197 878 1202
rect 1393 1197 1398 1202
rect 1473 1197 1478 1202
rect 1561 1202 1590 1207
rect 1817 1202 1926 1207
rect 2049 1202 2118 1207
rect 1561 1197 1566 1202
rect 2129 1197 2134 1212
rect 2177 1202 2238 1207
rect 2457 1202 2566 1207
rect 297 1192 366 1197
rect 449 1192 734 1197
rect 873 1192 1006 1197
rect 1105 1192 1134 1197
rect 1233 1192 1294 1197
rect 1393 1192 1454 1197
rect 1473 1192 1566 1197
rect 1889 1192 1990 1197
rect 2097 1192 2134 1197
rect 2153 1192 2310 1197
rect 2481 1192 2606 1197
rect 1001 1187 1110 1192
rect 105 1182 158 1187
rect 313 1182 710 1187
rect 761 1182 926 1187
rect 937 1182 982 1187
rect 1841 1182 1910 1187
rect 1929 1182 1966 1187
rect 2081 1182 2238 1187
rect 2265 1182 2318 1187
rect 2593 1182 2662 1187
rect 1905 1177 1910 1182
rect 97 1172 150 1177
rect 177 1172 326 1177
rect 337 1172 430 1177
rect 489 1172 550 1177
rect 577 1172 694 1177
rect 713 1172 950 1177
rect 1001 1172 1126 1177
rect 1153 1172 1582 1177
rect 1905 1172 2166 1177
rect 2265 1172 2574 1177
rect 577 1167 582 1172
rect 1001 1167 1006 1172
rect 297 1162 326 1167
rect 441 1162 582 1167
rect 601 1162 622 1167
rect 665 1162 846 1167
rect 953 1162 1006 1167
rect 1121 1167 1126 1172
rect 2161 1167 2270 1172
rect 1121 1162 1150 1167
rect 1881 1162 1990 1167
rect 2081 1162 2142 1167
rect 321 1157 326 1162
rect 1985 1157 2086 1162
rect 81 1152 190 1157
rect 265 1152 310 1157
rect 321 1152 422 1157
rect 529 1152 790 1157
rect 801 1152 1238 1157
rect 1249 1152 1294 1157
rect 1513 1152 1550 1157
rect 1601 1152 1710 1157
rect 1833 1152 1870 1157
rect 305 1147 310 1152
rect 113 1142 142 1147
rect 201 1142 286 1147
rect 305 1142 398 1147
rect 113 1127 118 1142
rect 417 1137 422 1152
rect 465 1142 494 1147
rect 505 1142 566 1147
rect 593 1142 622 1147
rect 633 1142 702 1147
rect 793 1142 878 1147
rect 961 1142 1038 1147
rect 617 1137 622 1142
rect 1233 1137 1238 1152
rect 1601 1147 1606 1152
rect 1257 1142 1358 1147
rect 1433 1142 1518 1147
rect 1537 1142 1606 1147
rect 1705 1147 1710 1152
rect 1865 1147 1870 1152
rect 1937 1152 1966 1157
rect 2105 1152 2246 1157
rect 1937 1147 1942 1152
rect 1705 1142 1734 1147
rect 1865 1142 1942 1147
rect 2057 1142 2094 1147
rect 129 1132 326 1137
rect 417 1132 518 1137
rect 617 1132 662 1137
rect 785 1132 1086 1137
rect 1233 1132 1710 1137
rect 513 1127 598 1132
rect 2089 1127 2094 1142
rect 2225 1142 2254 1147
rect 2225 1127 2230 1142
rect 113 1122 142 1127
rect 153 1122 454 1127
rect 473 1122 494 1127
rect 593 1122 806 1127
rect 913 1122 1006 1127
rect 1129 1122 1206 1127
rect 1273 1122 1462 1127
rect 2089 1122 2230 1127
rect 2289 1122 2358 1127
rect 449 1117 454 1122
rect 1129 1117 1134 1122
rect 345 1112 382 1117
rect 449 1112 774 1117
rect 801 1112 830 1117
rect 849 1112 974 1117
rect 1057 1112 1134 1117
rect 1201 1117 1206 1122
rect 2289 1117 2294 1122
rect 1201 1112 1230 1117
rect 1361 1112 1454 1117
rect 1529 1112 1598 1117
rect 1833 1112 1918 1117
rect 2265 1112 2294 1117
rect 2353 1117 2358 1122
rect 2353 1112 2422 1117
rect 97 1102 134 1107
rect 361 1102 630 1107
rect 697 1102 766 1107
rect 841 1102 1046 1107
rect 1249 1102 1342 1107
rect 1577 1102 1718 1107
rect 1065 1097 1254 1102
rect 1337 1097 1342 1102
rect 89 1092 430 1097
rect 465 1092 502 1097
rect 545 1092 590 1097
rect 601 1092 630 1097
rect 657 1092 1070 1097
rect 1337 1092 1398 1097
rect 2281 1092 2342 1097
rect 337 1082 678 1087
rect 689 1082 1390 1087
rect 1521 1082 1694 1087
rect 217 1077 318 1082
rect 161 1072 222 1077
rect 313 1072 414 1077
rect 433 1072 606 1077
rect 753 1072 814 1077
rect 889 1072 1038 1077
rect 1129 1072 1350 1077
rect 625 1067 734 1072
rect 1345 1067 1350 1072
rect 1409 1072 1510 1077
rect 1409 1067 1414 1072
rect 185 1062 302 1067
rect 401 1062 630 1067
rect 729 1062 1270 1067
rect 1345 1062 1414 1067
rect 1505 1067 1510 1072
rect 1705 1072 1790 1077
rect 1505 1062 1582 1067
rect 297 1057 406 1062
rect 1577 1057 1582 1062
rect 1705 1057 1710 1072
rect 1921 1062 1958 1067
rect 233 1052 278 1057
rect 425 1052 454 1057
rect 505 1052 558 1057
rect 585 1052 662 1057
rect 689 1052 982 1057
rect 1001 1052 1326 1057
rect 1577 1052 1710 1057
rect 1825 1052 1902 1057
rect 1825 1047 1830 1052
rect 17 1042 110 1047
rect 177 1042 230 1047
rect 289 1042 334 1047
rect 353 1042 550 1047
rect 561 1042 678 1047
rect 777 1042 950 1047
rect 985 1042 1046 1047
rect 1057 1042 1310 1047
rect 1801 1042 1830 1047
rect 1897 1047 1902 1052
rect 1897 1042 1926 1047
rect 17 877 22 1042
rect 1057 1037 1062 1042
rect 65 1032 302 1037
rect 321 1032 518 1037
rect 569 1032 622 1037
rect 633 1032 790 1037
rect 801 1032 862 1037
rect 897 1032 942 1037
rect 993 1032 1062 1037
rect 1073 1032 1422 1037
rect 1489 1032 1558 1037
rect 1817 1032 1886 1037
rect 2049 1032 2094 1037
rect 513 1027 518 1032
rect 993 1027 998 1032
rect 313 1022 446 1027
rect 473 1022 502 1027
rect 513 1022 998 1027
rect 1009 1022 1126 1027
rect 1145 1022 1182 1027
rect 1273 1022 1350 1027
rect 1481 1022 1606 1027
rect 1705 1022 1982 1027
rect 2017 1022 2150 1027
rect 2161 1022 2286 1027
rect 2561 1022 2622 1027
rect 209 1017 294 1022
rect 497 1017 502 1022
rect 65 1012 214 1017
rect 289 1012 350 1017
rect 369 1007 374 1017
rect 225 1002 286 1007
rect 305 1002 374 1007
rect 385 1007 390 1017
rect 425 1012 486 1017
rect 497 1012 518 1017
rect 553 1012 670 1017
rect 721 1012 766 1017
rect 881 1012 934 1017
rect 945 1012 1014 1017
rect 1113 1012 1262 1017
rect 385 1002 438 1007
rect 481 1002 486 1012
rect 945 1007 950 1012
rect 1009 1007 1014 1012
rect 1257 1007 1262 1012
rect 1345 1012 1462 1017
rect 2481 1012 2582 1017
rect 1345 1007 1350 1012
rect 1481 1007 1950 1012
rect 529 1002 550 1007
rect 625 1002 686 1007
rect 849 1002 902 1007
rect 921 1002 950 1007
rect 961 1002 998 1007
rect 1009 1002 1086 1007
rect 225 992 230 1002
rect 545 997 550 1002
rect 1121 997 1126 1007
rect 1257 1002 1350 1007
rect 1369 1002 1486 1007
rect 1945 1002 2166 1007
rect 273 992 526 997
rect 545 992 582 997
rect 593 992 830 997
rect 857 992 918 997
rect 937 992 1022 997
rect 1057 992 1190 997
rect 1489 992 1550 997
rect 1569 992 1790 997
rect 1801 992 1982 997
rect 2161 992 2166 1002
rect 1785 987 1790 992
rect 81 982 134 987
rect 209 982 270 987
rect 297 982 430 987
rect 577 982 606 987
rect 617 982 638 987
rect 673 982 862 987
rect 881 982 926 987
rect 969 982 1150 987
rect 1313 982 1774 987
rect 1785 982 2070 987
rect 2441 982 2598 987
rect 881 977 886 982
rect 201 972 254 977
rect 281 972 486 977
rect 537 972 702 977
rect 753 972 814 977
rect 825 972 854 977
rect 865 972 886 977
rect 929 972 982 977
rect 1105 972 1182 977
rect 1225 972 1350 977
rect 1481 972 1534 977
rect 1721 972 1822 977
rect 1937 972 2038 977
rect 33 962 166 967
rect 257 962 390 967
rect 425 962 702 967
rect 737 962 1086 967
rect 33 907 38 962
rect 1345 957 1350 972
rect 1553 967 1702 972
rect 1937 967 1942 972
rect 2385 967 2478 972
rect 1521 962 1558 967
rect 1697 962 1814 967
rect 1841 962 1942 967
rect 1953 962 2326 967
rect 2361 962 2390 967
rect 2473 962 2502 967
rect 49 952 94 957
rect 185 952 246 957
rect 257 952 310 957
rect 377 952 934 957
rect 945 952 1014 957
rect 1257 952 1326 957
rect 1345 952 1366 957
rect 1409 952 1478 957
rect 49 917 54 952
rect 929 947 934 952
rect 1521 947 1526 962
rect 1553 952 1654 957
rect 1681 952 2006 957
rect 2393 952 2494 957
rect 2593 952 2614 957
rect 1681 947 1686 952
rect 289 942 406 947
rect 417 942 494 947
rect 505 942 534 947
rect 321 932 358 937
rect 73 922 134 927
rect 145 922 206 927
rect 225 922 342 927
rect 361 922 382 927
rect 417 922 422 942
rect 529 937 534 942
rect 449 932 486 937
rect 529 932 566 937
rect 481 922 486 932
rect 641 927 646 947
rect 729 937 734 947
rect 777 942 822 947
rect 841 942 910 947
rect 929 942 950 947
rect 961 942 1118 947
rect 1345 942 1526 947
rect 1537 942 1606 947
rect 1633 942 1686 947
rect 1705 942 1734 947
rect 945 937 950 942
rect 1345 937 1350 942
rect 729 932 798 937
rect 817 932 894 937
rect 641 922 686 927
rect 769 922 774 932
rect 929 927 934 937
rect 945 932 1142 937
rect 1153 932 1350 937
rect 1361 932 1622 937
rect 1633 932 1638 942
rect 1729 937 1734 942
rect 1649 932 1694 937
rect 1713 932 1734 937
rect 1809 942 1830 947
rect 1929 942 1958 947
rect 2017 942 2094 947
rect 2297 942 2326 947
rect 2409 942 2510 947
rect 2561 942 2654 947
rect 801 922 934 927
rect 969 922 1046 927
rect 1089 922 1126 927
rect 49 912 110 917
rect 121 912 214 917
rect 297 912 446 917
rect 457 912 566 917
rect 601 912 766 917
rect 841 912 958 917
rect 985 912 1054 917
rect 1137 907 1142 932
rect 1193 922 1230 927
rect 1225 917 1230 922
rect 1321 922 1350 927
rect 1361 922 1366 932
rect 1713 927 1718 932
rect 1393 922 1678 927
rect 1697 922 1718 927
rect 1321 917 1326 922
rect 1225 912 1326 917
rect 1345 907 1350 922
rect 1809 917 1814 942
rect 1897 932 1998 937
rect 2009 932 2054 937
rect 2145 932 2286 937
rect 2345 932 2390 937
rect 2401 932 2454 937
rect 2601 932 2630 937
rect 2385 927 2390 932
rect 2449 927 2606 932
rect 1841 922 1862 927
rect 2273 922 2374 927
rect 2385 922 2430 927
rect 2369 917 2374 922
rect 1457 912 1558 917
rect 1569 912 1678 917
rect 1689 912 1790 917
rect 1809 912 1838 917
rect 1865 912 1942 917
rect 2041 912 2150 917
rect 2369 912 2454 917
rect 2473 912 2566 917
rect 33 902 62 907
rect 193 902 270 907
rect 305 902 342 907
rect 393 902 534 907
rect 545 902 582 907
rect 593 902 622 907
rect 649 902 678 907
rect 721 902 934 907
rect 945 902 1102 907
rect 1137 902 1206 907
rect 1345 902 1502 907
rect 57 897 198 902
rect 217 892 518 897
rect 561 892 614 897
rect 625 892 670 897
rect 705 892 758 897
rect 785 892 830 897
rect 865 892 886 897
rect 897 892 1038 897
rect 1497 892 1526 897
rect 1553 892 1558 912
rect 1577 902 1670 907
rect 1681 902 1710 907
rect 1721 902 1894 907
rect 2449 897 2454 912
rect 2521 902 2550 907
rect 2521 897 2526 902
rect 1713 892 1782 897
rect 1929 892 1958 897
rect 2449 892 2526 897
rect 1329 887 1422 892
rect 1553 887 1694 892
rect 145 882 278 887
rect 353 882 926 887
rect 937 882 982 887
rect 1089 882 1278 887
rect 1305 882 1334 887
rect 1417 882 1446 887
rect 1481 882 1542 887
rect 1689 882 1806 887
rect 1817 882 1878 887
rect 145 877 150 882
rect 1089 877 1094 882
rect 17 872 150 877
rect 249 872 510 877
rect 585 872 718 877
rect 929 872 966 877
rect 1065 872 1094 877
rect 1273 877 1278 882
rect 1273 872 1750 877
rect 1769 872 1998 877
rect 737 867 910 872
rect 1129 867 1238 872
rect 233 862 462 867
rect 497 862 646 867
rect 681 862 742 867
rect 905 862 1006 867
rect 1105 862 1134 867
rect 1233 862 1262 867
rect 1385 862 1478 867
rect 1577 862 1606 867
rect 1753 862 1950 867
rect 1473 857 1582 862
rect 1641 857 1734 862
rect 169 852 398 857
rect 409 852 654 857
rect 689 852 758 857
rect 769 852 910 857
rect 1009 852 1294 857
rect 1409 852 1454 857
rect 1617 852 1646 857
rect 1729 852 1870 857
rect 1409 847 1414 852
rect 137 842 1022 847
rect 1089 842 1166 847
rect 1257 842 1414 847
rect 1425 842 1518 847
rect 1657 842 1774 847
rect 1809 842 1886 847
rect 1921 842 2006 847
rect 2017 842 2182 847
rect 2361 842 2494 847
rect 2553 842 2622 847
rect 2553 837 2558 842
rect 241 832 382 837
rect 441 832 534 837
rect 569 832 734 837
rect 777 832 838 837
rect 873 832 894 837
rect 953 832 1030 837
rect 1049 832 1102 837
rect 1137 832 1334 837
rect 1393 832 1510 837
rect 1553 832 1646 837
rect 1705 832 1878 837
rect 1937 832 1990 837
rect 2313 832 2358 837
rect 2529 832 2558 837
rect 2617 837 2622 842
rect 2617 832 2646 837
rect 249 822 366 827
rect 457 822 702 827
rect 713 822 846 827
rect 873 822 926 827
rect 1049 822 1142 827
rect 1169 822 1198 827
rect 1481 822 1526 827
rect 1577 822 1670 827
rect 1681 822 1742 827
rect 1793 822 1862 827
rect 1881 822 1934 827
rect 1977 822 2070 827
rect 2145 822 2174 827
rect 2417 822 2462 827
rect 361 817 462 822
rect 225 812 286 817
rect 305 812 342 817
rect 481 812 974 817
rect 993 812 1014 817
rect 1073 812 1118 817
rect 1137 812 1142 822
rect 1681 817 1686 822
rect 1857 817 1862 822
rect 1185 812 1342 817
rect 1433 812 1686 817
rect 1769 812 1822 817
rect 1857 812 1918 817
rect 1985 812 2014 817
rect 2161 812 2254 817
rect 2409 812 2470 817
rect 2537 812 2638 817
rect 281 807 286 812
rect 993 807 998 812
rect 1185 807 1190 812
rect 1985 807 1990 812
rect 281 802 302 807
rect 345 802 390 807
rect 425 802 470 807
rect 505 802 614 807
rect 641 802 798 807
rect 849 802 918 807
rect 929 802 998 807
rect 1009 802 1190 807
rect 1209 802 1262 807
rect 1369 802 1470 807
rect 1505 802 1598 807
rect 1609 802 1630 807
rect 1641 802 1678 807
rect 1849 802 1990 807
rect 2009 802 2126 807
rect 2353 802 2382 807
rect 2449 802 2534 807
rect 2617 802 2662 807
rect 641 797 646 802
rect 929 797 934 802
rect 97 792 134 797
rect 273 792 558 797
rect 625 792 646 797
rect 713 792 934 797
rect 1025 792 1094 797
rect 1201 792 1414 797
rect 1441 792 1494 797
rect 1025 787 1030 792
rect 1505 787 1510 802
rect 1609 797 1614 802
rect 2353 797 2358 802
rect 1521 792 1630 797
rect 105 782 190 787
rect 281 782 422 787
rect 433 782 486 787
rect 497 782 550 787
rect 593 782 654 787
rect 737 782 1030 787
rect 1041 782 1366 787
rect 1393 782 1510 787
rect 1625 787 1630 792
rect 1689 792 1774 797
rect 1785 792 2030 797
rect 2209 792 2238 797
rect 2321 792 2358 797
rect 2497 792 2638 797
rect 1689 787 1694 792
rect 1625 782 1694 787
rect 1713 782 1766 787
rect 1793 782 1990 787
rect 2241 777 2326 782
rect 369 772 638 777
rect 665 772 1310 777
rect 1393 772 1462 777
rect 1505 772 1558 777
rect 1737 772 1790 777
rect 1857 772 1966 777
rect 2145 772 2246 777
rect 2321 772 2374 777
rect 2369 767 2374 772
rect 313 762 438 767
rect 513 762 694 767
rect 777 762 806 767
rect 849 762 1006 767
rect 1025 762 1062 767
rect 1097 762 1150 767
rect 1497 762 1782 767
rect 2257 762 2326 767
rect 2369 762 2478 767
rect 1025 757 1030 762
rect 1849 757 1950 762
rect 265 752 502 757
rect 537 752 622 757
rect 633 752 1030 757
rect 1097 752 1326 757
rect 1385 752 1478 757
rect 1825 752 1854 757
rect 1945 752 1974 757
rect 1385 747 1390 752
rect 1473 747 1550 752
rect 193 742 254 747
rect 401 742 622 747
rect 705 742 742 747
rect 769 742 934 747
rect 985 742 1038 747
rect 1073 742 1390 747
rect 1545 742 1662 747
rect 1777 742 1806 747
rect 249 737 406 742
rect 617 737 710 742
rect 1825 737 1830 752
rect 1889 742 1934 747
rect 1945 742 2054 747
rect 2209 742 2294 747
rect 2425 742 2510 747
rect 2529 742 2574 747
rect 2593 742 2670 747
rect 2425 737 2430 742
rect 521 732 598 737
rect 729 732 1278 737
rect 1401 732 1534 737
rect 1713 732 1830 737
rect 1841 732 1998 737
rect 2401 732 2430 737
rect 2505 737 2510 742
rect 2505 732 2550 737
rect 425 727 502 732
rect 129 722 182 727
rect 177 717 182 722
rect 281 722 430 727
rect 497 722 1086 727
rect 1113 722 1262 727
rect 1321 722 1686 727
rect 1697 722 1878 727
rect 2433 722 2470 727
rect 2529 722 2614 727
rect 281 717 286 722
rect 1681 717 1686 722
rect 2433 717 2438 722
rect 177 712 286 717
rect 441 712 550 717
rect 561 712 926 717
rect 945 712 1046 717
rect 1089 712 1198 717
rect 1217 712 1302 717
rect 1313 712 1574 717
rect 1681 712 1974 717
rect 2217 712 2438 717
rect 2457 712 2486 717
rect 561 707 566 712
rect 1569 707 1662 712
rect 321 702 566 707
rect 593 702 1174 707
rect 1281 702 1350 707
rect 1401 702 1550 707
rect 1657 702 1838 707
rect 2449 702 2550 707
rect 1169 697 1270 702
rect 305 692 558 697
rect 625 692 806 697
rect 817 692 886 697
rect 929 692 1014 697
rect 1041 692 1150 697
rect 1265 692 1366 697
rect 1481 692 1526 697
rect 1553 692 1670 697
rect 1721 692 1870 697
rect 2161 692 2206 697
rect 881 687 886 692
rect 1361 687 1438 692
rect 2201 687 2206 692
rect 2265 692 2294 697
rect 2265 687 2270 692
rect 265 682 294 687
rect 289 677 294 682
rect 425 682 590 687
rect 689 682 742 687
rect 785 682 846 687
rect 881 682 998 687
rect 1025 682 1318 687
rect 1433 682 1534 687
rect 1545 682 1814 687
rect 2201 682 2270 687
rect 425 677 430 682
rect 289 672 430 677
rect 585 672 918 677
rect 969 672 1102 677
rect 1137 672 1198 677
rect 1361 672 1422 677
rect 1497 672 1566 677
rect 1785 672 1902 677
rect 473 667 566 672
rect 1681 667 1766 672
rect 449 662 478 667
rect 561 662 606 667
rect 625 662 662 667
rect 761 662 790 667
rect 873 662 910 667
rect 961 662 1254 667
rect 1297 662 1326 667
rect 1401 662 1686 667
rect 1761 662 1822 667
rect 1841 662 1894 667
rect 1841 657 1846 662
rect 513 652 870 657
rect 881 652 1038 657
rect 1185 652 1542 657
rect 1697 652 1726 657
rect 1753 652 1846 657
rect 1857 652 1966 657
rect 2249 652 2494 657
rect 409 642 614 647
rect 761 642 814 647
rect 849 642 910 647
rect 961 642 1126 647
rect 1169 642 1238 647
rect 1305 642 1382 647
rect 1393 642 1422 647
rect 1633 642 1710 647
rect 1761 642 1982 647
rect 2129 642 2278 647
rect 633 637 742 642
rect 401 632 462 637
rect 489 632 558 637
rect 593 632 638 637
rect 737 632 886 637
rect 897 632 950 637
rect 993 632 1046 637
rect 1057 632 1158 637
rect 1329 632 1454 637
rect 1473 632 1590 637
rect 1609 632 1814 637
rect 1953 632 1998 637
rect 2017 632 2094 637
rect 2193 632 2254 637
rect 881 627 886 632
rect 1473 627 1478 632
rect 281 622 326 627
rect 433 622 510 627
rect 537 622 638 627
rect 681 622 726 627
rect 793 622 854 627
rect 881 622 926 627
rect 1017 622 1150 627
rect 1281 622 1478 627
rect 1585 627 1590 632
rect 2017 627 2022 632
rect 1585 622 2022 627
rect 2089 627 2094 632
rect 2089 622 2118 627
rect 2177 622 2198 627
rect 2217 622 2270 627
rect 2473 622 2614 627
rect 385 612 550 617
rect 713 612 902 617
rect 945 612 1030 617
rect 1041 612 1270 617
rect 1289 612 1342 617
rect 1353 612 1374 617
rect 1441 612 1782 617
rect 1817 612 1918 617
rect 2105 612 2214 617
rect 385 607 390 612
rect 297 602 390 607
rect 409 602 478 607
rect 489 602 534 607
rect 641 602 694 607
rect 745 602 774 607
rect 865 602 894 607
rect 945 597 950 612
rect 1265 607 1270 612
rect 985 602 1022 607
rect 1089 602 1222 607
rect 1265 602 1606 607
rect 1641 602 1686 607
rect 1761 602 1830 607
rect 1977 602 2046 607
rect 2377 602 2518 607
rect 1217 597 1222 602
rect 233 592 294 597
rect 345 592 814 597
rect 897 592 950 597
rect 969 592 1014 597
rect 1057 592 1174 597
rect 1217 592 1326 597
rect 1393 592 1510 597
rect 1529 592 1702 597
rect 1721 592 1766 597
rect 1785 592 1870 597
rect 1929 592 2094 597
rect 2105 592 2182 597
rect 897 587 902 592
rect 1057 587 1062 592
rect 1761 587 1766 592
rect 393 582 542 587
rect 577 582 662 587
rect 721 582 902 587
rect 921 582 1062 587
rect 1073 582 1158 587
rect 1169 582 1214 587
rect 1329 582 1422 587
rect 1449 582 1486 587
rect 1569 582 1622 587
rect 1665 582 1742 587
rect 1761 582 1894 587
rect 1985 582 2158 587
rect 2233 582 2326 587
rect 1073 577 1078 582
rect 273 572 614 577
rect 713 572 966 577
rect 1025 572 1078 577
rect 1097 572 1390 577
rect 609 567 718 572
rect 961 567 966 572
rect 1417 567 1422 577
rect 1433 572 1734 577
rect 1785 572 1878 577
rect 2337 572 2446 577
rect 185 562 590 567
rect 753 562 846 567
rect 961 562 998 567
rect 1065 562 1358 567
rect 1417 562 1566 567
rect 1649 562 1742 567
rect 225 552 326 557
rect 361 552 406 557
rect 465 552 534 557
rect 657 552 718 557
rect 809 552 942 557
rect 969 552 1014 557
rect 1065 552 1214 557
rect 1249 552 1302 557
rect 1345 552 1422 557
rect 1433 552 1470 557
rect 1481 552 1550 557
rect 1009 547 1014 552
rect 1417 547 1422 552
rect 665 542 710 547
rect 897 542 990 547
rect 1009 542 1102 547
rect 1113 542 1190 547
rect 1281 542 1406 547
rect 1417 542 1558 547
rect 1649 537 1654 562
rect 1737 557 1742 562
rect 1889 562 2102 567
rect 1889 557 1894 562
rect 1673 552 1718 557
rect 1737 552 1894 557
rect 2433 552 2470 557
rect 2025 542 2134 547
rect 2489 542 2590 547
rect 297 532 390 537
rect 497 532 558 537
rect 601 532 630 537
rect 785 532 1222 537
rect 1241 532 1270 537
rect 1369 532 1518 537
rect 1569 532 1654 537
rect 1721 532 1838 537
rect 1857 532 1910 537
rect 561 522 686 527
rect 945 522 1046 527
rect 1057 522 1206 527
rect 945 517 950 522
rect 1041 517 1046 522
rect 305 512 350 517
rect 449 512 606 517
rect 697 512 950 517
rect 961 512 1022 517
rect 1041 512 1166 517
rect 601 507 702 512
rect 1217 507 1222 532
rect 1265 527 1270 532
rect 1857 527 1862 532
rect 1265 522 1294 527
rect 1377 522 1422 527
rect 1433 522 1622 527
rect 1825 522 1862 527
rect 1641 517 1830 522
rect 1977 517 1982 537
rect 2121 532 2182 537
rect 1273 512 1526 517
rect 1577 512 1646 517
rect 1881 512 1950 517
rect 1977 512 1990 517
rect 2001 512 2078 517
rect 329 502 550 507
rect 721 502 1086 507
rect 1217 502 1310 507
rect 1321 502 1430 507
rect 1457 502 1806 507
rect 1825 502 1902 507
rect 1985 502 1990 512
rect 625 492 694 497
rect 841 492 1350 497
rect 1401 492 1502 497
rect 1513 492 1654 497
rect 1753 492 1814 497
rect 1889 492 2030 497
rect 1513 487 1518 492
rect 1649 487 1758 492
rect 521 482 558 487
rect 713 482 822 487
rect 881 482 1134 487
rect 1225 482 1518 487
rect 1777 482 1910 487
rect 577 477 718 482
rect 817 477 822 482
rect 1537 477 1630 482
rect 65 472 582 477
rect 817 472 870 477
rect 937 472 1054 477
rect 1065 472 1286 477
rect 1433 472 1542 477
rect 1625 472 1710 477
rect 1281 467 1286 472
rect 1705 467 1710 472
rect 1801 472 1830 477
rect 1841 472 2014 477
rect 1801 467 1806 472
rect 577 462 1254 467
rect 1281 462 1382 467
rect 1393 462 1494 467
rect 1553 462 1614 467
rect 1705 462 1806 467
rect 1857 462 2142 467
rect 1377 457 1382 462
rect 665 452 1262 457
rect 1377 452 1462 457
rect 1585 452 1686 457
rect 2017 452 2078 457
rect 449 442 486 447
rect 537 442 670 447
rect 689 442 1086 447
rect 1105 442 1582 447
rect 1617 442 1654 447
rect 1841 442 2014 447
rect 1105 437 1110 442
rect 537 432 630 437
rect 657 432 710 437
rect 801 432 854 437
rect 865 432 1110 437
rect 1137 432 1390 437
rect 1425 432 1454 437
rect 1569 432 1646 437
rect 1841 427 1846 442
rect 1961 432 2030 437
rect 289 417 294 427
rect 489 422 638 427
rect 785 422 1102 427
rect 1233 422 1270 427
rect 1305 422 1622 427
rect 1633 417 1638 427
rect 1785 422 1846 427
rect 1929 422 1958 427
rect 1953 417 1958 422
rect 2561 422 2614 427
rect 2561 417 2566 422
rect 289 412 358 417
rect 369 412 550 417
rect 673 412 1262 417
rect 1377 412 1486 417
rect 1497 412 1638 417
rect 1785 412 1846 417
rect 1873 412 1926 417
rect 1953 412 1998 417
rect 2273 412 2422 417
rect 2441 412 2566 417
rect 2417 407 2422 412
rect 457 402 534 407
rect 713 402 750 407
rect 913 402 982 407
rect 993 402 1062 407
rect 1081 402 1254 407
rect 1457 402 1526 407
rect 1729 402 1774 407
rect 1977 402 2006 407
rect 2417 402 2486 407
rect 913 397 918 402
rect 1545 397 1614 402
rect 1729 397 1734 402
rect 177 392 246 397
rect 329 392 382 397
rect 409 392 438 397
rect 433 387 438 392
rect 529 392 558 397
rect 657 392 782 397
rect 793 392 918 397
rect 929 392 1006 397
rect 1041 392 1078 397
rect 1169 392 1334 397
rect 1417 392 1550 397
rect 1609 392 1734 397
rect 1897 392 2022 397
rect 2137 392 2230 397
rect 2249 392 2334 397
rect 529 387 534 392
rect 1169 387 1174 392
rect 2225 387 2230 392
rect 281 382 342 387
rect 433 382 534 387
rect 601 382 630 387
rect 681 382 726 387
rect 761 382 1174 387
rect 1337 382 1430 387
rect 1505 382 1598 387
rect 1833 382 1934 387
rect 2009 382 2086 387
rect 2225 382 2590 387
rect 1217 377 1318 382
rect 785 372 1222 377
rect 1313 372 1366 377
rect 1513 372 1566 377
rect 1641 372 1742 377
rect 1881 372 1942 377
rect 2313 372 2366 377
rect 729 362 1334 367
rect 1353 362 1382 367
rect 1569 362 1662 367
rect 1777 362 1878 367
rect 1905 362 1926 367
rect 1953 362 2030 367
rect 1473 357 1574 362
rect 1953 357 1958 362
rect 225 352 326 357
rect 393 352 462 357
rect 641 352 710 357
rect 865 352 934 357
rect 977 352 1054 357
rect 1073 352 1166 357
rect 1209 352 1254 357
rect 1393 352 1478 357
rect 1585 352 1806 357
rect 1913 352 1958 357
rect 2369 352 2510 357
rect 729 347 846 352
rect 297 342 382 347
rect 377 337 382 342
rect 441 342 470 347
rect 593 342 734 347
rect 841 342 1022 347
rect 1369 342 1430 347
rect 1481 342 1622 347
rect 1809 342 1950 347
rect 1993 342 2070 347
rect 2185 342 2302 347
rect 2449 342 2478 347
rect 441 337 446 342
rect 2449 337 2454 342
rect 305 332 350 337
rect 377 332 446 337
rect 521 332 838 337
rect 897 332 982 337
rect 1241 332 1310 337
rect 1321 332 1446 337
rect 1497 332 1550 337
rect 1561 332 1686 337
rect 1921 332 1990 337
rect 2345 332 2454 337
rect 2465 332 2574 337
rect 481 322 534 327
rect 657 322 758 327
rect 857 322 902 327
rect 969 322 1038 327
rect 1241 322 1270 327
rect 1337 322 1406 327
rect 1425 322 1478 327
rect 1833 322 1886 327
rect 2265 322 2294 327
rect 2329 322 2382 327
rect 2457 322 2638 327
rect 753 317 758 322
rect 449 312 502 317
rect 753 312 838 317
rect 977 312 1014 317
rect 1121 312 1190 317
rect 1297 312 1358 317
rect 1673 312 1750 317
rect 1761 312 1814 317
rect 1961 312 2006 317
rect 2017 312 2126 317
rect 2257 312 2374 317
rect 2473 312 2534 317
rect 2545 312 2622 317
rect 633 307 734 312
rect 273 302 350 307
rect 505 302 638 307
rect 729 302 1006 307
rect 1025 302 1078 307
rect 1281 302 1406 307
rect 1417 302 1454 307
rect 1649 302 1710 307
rect 1985 302 2030 307
rect 2241 302 2446 307
rect 2537 302 2566 307
rect 649 292 878 297
rect 985 292 1030 297
rect 1057 292 1142 297
rect 1465 292 1510 297
rect 1609 292 1646 297
rect 1657 292 1702 297
rect 2329 292 2670 297
rect 529 282 630 287
rect 729 282 782 287
rect 801 282 1094 287
rect 1177 282 1638 287
rect 1729 282 1806 287
rect 2281 282 2382 287
rect 529 277 534 282
rect 625 277 710 282
rect 393 272 534 277
rect 705 272 734 277
rect 761 272 830 277
rect 889 272 1070 277
rect 1089 272 1094 282
rect 1729 277 1734 282
rect 1689 272 1734 277
rect 1801 277 1806 282
rect 2377 277 2382 282
rect 2465 282 2494 287
rect 2465 277 2470 282
rect 1801 272 2014 277
rect 2161 272 2270 277
rect 1089 267 1214 272
rect 1505 267 1582 272
rect 2265 267 2270 272
rect 2329 272 2358 277
rect 2377 272 2470 277
rect 2329 267 2334 272
rect 545 262 750 267
rect 977 262 1014 267
rect 1209 262 1262 267
rect 1305 262 1390 267
rect 1481 262 1510 267
rect 1577 262 1678 267
rect 1305 257 1310 262
rect 689 252 838 257
rect 961 252 1214 257
rect 1281 252 1310 257
rect 1385 257 1390 262
rect 1673 257 1678 262
rect 1745 262 1790 267
rect 2265 262 2334 267
rect 1745 257 1750 262
rect 1385 252 1470 257
rect 689 247 694 252
rect 1465 247 1470 252
rect 1537 252 1566 257
rect 1673 252 1750 257
rect 1537 247 1542 252
rect 369 242 694 247
rect 761 242 1078 247
rect 1225 242 1438 247
rect 1465 242 1542 247
rect 1601 242 1622 247
rect 2377 242 2430 247
rect 1073 237 1166 242
rect 1225 237 1230 242
rect 721 232 774 237
rect 809 232 870 237
rect 1017 232 1054 237
rect 1161 232 1230 237
rect 1289 232 1334 237
rect 1601 232 1606 242
rect 1625 232 1702 237
rect 1785 232 1966 237
rect 2129 232 2238 237
rect 2257 232 2310 237
rect 2521 232 2558 237
rect 449 222 550 227
rect 705 222 806 227
rect 817 222 910 227
rect 921 222 1022 227
rect 1041 222 1142 227
rect 1321 222 1766 227
rect 545 217 550 222
rect 801 217 806 222
rect 361 212 414 217
rect 545 212 574 217
rect 801 212 854 217
rect 905 212 990 217
rect 289 202 358 207
rect 385 202 534 207
rect 689 202 742 207
rect 1017 202 1046 207
rect 441 192 462 197
rect 577 192 838 197
rect 913 192 998 197
rect 913 187 918 192
rect 393 182 918 187
rect 993 187 998 192
rect 1025 192 1062 197
rect 1025 187 1030 192
rect 1073 187 1078 222
rect 1785 217 1790 232
rect 1177 212 1302 217
rect 1609 212 1790 217
rect 1961 217 1966 232
rect 2417 222 2486 227
rect 2513 222 2574 227
rect 2417 217 2422 222
rect 1961 212 2070 217
rect 2201 212 2270 217
rect 2313 212 2422 217
rect 2457 212 2494 217
rect 1401 207 1590 212
rect 1137 202 1278 207
rect 1377 202 1406 207
rect 1585 202 1686 207
rect 1705 202 1758 207
rect 1769 202 1806 207
rect 1817 202 1982 207
rect 1249 192 1438 197
rect 1489 192 1862 197
rect 2209 192 2326 197
rect 2553 192 2614 197
rect 1489 187 1494 192
rect 993 182 1030 187
rect 1049 182 1134 187
rect 1361 182 1494 187
rect 1577 182 1718 187
rect 1785 182 1806 187
rect 2289 182 2470 187
rect 1713 177 1718 182
rect 345 172 726 177
rect 721 167 726 172
rect 929 172 1150 177
rect 1177 172 1374 177
rect 929 167 934 172
rect 1369 167 1374 172
rect 1513 172 1614 177
rect 1673 172 1702 177
rect 1713 172 1950 177
rect 1513 167 1518 172
rect 265 162 334 167
rect 329 157 334 162
rect 401 162 478 167
rect 569 162 702 167
rect 721 162 934 167
rect 1065 162 1142 167
rect 1369 162 1518 167
rect 1777 162 1846 167
rect 401 157 406 162
rect 473 157 574 162
rect 1561 157 1670 162
rect 329 152 406 157
rect 593 152 646 157
rect 1025 152 1350 157
rect 1537 152 1566 157
rect 1665 152 1694 157
rect 241 142 270 147
rect 265 137 270 142
rect 425 142 470 147
rect 489 142 534 147
rect 561 142 870 147
rect 961 142 1158 147
rect 425 137 430 142
rect 265 132 430 137
rect 465 107 470 142
rect 1537 137 1542 152
rect 1561 142 1590 147
rect 537 132 566 137
rect 561 127 566 132
rect 881 132 1542 137
rect 1585 137 1590 142
rect 1649 142 1766 147
rect 1649 137 1654 142
rect 1585 132 1654 137
rect 1761 137 1766 142
rect 1857 142 2046 147
rect 1857 137 1862 142
rect 1761 132 1862 137
rect 881 127 886 132
rect 561 122 886 127
rect 937 122 966 127
rect 1001 122 1030 127
rect 937 107 942 122
rect 1025 117 1030 122
rect 1161 122 1190 127
rect 1265 122 1366 127
rect 1161 117 1166 122
rect 1025 112 1166 117
rect 465 102 942 107
rect 889 72 1246 77
use AND2X2  AND2X2_0
timestamp 1710899220
transform 1 0 272 0 1 2170
box -8 -3 40 105
use AND2X2  AND2X2_1
timestamp 1710899220
transform 1 0 384 0 1 2170
box -8 -3 40 105
use AND2X2  AND2X2_2
timestamp 1710899220
transform 1 0 488 0 1 2170
box -8 -3 40 105
use AND2X2  AND2X2_3
timestamp 1710899220
transform 1 0 1288 0 -1 2170
box -8 -3 40 105
use AND2X2  AND2X2_4
timestamp 1710899220
transform 1 0 216 0 -1 1370
box -8 -3 40 105
use AND2X2  AND2X2_5
timestamp 1710899220
transform 1 0 96 0 1 770
box -8 -3 40 105
use AND2X2  AND2X2_6
timestamp 1710899220
transform 1 0 1184 0 1 770
box -8 -3 40 105
use AND2X2  AND2X2_7
timestamp 1710899220
transform 1 0 168 0 1 2170
box -8 -3 40 105
use AND2X2  AND2X2_8
timestamp 1710899220
transform 1 0 2016 0 1 1170
box -8 -3 40 105
use AND2X2  AND2X2_9
timestamp 1710899220
transform 1 0 2032 0 -1 1570
box -8 -3 40 105
use AND2X2  AND2X2_10
timestamp 1710899220
transform 1 0 2216 0 -1 1570
box -8 -3 40 105
use AND2X2  AND2X2_11
timestamp 1710899220
transform 1 0 2192 0 -1 1770
box -8 -3 40 105
use AND2X2  AND2X2_12
timestamp 1710899220
transform 1 0 2000 0 1 1770
box -8 -3 40 105
use AND2X2  AND2X2_13
timestamp 1710899220
transform 1 0 1984 0 -1 1770
box -8 -3 40 105
use AND2X2  AND2X2_14
timestamp 1710899220
transform 1 0 2192 0 1 570
box -8 -3 40 105
use AND2X2  AND2X2_15
timestamp 1710899220
transform 1 0 1256 0 1 370
box -8 -3 40 105
use AND2X2  AND2X2_16
timestamp 1710899220
transform 1 0 856 0 1 1170
box -8 -3 40 105
use AND2X2  AND2X2_17
timestamp 1710899220
transform 1 0 2248 0 1 170
box -8 -3 40 105
use AND2X2  AND2X2_18
timestamp 1710899220
transform 1 0 2592 0 -1 770
box -8 -3 40 105
use AND2X2  AND2X2_19
timestamp 1710899220
transform 1 0 2352 0 1 770
box -8 -3 40 105
use AOI21X1  AOI21X1_0
timestamp 1710899220
transform 1 0 512 0 -1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_1
timestamp 1710899220
transform 1 0 1608 0 -1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_2
timestamp 1710899220
transform 1 0 2008 0 1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_3
timestamp 1710899220
transform 1 0 1976 0 1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_4
timestamp 1710899220
transform 1 0 1784 0 1 570
box -7 -3 39 105
use AOI21X1  AOI21X1_5
timestamp 1710899220
transform 1 0 512 0 1 570
box -7 -3 39 105
use AOI21X1  AOI21X1_6
timestamp 1710899220
transform 1 0 1592 0 -1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_7
timestamp 1710899220
transform 1 0 776 0 -1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_8
timestamp 1710899220
transform 1 0 824 0 1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_9
timestamp 1710899220
transform 1 0 936 0 1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_10
timestamp 1710899220
transform 1 0 952 0 -1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_11
timestamp 1710899220
transform 1 0 776 0 1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_12
timestamp 1710899220
transform 1 0 744 0 -1 1570
box -7 -3 39 105
use AOI21X1  AOI21X1_13
timestamp 1710899220
transform 1 0 256 0 1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_14
timestamp 1710899220
transform 1 0 288 0 1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_15
timestamp 1710899220
transform 1 0 240 0 1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_16
timestamp 1710899220
transform 1 0 224 0 -1 1570
box -7 -3 39 105
use AOI21X1  AOI21X1_17
timestamp 1710899220
transform 1 0 248 0 -1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_18
timestamp 1710899220
transform 1 0 216 0 -1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_19
timestamp 1710899220
transform 1 0 2416 0 -1 370
box -7 -3 39 105
use AOI21X1  AOI21X1_20
timestamp 1710899220
transform 1 0 2448 0 -1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_21
timestamp 1710899220
transform 1 0 2456 0 1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_22
timestamp 1710899220
transform 1 0 2520 0 -1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_23
timestamp 1710899220
transform 1 0 2368 0 -1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_24
timestamp 1710899220
transform 1 0 2320 0 1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_25
timestamp 1710899220
transform 1 0 2328 0 -1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_26
timestamp 1710899220
transform 1 0 2472 0 1 970
box -7 -3 39 105
use AOI22X1  AOI22X1_0
timestamp 1710899220
transform 1 0 1560 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_1
timestamp 1710899220
transform 1 0 1520 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_2
timestamp 1710899220
transform 1 0 2576 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_3
timestamp 1710899220
transform 1 0 2504 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_4
timestamp 1710899220
transform 1 0 2456 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_5
timestamp 1710899220
transform 1 0 2312 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_6
timestamp 1710899220
transform 1 0 2288 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_7
timestamp 1710899220
transform 1 0 2504 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_8
timestamp 1710899220
transform 1 0 2624 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_9
timestamp 1710899220
transform 1 0 2536 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_10
timestamp 1710899220
transform 1 0 2336 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_11
timestamp 1710899220
transform 1 0 2336 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_12
timestamp 1710899220
transform 1 0 2536 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_13
timestamp 1710899220
transform 1 0 2504 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_14
timestamp 1710899220
transform 1 0 2520 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_15
timestamp 1710899220
transform 1 0 2520 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_16
timestamp 1710899220
transform 1 0 2320 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_17
timestamp 1710899220
transform 1 0 2520 0 -1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_18
timestamp 1710899220
transform 1 0 2560 0 1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_19
timestamp 1710899220
transform 1 0 2360 0 1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_20
timestamp 1710899220
transform 1 0 2280 0 1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_21
timestamp 1710899220
transform 1 0 2248 0 -1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_22
timestamp 1710899220
transform 1 0 2000 0 -1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_23
timestamp 1710899220
transform 1 0 2144 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_24
timestamp 1710899220
transform 1 0 1944 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_25
timestamp 1710899220
transform 1 0 1928 0 1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_26
timestamp 1710899220
transform 1 0 1928 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_27
timestamp 1710899220
transform 1 0 1888 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_28
timestamp 1710899220
transform 1 0 1928 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_29
timestamp 1710899220
transform 1 0 2104 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_30
timestamp 1710899220
transform 1 0 2160 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_31
timestamp 1710899220
transform 1 0 2136 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_32
timestamp 1710899220
transform 1 0 2272 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_33
timestamp 1710899220
transform 1 0 2264 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_34
timestamp 1710899220
transform 1 0 432 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_35
timestamp 1710899220
transform 1 0 544 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_36
timestamp 1710899220
transform 1 0 1848 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_37
timestamp 1710899220
transform 1 0 1504 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_38
timestamp 1710899220
transform 1 0 864 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_39
timestamp 1710899220
transform 1 0 704 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_40
timestamp 1710899220
transform 1 0 1560 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_41
timestamp 1710899220
transform 1 0 1024 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_42
timestamp 1710899220
transform 1 0 1552 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_43
timestamp 1710899220
transform 1 0 1568 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_44
timestamp 1710899220
transform 1 0 928 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_45
timestamp 1710899220
transform 1 0 888 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_46
timestamp 1710899220
transform 1 0 456 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_47
timestamp 1710899220
transform 1 0 984 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_48
timestamp 1710899220
transform 1 0 968 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_49
timestamp 1710899220
transform 1 0 928 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_50
timestamp 1710899220
transform 1 0 520 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_51
timestamp 1710899220
transform 1 0 392 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_52
timestamp 1710899220
transform 1 0 1416 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_53
timestamp 1710899220
transform 1 0 1416 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_54
timestamp 1710899220
transform 1 0 904 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_55
timestamp 1710899220
transform 1 0 840 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_56
timestamp 1710899220
transform 1 0 968 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_57
timestamp 1710899220
transform 1 0 992 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_58
timestamp 1710899220
transform 1 0 896 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_59
timestamp 1710899220
transform 1 0 784 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_60
timestamp 1710899220
transform 1 0 1016 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_61
timestamp 1710899220
transform 1 0 888 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_62
timestamp 1710899220
transform 1 0 840 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_63
timestamp 1710899220
transform 1 0 1032 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_64
timestamp 1710899220
transform 1 0 880 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_65
timestamp 1710899220
transform 1 0 928 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_66
timestamp 1710899220
transform 1 0 784 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_67
timestamp 1710899220
transform 1 0 688 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_68
timestamp 1710899220
transform 1 0 696 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_69
timestamp 1710899220
transform 1 0 848 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_70
timestamp 1710899220
transform 1 0 680 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_71
timestamp 1710899220
transform 1 0 688 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_72
timestamp 1710899220
transform 1 0 776 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_73
timestamp 1710899220
transform 1 0 224 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_74
timestamp 1710899220
transform 1 0 144 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_75
timestamp 1710899220
transform 1 0 176 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_76
timestamp 1710899220
transform 1 0 2400 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_77
timestamp 1710899220
transform 1 0 2584 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_78
timestamp 1710899220
transform 1 0 2544 0 -1 970
box -8 -3 46 105
use BUFX2  BUFX2_0
timestamp 1710899220
transform 1 0 2008 0 -1 1370
box -5 -3 28 105
use BUFX2  BUFX2_1
timestamp 1710899220
transform 1 0 1800 0 -1 1370
box -5 -3 28 105
use BUFX2  BUFX2_2
timestamp 1710899220
transform 1 0 1824 0 -1 1370
box -5 -3 28 105
use BUFX2  BUFX2_3
timestamp 1710899220
transform 1 0 2304 0 1 970
box -5 -3 28 105
use BUFX2  BUFX2_4
timestamp 1710899220
transform 1 0 1912 0 -1 1370
box -5 -3 28 105
use BUFX2  BUFX2_5
timestamp 1710899220
transform 1 0 1936 0 -1 1370
box -5 -3 28 105
use BUFX2  BUFX2_6
timestamp 1710899220
transform 1 0 1928 0 1 1770
box -5 -3 28 105
use BUFX2  BUFX2_7
timestamp 1710899220
transform 1 0 1888 0 1 970
box -5 -3 28 105
use BUFX2  BUFX2_8
timestamp 1710899220
transform 1 0 1904 0 1 1770
box -5 -3 28 105
use BUFX2  BUFX2_9
timestamp 1710899220
transform 1 0 2264 0 -1 1570
box -5 -3 28 105
use BUFX2  BUFX2_10
timestamp 1710899220
transform 1 0 2104 0 1 1370
box -5 -3 28 105
use BUFX2  BUFX2_11
timestamp 1710899220
transform 1 0 2040 0 -1 1170
box -5 -3 28 105
use BUFX2  BUFX2_12
timestamp 1710899220
transform 1 0 1216 0 -1 770
box -5 -3 28 105
use BUFX2  BUFX2_13
timestamp 1710899220
transform 1 0 1296 0 -1 770
box -5 -3 28 105
use BUFX2  BUFX2_14
timestamp 1710899220
transform 1 0 1240 0 -1 770
box -5 -3 28 105
use BUFX2  BUFX2_15
timestamp 1710899220
transform 1 0 1776 0 1 1370
box -5 -3 28 105
use BUFX2  BUFX2_16
timestamp 1710899220
transform 1 0 1744 0 1 1370
box -5 -3 28 105
use BUFX2  BUFX2_17
timestamp 1710899220
transform 1 0 1800 0 1 1370
box -5 -3 28 105
use BUFX2  BUFX2_18
timestamp 1710899220
transform 1 0 1688 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_19
timestamp 1710899220
transform 1 0 1440 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_20
timestamp 1710899220
transform 1 0 1296 0 -1 570
box -5 -3 28 105
use BUFX2  BUFX2_21
timestamp 1710899220
transform 1 0 1248 0 -1 570
box -5 -3 28 105
use BUFX2  BUFX2_22
timestamp 1710899220
transform 1 0 1528 0 -1 570
box -5 -3 28 105
use BUFX2  BUFX2_23
timestamp 1710899220
transform 1 0 1272 0 -1 570
box -5 -3 28 105
use BUFX2  BUFX2_24
timestamp 1710899220
transform 1 0 1840 0 -1 770
box -5 -3 28 105
use BUFX2  BUFX2_25
timestamp 1710899220
transform 1 0 720 0 1 570
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_0
timestamp 1710899220
transform 1 0 2144 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_1
timestamp 1710899220
transform 1 0 1400 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_2
timestamp 1710899220
transform 1 0 1592 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_3
timestamp 1710899220
transform 1 0 1672 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_4
timestamp 1710899220
transform 1 0 1224 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_5
timestamp 1710899220
transform 1 0 1840 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_6
timestamp 1710899220
transform 1 0 1432 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_7
timestamp 1710899220
transform 1 0 1752 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_8
timestamp 1710899220
transform 1 0 1632 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_9
timestamp 1710899220
transform 1 0 1792 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_10
timestamp 1710899220
transform 1 0 1760 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_11
timestamp 1710899220
transform 1 0 1024 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_12
timestamp 1710899220
transform 1 0 1136 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_13
timestamp 1710899220
transform 1 0 984 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_14
timestamp 1710899220
transform 1 0 1008 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_15
timestamp 1710899220
transform 1 0 1432 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_16
timestamp 1710899220
transform 1 0 744 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_17
timestamp 1710899220
transform 1 0 1192 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_18
timestamp 1710899220
transform 1 0 528 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_19
timestamp 1710899220
transform 1 0 464 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_20
timestamp 1710899220
transform 1 0 808 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_21
timestamp 1710899220
transform 1 0 936 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_22
timestamp 1710899220
transform 1 0 688 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_23
timestamp 1710899220
transform 1 0 768 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_24
timestamp 1710899220
transform 1 0 832 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_25
timestamp 1710899220
transform 1 0 872 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_26
timestamp 1710899220
transform 1 0 912 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_27
timestamp 1710899220
transform 1 0 1216 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_28
timestamp 1710899220
transform 1 0 1384 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_29
timestamp 1710899220
transform 1 0 1576 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_30
timestamp 1710899220
transform 1 0 1872 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_31
timestamp 1710899220
transform 1 0 1888 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_32
timestamp 1710899220
transform 1 0 2032 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_33
timestamp 1710899220
transform 1 0 2128 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_34
timestamp 1710899220
transform 1 0 2168 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_35
timestamp 1710899220
transform 1 0 1936 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_36
timestamp 1710899220
transform 1 0 2328 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_37
timestamp 1710899220
transform 1 0 1200 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_38
timestamp 1710899220
transform 1 0 1352 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_39
timestamp 1710899220
transform 1 0 1216 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_40
timestamp 1710899220
transform 1 0 1096 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_41
timestamp 1710899220
transform 1 0 1104 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_42
timestamp 1710899220
transform 1 0 568 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_43
timestamp 1710899220
transform 1 0 544 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_44
timestamp 1710899220
transform 1 0 400 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_45
timestamp 1710899220
transform 1 0 440 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_46
timestamp 1710899220
transform 1 0 1152 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_47
timestamp 1710899220
transform 1 0 848 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_48
timestamp 1710899220
transform 1 0 736 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_49
timestamp 1710899220
transform 1 0 552 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_50
timestamp 1710899220
transform 1 0 656 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_51
timestamp 1710899220
transform 1 0 752 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_52
timestamp 1710899220
transform 1 0 856 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_53
timestamp 1710899220
transform 1 0 1064 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_54
timestamp 1710899220
transform 1 0 1256 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_55
timestamp 1710899220
transform 1 0 1456 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_56
timestamp 1710899220
transform 1 0 1512 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_57
timestamp 1710899220
transform 1 0 1352 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_58
timestamp 1710899220
transform 1 0 1760 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_59
timestamp 1710899220
transform 1 0 1848 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_60
timestamp 1710899220
transform 1 0 1840 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_61
timestamp 1710899220
transform 1 0 1424 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_62
timestamp 1710899220
transform 1 0 1424 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_63
timestamp 1710899220
transform 1 0 1552 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_64
timestamp 1710899220
transform 1 0 1832 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_65
timestamp 1710899220
transform 1 0 1960 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_66
timestamp 1710899220
transform 1 0 1456 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_67
timestamp 1710899220
transform 1 0 584 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_68
timestamp 1710899220
transform 1 0 232 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_69
timestamp 1710899220
transform 1 0 168 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_70
timestamp 1710899220
transform 1 0 176 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_71
timestamp 1710899220
transform 1 0 1160 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_72
timestamp 1710899220
transform 1 0 912 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_73
timestamp 1710899220
transform 1 0 816 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_74
timestamp 1710899220
transform 1 0 440 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_75
timestamp 1710899220
transform 1 0 168 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_76
timestamp 1710899220
transform 1 0 232 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_77
timestamp 1710899220
transform 1 0 952 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_78
timestamp 1710899220
transform 1 0 1048 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_79
timestamp 1710899220
transform 1 0 1144 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_80
timestamp 1710899220
transform 1 0 1712 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_81
timestamp 1710899220
transform 1 0 1552 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_82
timestamp 1710899220
transform 1 0 1664 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_83
timestamp 1710899220
transform 1 0 2040 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_84
timestamp 1710899220
transform 1 0 2032 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_85
timestamp 1710899220
transform 1 0 1944 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_86
timestamp 1710899220
transform 1 0 1560 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_87
timestamp 1710899220
transform 1 0 1664 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_88
timestamp 1710899220
transform 1 0 1904 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_89
timestamp 1710899220
transform 1 0 2008 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_90
timestamp 1710899220
transform 1 0 2032 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_91
timestamp 1710899220
transform 1 0 2056 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_92
timestamp 1710899220
transform 1 0 2056 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_93
timestamp 1710899220
transform 1 0 1952 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_94
timestamp 1710899220
transform 1 0 2152 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_95
timestamp 1710899220
transform 1 0 2336 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_96
timestamp 1710899220
transform 1 0 2024 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_97
timestamp 1710899220
transform 1 0 2240 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_98
timestamp 1710899220
transform 1 0 1984 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_99
timestamp 1710899220
transform 1 0 1816 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_100
timestamp 1710899220
transform 1 0 1760 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_101
timestamp 1710899220
transform 1 0 1816 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_102
timestamp 1710899220
transform 1 0 1816 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_103
timestamp 1710899220
transform 1 0 1832 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_104
timestamp 1710899220
transform 1 0 2200 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_105
timestamp 1710899220
transform 1 0 2056 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_106
timestamp 1710899220
transform 1 0 2320 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_107
timestamp 1710899220
transform 1 0 2296 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_108
timestamp 1710899220
transform 1 0 2424 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_109
timestamp 1710899220
transform 1 0 2552 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_110
timestamp 1710899220
transform 1 0 2576 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_111
timestamp 1710899220
transform 1 0 2408 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_112
timestamp 1710899220
transform 1 0 2560 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_113
timestamp 1710899220
transform 1 0 2576 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_114
timestamp 1710899220
transform 1 0 2560 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_115
timestamp 1710899220
transform 1 0 2576 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_116
timestamp 1710899220
transform 1 0 2224 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_117
timestamp 1710899220
transform 1 0 2224 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_118
timestamp 1710899220
transform 1 0 2576 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_119
timestamp 1710899220
transform 1 0 2528 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_120
timestamp 1710899220
transform 1 0 2408 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_121
timestamp 1710899220
transform 1 0 2272 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_122
timestamp 1710899220
transform 1 0 2280 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_123
timestamp 1710899220
transform 1 0 2464 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_124
timestamp 1710899220
transform 1 0 2576 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_125
timestamp 1710899220
transform 1 0 2560 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_126
timestamp 1710899220
transform 1 0 1832 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_127
timestamp 1710899220
transform 1 0 1880 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_128
timestamp 1710899220
transform 1 0 2240 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_129
timestamp 1710899220
transform 1 0 2152 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_130
timestamp 1710899220
transform 1 0 2480 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_131
timestamp 1710899220
transform 1 0 2432 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_132
timestamp 1710899220
transform 1 0 2528 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_133
timestamp 1710899220
transform 1 0 2384 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_134
timestamp 1710899220
transform 1 0 2576 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_135
timestamp 1710899220
transform 1 0 2328 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_136
timestamp 1710899220
transform 1 0 2576 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_137
timestamp 1710899220
transform 1 0 2288 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_138
timestamp 1710899220
transform 1 0 2088 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_139
timestamp 1710899220
transform 1 0 2192 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_140
timestamp 1710899220
transform 1 0 2128 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_141
timestamp 1710899220
transform 1 0 2072 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_142
timestamp 1710899220
transform 1 0 2576 0 1 170
box -8 -3 104 105
use FAX1  FAX1_0
timestamp 1710899220
transform 1 0 784 0 -1 2370
box -5 -3 126 105
use FAX1  FAX1_1
timestamp 1710899220
transform 1 0 992 0 -1 2370
box -5 -3 126 105
use FAX1  FAX1_2
timestamp 1710899220
transform 1 0 1144 0 -1 2370
box -5 -3 126 105
use FAX1  FAX1_3
timestamp 1710899220
transform 1 0 1232 0 1 2170
box -5 -3 126 105
use FAX1  FAX1_4
timestamp 1710899220
transform 1 0 104 0 -1 2170
box -5 -3 126 105
use FAX1  FAX1_5
timestamp 1710899220
transform 1 0 232 0 -1 2170
box -5 -3 126 105
use FAX1  FAX1_6
timestamp 1710899220
transform 1 0 376 0 -1 2170
box -5 -3 126 105
use FAX1  FAX1_7
timestamp 1710899220
transform 1 0 528 0 1 2170
box -5 -3 126 105
use FAX1  FAX1_8
timestamp 1710899220
transform 1 0 848 0 1 2170
box -5 -3 126 105
use FAX1  FAX1_9
timestamp 1710899220
transform 1 0 968 0 1 2170
box -5 -3 126 105
use FAX1  FAX1_10
timestamp 1710899220
transform 1 0 1088 0 1 2170
box -5 -3 126 105
use FAX1  FAX1_11
timestamp 1710899220
transform 1 0 128 0 -1 1970
box -5 -3 126 105
use FAX1  FAX1_12
timestamp 1710899220
transform 1 0 304 0 1 1970
box -5 -3 126 105
use FAX1  FAX1_13
timestamp 1710899220
transform 1 0 304 0 -1 1970
box -5 -3 126 105
use FAX1  FAX1_14
timestamp 1710899220
transform 1 0 520 0 -1 2170
box -5 -3 126 105
use FAX1  FAX1_15
timestamp 1710899220
transform 1 0 528 0 1 1970
box -5 -3 126 105
use FAX1  FAX1_16
timestamp 1710899220
transform 1 0 728 0 1 2170
box -5 -3 126 105
use FAX1  FAX1_17
timestamp 1710899220
transform 1 0 776 0 -1 2170
box -5 -3 126 105
use FAX1  FAX1_18
timestamp 1710899220
transform 1 0 928 0 -1 2170
box -5 -3 126 105
use FILL  FILL_0
timestamp 1710899220
transform 1 0 2664 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1
timestamp 1710899220
transform 1 0 2656 0 -1 2570
box -8 -3 16 105
use FILL  FILL_2
timestamp 1710899220
transform 1 0 2648 0 -1 2570
box -8 -3 16 105
use FILL  FILL_3
timestamp 1710899220
transform 1 0 2544 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4
timestamp 1710899220
transform 1 0 2536 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5
timestamp 1710899220
transform 1 0 2528 0 -1 2570
box -8 -3 16 105
use FILL  FILL_6
timestamp 1710899220
transform 1 0 2520 0 -1 2570
box -8 -3 16 105
use FILL  FILL_7
timestamp 1710899220
transform 1 0 2416 0 -1 2570
box -8 -3 16 105
use FILL  FILL_8
timestamp 1710899220
transform 1 0 2408 0 -1 2570
box -8 -3 16 105
use FILL  FILL_9
timestamp 1710899220
transform 1 0 2664 0 1 2370
box -8 -3 16 105
use FILL  FILL_10
timestamp 1710899220
transform 1 0 2656 0 1 2370
box -8 -3 16 105
use FILL  FILL_11
timestamp 1710899220
transform 1 0 2648 0 1 2370
box -8 -3 16 105
use FILL  FILL_12
timestamp 1710899220
transform 1 0 2640 0 1 2370
box -8 -3 16 105
use FILL  FILL_13
timestamp 1710899220
transform 1 0 2632 0 1 2370
box -8 -3 16 105
use FILL  FILL_14
timestamp 1710899220
transform 1 0 2624 0 1 2370
box -8 -3 16 105
use FILL  FILL_15
timestamp 1710899220
transform 1 0 2616 0 1 2370
box -8 -3 16 105
use FILL  FILL_16
timestamp 1710899220
transform 1 0 2352 0 1 2370
box -8 -3 16 105
use FILL  FILL_17
timestamp 1710899220
transform 1 0 2344 0 1 2370
box -8 -3 16 105
use FILL  FILL_18
timestamp 1710899220
transform 1 0 2336 0 1 2370
box -8 -3 16 105
use FILL  FILL_19
timestamp 1710899220
transform 1 0 2192 0 1 2370
box -8 -3 16 105
use FILL  FILL_20
timestamp 1710899220
transform 1 0 2184 0 1 2370
box -8 -3 16 105
use FILL  FILL_21
timestamp 1710899220
transform 1 0 2176 0 1 2370
box -8 -3 16 105
use FILL  FILL_22
timestamp 1710899220
transform 1 0 2168 0 1 2370
box -8 -3 16 105
use FILL  FILL_23
timestamp 1710899220
transform 1 0 2160 0 1 2370
box -8 -3 16 105
use FILL  FILL_24
timestamp 1710899220
transform 1 0 2152 0 1 2370
box -8 -3 16 105
use FILL  FILL_25
timestamp 1710899220
transform 1 0 2144 0 1 2370
box -8 -3 16 105
use FILL  FILL_26
timestamp 1710899220
transform 1 0 2136 0 1 2370
box -8 -3 16 105
use FILL  FILL_27
timestamp 1710899220
transform 1 0 2128 0 1 2370
box -8 -3 16 105
use FILL  FILL_28
timestamp 1710899220
transform 1 0 2120 0 1 2370
box -8 -3 16 105
use FILL  FILL_29
timestamp 1710899220
transform 1 0 2112 0 1 2370
box -8 -3 16 105
use FILL  FILL_30
timestamp 1710899220
transform 1 0 2104 0 1 2370
box -8 -3 16 105
use FILL  FILL_31
timestamp 1710899220
transform 1 0 2096 0 1 2370
box -8 -3 16 105
use FILL  FILL_32
timestamp 1710899220
transform 1 0 2088 0 1 2370
box -8 -3 16 105
use FILL  FILL_33
timestamp 1710899220
transform 1 0 2080 0 1 2370
box -8 -3 16 105
use FILL  FILL_34
timestamp 1710899220
transform 1 0 2072 0 1 2370
box -8 -3 16 105
use FILL  FILL_35
timestamp 1710899220
transform 1 0 2064 0 1 2370
box -8 -3 16 105
use FILL  FILL_36
timestamp 1710899220
transform 1 0 2056 0 1 2370
box -8 -3 16 105
use FILL  FILL_37
timestamp 1710899220
transform 1 0 2048 0 1 2370
box -8 -3 16 105
use FILL  FILL_38
timestamp 1710899220
transform 1 0 1808 0 1 2370
box -8 -3 16 105
use FILL  FILL_39
timestamp 1710899220
transform 1 0 1800 0 1 2370
box -8 -3 16 105
use FILL  FILL_40
timestamp 1710899220
transform 1 0 1792 0 1 2370
box -8 -3 16 105
use FILL  FILL_41
timestamp 1710899220
transform 1 0 1784 0 1 2370
box -8 -3 16 105
use FILL  FILL_42
timestamp 1710899220
transform 1 0 1776 0 1 2370
box -8 -3 16 105
use FILL  FILL_43
timestamp 1710899220
transform 1 0 1768 0 1 2370
box -8 -3 16 105
use FILL  FILL_44
timestamp 1710899220
transform 1 0 1760 0 1 2370
box -8 -3 16 105
use FILL  FILL_45
timestamp 1710899220
transform 1 0 1752 0 1 2370
box -8 -3 16 105
use FILL  FILL_46
timestamp 1710899220
transform 1 0 1744 0 1 2370
box -8 -3 16 105
use FILL  FILL_47
timestamp 1710899220
transform 1 0 1672 0 1 2370
box -8 -3 16 105
use FILL  FILL_48
timestamp 1710899220
transform 1 0 1584 0 1 2370
box -8 -3 16 105
use FILL  FILL_49
timestamp 1710899220
transform 1 0 1576 0 1 2370
box -8 -3 16 105
use FILL  FILL_50
timestamp 1710899220
transform 1 0 1568 0 1 2370
box -8 -3 16 105
use FILL  FILL_51
timestamp 1710899220
transform 1 0 1544 0 1 2370
box -8 -3 16 105
use FILL  FILL_52
timestamp 1710899220
transform 1 0 1536 0 1 2370
box -8 -3 16 105
use FILL  FILL_53
timestamp 1710899220
transform 1 0 1464 0 1 2370
box -8 -3 16 105
use FILL  FILL_54
timestamp 1710899220
transform 1 0 1456 0 1 2370
box -8 -3 16 105
use FILL  FILL_55
timestamp 1710899220
transform 1 0 1448 0 1 2370
box -8 -3 16 105
use FILL  FILL_56
timestamp 1710899220
transform 1 0 1360 0 1 2370
box -8 -3 16 105
use FILL  FILL_57
timestamp 1710899220
transform 1 0 1352 0 1 2370
box -8 -3 16 105
use FILL  FILL_58
timestamp 1710899220
transform 1 0 1320 0 1 2370
box -8 -3 16 105
use FILL  FILL_59
timestamp 1710899220
transform 1 0 1312 0 1 2370
box -8 -3 16 105
use FILL  FILL_60
timestamp 1710899220
transform 1 0 1288 0 1 2370
box -8 -3 16 105
use FILL  FILL_61
timestamp 1710899220
transform 1 0 1280 0 1 2370
box -8 -3 16 105
use FILL  FILL_62
timestamp 1710899220
transform 1 0 1272 0 1 2370
box -8 -3 16 105
use FILL  FILL_63
timestamp 1710899220
transform 1 0 1200 0 1 2370
box -8 -3 16 105
use FILL  FILL_64
timestamp 1710899220
transform 1 0 1144 0 1 2370
box -8 -3 16 105
use FILL  FILL_65
timestamp 1710899220
transform 1 0 1080 0 1 2370
box -8 -3 16 105
use FILL  FILL_66
timestamp 1710899220
transform 1 0 1032 0 1 2370
box -8 -3 16 105
use FILL  FILL_67
timestamp 1710899220
transform 1 0 1024 0 1 2370
box -8 -3 16 105
use FILL  FILL_68
timestamp 1710899220
transform 1 0 1016 0 1 2370
box -8 -3 16 105
use FILL  FILL_69
timestamp 1710899220
transform 1 0 1008 0 1 2370
box -8 -3 16 105
use FILL  FILL_70
timestamp 1710899220
transform 1 0 888 0 1 2370
box -8 -3 16 105
use FILL  FILL_71
timestamp 1710899220
transform 1 0 880 0 1 2370
box -8 -3 16 105
use FILL  FILL_72
timestamp 1710899220
transform 1 0 848 0 1 2370
box -8 -3 16 105
use FILL  FILL_73
timestamp 1710899220
transform 1 0 776 0 1 2370
box -8 -3 16 105
use FILL  FILL_74
timestamp 1710899220
transform 1 0 672 0 1 2370
box -8 -3 16 105
use FILL  FILL_75
timestamp 1710899220
transform 1 0 664 0 1 2370
box -8 -3 16 105
use FILL  FILL_76
timestamp 1710899220
transform 1 0 656 0 1 2370
box -8 -3 16 105
use FILL  FILL_77
timestamp 1710899220
transform 1 0 584 0 1 2370
box -8 -3 16 105
use FILL  FILL_78
timestamp 1710899220
transform 1 0 576 0 1 2370
box -8 -3 16 105
use FILL  FILL_79
timestamp 1710899220
transform 1 0 488 0 1 2370
box -8 -3 16 105
use FILL  FILL_80
timestamp 1710899220
transform 1 0 424 0 1 2370
box -8 -3 16 105
use FILL  FILL_81
timestamp 1710899220
transform 1 0 392 0 1 2370
box -8 -3 16 105
use FILL  FILL_82
timestamp 1710899220
transform 1 0 384 0 1 2370
box -8 -3 16 105
use FILL  FILL_83
timestamp 1710899220
transform 1 0 376 0 1 2370
box -8 -3 16 105
use FILL  FILL_84
timestamp 1710899220
transform 1 0 368 0 1 2370
box -8 -3 16 105
use FILL  FILL_85
timestamp 1710899220
transform 1 0 312 0 1 2370
box -8 -3 16 105
use FILL  FILL_86
timestamp 1710899220
transform 1 0 304 0 1 2370
box -8 -3 16 105
use FILL  FILL_87
timestamp 1710899220
transform 1 0 296 0 1 2370
box -8 -3 16 105
use FILL  FILL_88
timestamp 1710899220
transform 1 0 288 0 1 2370
box -8 -3 16 105
use FILL  FILL_89
timestamp 1710899220
transform 1 0 264 0 1 2370
box -8 -3 16 105
use FILL  FILL_90
timestamp 1710899220
transform 1 0 240 0 1 2370
box -8 -3 16 105
use FILL  FILL_91
timestamp 1710899220
transform 1 0 232 0 1 2370
box -8 -3 16 105
use FILL  FILL_92
timestamp 1710899220
transform 1 0 176 0 1 2370
box -8 -3 16 105
use FILL  FILL_93
timestamp 1710899220
transform 1 0 168 0 1 2370
box -8 -3 16 105
use FILL  FILL_94
timestamp 1710899220
transform 1 0 160 0 1 2370
box -8 -3 16 105
use FILL  FILL_95
timestamp 1710899220
transform 1 0 152 0 1 2370
box -8 -3 16 105
use FILL  FILL_96
timestamp 1710899220
transform 1 0 2432 0 -1 2370
box -8 -3 16 105
use FILL  FILL_97
timestamp 1710899220
transform 1 0 2424 0 -1 2370
box -8 -3 16 105
use FILL  FILL_98
timestamp 1710899220
transform 1 0 2416 0 -1 2370
box -8 -3 16 105
use FILL  FILL_99
timestamp 1710899220
transform 1 0 2312 0 -1 2370
box -8 -3 16 105
use FILL  FILL_100
timestamp 1710899220
transform 1 0 2304 0 -1 2370
box -8 -3 16 105
use FILL  FILL_101
timestamp 1710899220
transform 1 0 2240 0 -1 2370
box -8 -3 16 105
use FILL  FILL_102
timestamp 1710899220
transform 1 0 2232 0 -1 2370
box -8 -3 16 105
use FILL  FILL_103
timestamp 1710899220
transform 1 0 2144 0 -1 2370
box -8 -3 16 105
use FILL  FILL_104
timestamp 1710899220
transform 1 0 2056 0 -1 2370
box -8 -3 16 105
use FILL  FILL_105
timestamp 1710899220
transform 1 0 1992 0 -1 2370
box -8 -3 16 105
use FILL  FILL_106
timestamp 1710899220
transform 1 0 1984 0 -1 2370
box -8 -3 16 105
use FILL  FILL_107
timestamp 1710899220
transform 1 0 1976 0 -1 2370
box -8 -3 16 105
use FILL  FILL_108
timestamp 1710899220
transform 1 0 1968 0 -1 2370
box -8 -3 16 105
use FILL  FILL_109
timestamp 1710899220
transform 1 0 1960 0 -1 2370
box -8 -3 16 105
use FILL  FILL_110
timestamp 1710899220
transform 1 0 1952 0 -1 2370
box -8 -3 16 105
use FILL  FILL_111
timestamp 1710899220
transform 1 0 1944 0 -1 2370
box -8 -3 16 105
use FILL  FILL_112
timestamp 1710899220
transform 1 0 1936 0 -1 2370
box -8 -3 16 105
use FILL  FILL_113
timestamp 1710899220
transform 1 0 1928 0 -1 2370
box -8 -3 16 105
use FILL  FILL_114
timestamp 1710899220
transform 1 0 1920 0 -1 2370
box -8 -3 16 105
use FILL  FILL_115
timestamp 1710899220
transform 1 0 1912 0 -1 2370
box -8 -3 16 105
use FILL  FILL_116
timestamp 1710899220
transform 1 0 1904 0 -1 2370
box -8 -3 16 105
use FILL  FILL_117
timestamp 1710899220
transform 1 0 1896 0 -1 2370
box -8 -3 16 105
use FILL  FILL_118
timestamp 1710899220
transform 1 0 1888 0 -1 2370
box -8 -3 16 105
use FILL  FILL_119
timestamp 1710899220
transform 1 0 1880 0 -1 2370
box -8 -3 16 105
use FILL  FILL_120
timestamp 1710899220
transform 1 0 1872 0 -1 2370
box -8 -3 16 105
use FILL  FILL_121
timestamp 1710899220
transform 1 0 1864 0 -1 2370
box -8 -3 16 105
use FILL  FILL_122
timestamp 1710899220
transform 1 0 1856 0 -1 2370
box -8 -3 16 105
use FILL  FILL_123
timestamp 1710899220
transform 1 0 1848 0 -1 2370
box -8 -3 16 105
use FILL  FILL_124
timestamp 1710899220
transform 1 0 1840 0 -1 2370
box -8 -3 16 105
use FILL  FILL_125
timestamp 1710899220
transform 1 0 1832 0 -1 2370
box -8 -3 16 105
use FILL  FILL_126
timestamp 1710899220
transform 1 0 1744 0 -1 2370
box -8 -3 16 105
use FILL  FILL_127
timestamp 1710899220
transform 1 0 1736 0 -1 2370
box -8 -3 16 105
use FILL  FILL_128
timestamp 1710899220
transform 1 0 1648 0 -1 2370
box -8 -3 16 105
use FILL  FILL_129
timestamp 1710899220
transform 1 0 1640 0 -1 2370
box -8 -3 16 105
use FILL  FILL_130
timestamp 1710899220
transform 1 0 1568 0 -1 2370
box -8 -3 16 105
use FILL  FILL_131
timestamp 1710899220
transform 1 0 1480 0 -1 2370
box -8 -3 16 105
use FILL  FILL_132
timestamp 1710899220
transform 1 0 1472 0 -1 2370
box -8 -3 16 105
use FILL  FILL_133
timestamp 1710899220
transform 1 0 1464 0 -1 2370
box -8 -3 16 105
use FILL  FILL_134
timestamp 1710899220
transform 1 0 1456 0 -1 2370
box -8 -3 16 105
use FILL  FILL_135
timestamp 1710899220
transform 1 0 1384 0 -1 2370
box -8 -3 16 105
use FILL  FILL_136
timestamp 1710899220
transform 1 0 1272 0 -1 2370
box -8 -3 16 105
use FILL  FILL_137
timestamp 1710899220
transform 1 0 1264 0 -1 2370
box -8 -3 16 105
use FILL  FILL_138
timestamp 1710899220
transform 1 0 1136 0 -1 2370
box -8 -3 16 105
use FILL  FILL_139
timestamp 1710899220
transform 1 0 1128 0 -1 2370
box -8 -3 16 105
use FILL  FILL_140
timestamp 1710899220
transform 1 0 1120 0 -1 2370
box -8 -3 16 105
use FILL  FILL_141
timestamp 1710899220
transform 1 0 1112 0 -1 2370
box -8 -3 16 105
use FILL  FILL_142
timestamp 1710899220
transform 1 0 984 0 -1 2370
box -8 -3 16 105
use FILL  FILL_143
timestamp 1710899220
transform 1 0 976 0 -1 2370
box -8 -3 16 105
use FILL  FILL_144
timestamp 1710899220
transform 1 0 968 0 -1 2370
box -8 -3 16 105
use FILL  FILL_145
timestamp 1710899220
transform 1 0 904 0 -1 2370
box -8 -3 16 105
use FILL  FILL_146
timestamp 1710899220
transform 1 0 776 0 -1 2370
box -8 -3 16 105
use FILL  FILL_147
timestamp 1710899220
transform 1 0 768 0 -1 2370
box -8 -3 16 105
use FILL  FILL_148
timestamp 1710899220
transform 1 0 760 0 -1 2370
box -8 -3 16 105
use FILL  FILL_149
timestamp 1710899220
transform 1 0 736 0 -1 2370
box -8 -3 16 105
use FILL  FILL_150
timestamp 1710899220
transform 1 0 728 0 -1 2370
box -8 -3 16 105
use FILL  FILL_151
timestamp 1710899220
transform 1 0 720 0 -1 2370
box -8 -3 16 105
use FILL  FILL_152
timestamp 1710899220
transform 1 0 712 0 -1 2370
box -8 -3 16 105
use FILL  FILL_153
timestamp 1710899220
transform 1 0 640 0 -1 2370
box -8 -3 16 105
use FILL  FILL_154
timestamp 1710899220
transform 1 0 576 0 -1 2370
box -8 -3 16 105
use FILL  FILL_155
timestamp 1710899220
transform 1 0 568 0 -1 2370
box -8 -3 16 105
use FILL  FILL_156
timestamp 1710899220
transform 1 0 560 0 -1 2370
box -8 -3 16 105
use FILL  FILL_157
timestamp 1710899220
transform 1 0 472 0 -1 2370
box -8 -3 16 105
use FILL  FILL_158
timestamp 1710899220
transform 1 0 448 0 -1 2370
box -8 -3 16 105
use FILL  FILL_159
timestamp 1710899220
transform 1 0 440 0 -1 2370
box -8 -3 16 105
use FILL  FILL_160
timestamp 1710899220
transform 1 0 368 0 -1 2370
box -8 -3 16 105
use FILL  FILL_161
timestamp 1710899220
transform 1 0 280 0 -1 2370
box -8 -3 16 105
use FILL  FILL_162
timestamp 1710899220
transform 1 0 208 0 -1 2370
box -8 -3 16 105
use FILL  FILL_163
timestamp 1710899220
transform 1 0 200 0 -1 2370
box -8 -3 16 105
use FILL  FILL_164
timestamp 1710899220
transform 1 0 112 0 -1 2370
box -8 -3 16 105
use FILL  FILL_165
timestamp 1710899220
transform 1 0 104 0 -1 2370
box -8 -3 16 105
use FILL  FILL_166
timestamp 1710899220
transform 1 0 96 0 -1 2370
box -8 -3 16 105
use FILL  FILL_167
timestamp 1710899220
transform 1 0 88 0 -1 2370
box -8 -3 16 105
use FILL  FILL_168
timestamp 1710899220
transform 1 0 80 0 -1 2370
box -8 -3 16 105
use FILL  FILL_169
timestamp 1710899220
transform 1 0 72 0 -1 2370
box -8 -3 16 105
use FILL  FILL_170
timestamp 1710899220
transform 1 0 2048 0 1 2170
box -8 -3 16 105
use FILL  FILL_171
timestamp 1710899220
transform 1 0 1808 0 1 2170
box -8 -3 16 105
use FILL  FILL_172
timestamp 1710899220
transform 1 0 1800 0 1 2170
box -8 -3 16 105
use FILL  FILL_173
timestamp 1710899220
transform 1 0 1712 0 1 2170
box -8 -3 16 105
use FILL  FILL_174
timestamp 1710899220
transform 1 0 1704 0 1 2170
box -8 -3 16 105
use FILL  FILL_175
timestamp 1710899220
transform 1 0 1696 0 1 2170
box -8 -3 16 105
use FILL  FILL_176
timestamp 1710899220
transform 1 0 1624 0 1 2170
box -8 -3 16 105
use FILL  FILL_177
timestamp 1710899220
transform 1 0 1616 0 1 2170
box -8 -3 16 105
use FILL  FILL_178
timestamp 1710899220
transform 1 0 1560 0 1 2170
box -8 -3 16 105
use FILL  FILL_179
timestamp 1710899220
transform 1 0 1552 0 1 2170
box -8 -3 16 105
use FILL  FILL_180
timestamp 1710899220
transform 1 0 1544 0 1 2170
box -8 -3 16 105
use FILL  FILL_181
timestamp 1710899220
transform 1 0 1360 0 1 2170
box -8 -3 16 105
use FILL  FILL_182
timestamp 1710899220
transform 1 0 1352 0 1 2170
box -8 -3 16 105
use FILL  FILL_183
timestamp 1710899220
transform 1 0 1224 0 1 2170
box -8 -3 16 105
use FILL  FILL_184
timestamp 1710899220
transform 1 0 1216 0 1 2170
box -8 -3 16 105
use FILL  FILL_185
timestamp 1710899220
transform 1 0 1208 0 1 2170
box -8 -3 16 105
use FILL  FILL_186
timestamp 1710899220
transform 1 0 520 0 1 2170
box -8 -3 16 105
use FILL  FILL_187
timestamp 1710899220
transform 1 0 480 0 1 2170
box -8 -3 16 105
use FILL  FILL_188
timestamp 1710899220
transform 1 0 416 0 1 2170
box -8 -3 16 105
use FILL  FILL_189
timestamp 1710899220
transform 1 0 376 0 1 2170
box -8 -3 16 105
use FILL  FILL_190
timestamp 1710899220
transform 1 0 368 0 1 2170
box -8 -3 16 105
use FILL  FILL_191
timestamp 1710899220
transform 1 0 304 0 1 2170
box -8 -3 16 105
use FILL  FILL_192
timestamp 1710899220
transform 1 0 264 0 1 2170
box -8 -3 16 105
use FILL  FILL_193
timestamp 1710899220
transform 1 0 256 0 1 2170
box -8 -3 16 105
use FILL  FILL_194
timestamp 1710899220
transform 1 0 160 0 1 2170
box -8 -3 16 105
use FILL  FILL_195
timestamp 1710899220
transform 1 0 152 0 1 2170
box -8 -3 16 105
use FILL  FILL_196
timestamp 1710899220
transform 1 0 2664 0 -1 2170
box -8 -3 16 105
use FILL  FILL_197
timestamp 1710899220
transform 1 0 2656 0 -1 2170
box -8 -3 16 105
use FILL  FILL_198
timestamp 1710899220
transform 1 0 2648 0 -1 2170
box -8 -3 16 105
use FILL  FILL_199
timestamp 1710899220
transform 1 0 2640 0 -1 2170
box -8 -3 16 105
use FILL  FILL_200
timestamp 1710899220
transform 1 0 2632 0 -1 2170
box -8 -3 16 105
use FILL  FILL_201
timestamp 1710899220
transform 1 0 2624 0 -1 2170
box -8 -3 16 105
use FILL  FILL_202
timestamp 1710899220
transform 1 0 2616 0 -1 2170
box -8 -3 16 105
use FILL  FILL_203
timestamp 1710899220
transform 1 0 2608 0 -1 2170
box -8 -3 16 105
use FILL  FILL_204
timestamp 1710899220
transform 1 0 2600 0 -1 2170
box -8 -3 16 105
use FILL  FILL_205
timestamp 1710899220
transform 1 0 2592 0 -1 2170
box -8 -3 16 105
use FILL  FILL_206
timestamp 1710899220
transform 1 0 2584 0 -1 2170
box -8 -3 16 105
use FILL  FILL_207
timestamp 1710899220
transform 1 0 2576 0 -1 2170
box -8 -3 16 105
use FILL  FILL_208
timestamp 1710899220
transform 1 0 2568 0 -1 2170
box -8 -3 16 105
use FILL  FILL_209
timestamp 1710899220
transform 1 0 2560 0 -1 2170
box -8 -3 16 105
use FILL  FILL_210
timestamp 1710899220
transform 1 0 2552 0 -1 2170
box -8 -3 16 105
use FILL  FILL_211
timestamp 1710899220
transform 1 0 2544 0 -1 2170
box -8 -3 16 105
use FILL  FILL_212
timestamp 1710899220
transform 1 0 2536 0 -1 2170
box -8 -3 16 105
use FILL  FILL_213
timestamp 1710899220
transform 1 0 2528 0 -1 2170
box -8 -3 16 105
use FILL  FILL_214
timestamp 1710899220
transform 1 0 2520 0 -1 2170
box -8 -3 16 105
use FILL  FILL_215
timestamp 1710899220
transform 1 0 2512 0 -1 2170
box -8 -3 16 105
use FILL  FILL_216
timestamp 1710899220
transform 1 0 2504 0 -1 2170
box -8 -3 16 105
use FILL  FILL_217
timestamp 1710899220
transform 1 0 2400 0 -1 2170
box -8 -3 16 105
use FILL  FILL_218
timestamp 1710899220
transform 1 0 2376 0 -1 2170
box -8 -3 16 105
use FILL  FILL_219
timestamp 1710899220
transform 1 0 2368 0 -1 2170
box -8 -3 16 105
use FILL  FILL_220
timestamp 1710899220
transform 1 0 2360 0 -1 2170
box -8 -3 16 105
use FILL  FILL_221
timestamp 1710899220
transform 1 0 2352 0 -1 2170
box -8 -3 16 105
use FILL  FILL_222
timestamp 1710899220
transform 1 0 2264 0 -1 2170
box -8 -3 16 105
use FILL  FILL_223
timestamp 1710899220
transform 1 0 2256 0 -1 2170
box -8 -3 16 105
use FILL  FILL_224
timestamp 1710899220
transform 1 0 2016 0 -1 2170
box -8 -3 16 105
use FILL  FILL_225
timestamp 1710899220
transform 1 0 1928 0 -1 2170
box -8 -3 16 105
use FILL  FILL_226
timestamp 1710899220
transform 1 0 1864 0 -1 2170
box -8 -3 16 105
use FILL  FILL_227
timestamp 1710899220
transform 1 0 1856 0 -1 2170
box -8 -3 16 105
use FILL  FILL_228
timestamp 1710899220
transform 1 0 1752 0 -1 2170
box -8 -3 16 105
use FILL  FILL_229
timestamp 1710899220
transform 1 0 1664 0 -1 2170
box -8 -3 16 105
use FILL  FILL_230
timestamp 1710899220
transform 1 0 1592 0 -1 2170
box -8 -3 16 105
use FILL  FILL_231
timestamp 1710899220
transform 1 0 1456 0 -1 2170
box -8 -3 16 105
use FILL  FILL_232
timestamp 1710899220
transform 1 0 1448 0 -1 2170
box -8 -3 16 105
use FILL  FILL_233
timestamp 1710899220
transform 1 0 1376 0 -1 2170
box -8 -3 16 105
use FILL  FILL_234
timestamp 1710899220
transform 1 0 1280 0 -1 2170
box -8 -3 16 105
use FILL  FILL_235
timestamp 1710899220
transform 1 0 1272 0 -1 2170
box -8 -3 16 105
use FILL  FILL_236
timestamp 1710899220
transform 1 0 1200 0 -1 2170
box -8 -3 16 105
use FILL  FILL_237
timestamp 1710899220
transform 1 0 1112 0 -1 2170
box -8 -3 16 105
use FILL  FILL_238
timestamp 1710899220
transform 1 0 1104 0 -1 2170
box -8 -3 16 105
use FILL  FILL_239
timestamp 1710899220
transform 1 0 1096 0 -1 2170
box -8 -3 16 105
use FILL  FILL_240
timestamp 1710899220
transform 1 0 1064 0 -1 2170
box -8 -3 16 105
use FILL  FILL_241
timestamp 1710899220
transform 1 0 1056 0 -1 2170
box -8 -3 16 105
use FILL  FILL_242
timestamp 1710899220
transform 1 0 1048 0 -1 2170
box -8 -3 16 105
use FILL  FILL_243
timestamp 1710899220
transform 1 0 920 0 -1 2170
box -8 -3 16 105
use FILL  FILL_244
timestamp 1710899220
transform 1 0 912 0 -1 2170
box -8 -3 16 105
use FILL  FILL_245
timestamp 1710899220
transform 1 0 904 0 -1 2170
box -8 -3 16 105
use FILL  FILL_246
timestamp 1710899220
transform 1 0 896 0 -1 2170
box -8 -3 16 105
use FILL  FILL_247
timestamp 1710899220
transform 1 0 768 0 -1 2170
box -8 -3 16 105
use FILL  FILL_248
timestamp 1710899220
transform 1 0 760 0 -1 2170
box -8 -3 16 105
use FILL  FILL_249
timestamp 1710899220
transform 1 0 752 0 -1 2170
box -8 -3 16 105
use FILL  FILL_250
timestamp 1710899220
transform 1 0 744 0 -1 2170
box -8 -3 16 105
use FILL  FILL_251
timestamp 1710899220
transform 1 0 736 0 -1 2170
box -8 -3 16 105
use FILL  FILL_252
timestamp 1710899220
transform 1 0 728 0 -1 2170
box -8 -3 16 105
use FILL  FILL_253
timestamp 1710899220
transform 1 0 672 0 -1 2170
box -8 -3 16 105
use FILL  FILL_254
timestamp 1710899220
transform 1 0 664 0 -1 2170
box -8 -3 16 105
use FILL  FILL_255
timestamp 1710899220
transform 1 0 656 0 -1 2170
box -8 -3 16 105
use FILL  FILL_256
timestamp 1710899220
transform 1 0 648 0 -1 2170
box -8 -3 16 105
use FILL  FILL_257
timestamp 1710899220
transform 1 0 640 0 -1 2170
box -8 -3 16 105
use FILL  FILL_258
timestamp 1710899220
transform 1 0 512 0 -1 2170
box -8 -3 16 105
use FILL  FILL_259
timestamp 1710899220
transform 1 0 504 0 -1 2170
box -8 -3 16 105
use FILL  FILL_260
timestamp 1710899220
transform 1 0 496 0 -1 2170
box -8 -3 16 105
use FILL  FILL_261
timestamp 1710899220
transform 1 0 368 0 -1 2170
box -8 -3 16 105
use FILL  FILL_262
timestamp 1710899220
transform 1 0 360 0 -1 2170
box -8 -3 16 105
use FILL  FILL_263
timestamp 1710899220
transform 1 0 352 0 -1 2170
box -8 -3 16 105
use FILL  FILL_264
timestamp 1710899220
transform 1 0 224 0 -1 2170
box -8 -3 16 105
use FILL  FILL_265
timestamp 1710899220
transform 1 0 96 0 -1 2170
box -8 -3 16 105
use FILL  FILL_266
timestamp 1710899220
transform 1 0 88 0 -1 2170
box -8 -3 16 105
use FILL  FILL_267
timestamp 1710899220
transform 1 0 80 0 -1 2170
box -8 -3 16 105
use FILL  FILL_268
timestamp 1710899220
transform 1 0 72 0 -1 2170
box -8 -3 16 105
use FILL  FILL_269
timestamp 1710899220
transform 1 0 2432 0 1 1970
box -8 -3 16 105
use FILL  FILL_270
timestamp 1710899220
transform 1 0 2328 0 1 1970
box -8 -3 16 105
use FILL  FILL_271
timestamp 1710899220
transform 1 0 2264 0 1 1970
box -8 -3 16 105
use FILL  FILL_272
timestamp 1710899220
transform 1 0 2256 0 1 1970
box -8 -3 16 105
use FILL  FILL_273
timestamp 1710899220
transform 1 0 2248 0 1 1970
box -8 -3 16 105
use FILL  FILL_274
timestamp 1710899220
transform 1 0 2160 0 1 1970
box -8 -3 16 105
use FILL  FILL_275
timestamp 1710899220
transform 1 0 2072 0 1 1970
box -8 -3 16 105
use FILL  FILL_276
timestamp 1710899220
transform 1 0 2064 0 1 1970
box -8 -3 16 105
use FILL  FILL_277
timestamp 1710899220
transform 1 0 2056 0 1 1970
box -8 -3 16 105
use FILL  FILL_278
timestamp 1710899220
transform 1 0 2048 0 1 1970
box -8 -3 16 105
use FILL  FILL_279
timestamp 1710899220
transform 1 0 1808 0 1 1970
box -8 -3 16 105
use FILL  FILL_280
timestamp 1710899220
transform 1 0 1800 0 1 1970
box -8 -3 16 105
use FILL  FILL_281
timestamp 1710899220
transform 1 0 1792 0 1 1970
box -8 -3 16 105
use FILL  FILL_282
timestamp 1710899220
transform 1 0 1784 0 1 1970
box -8 -3 16 105
use FILL  FILL_283
timestamp 1710899220
transform 1 0 1776 0 1 1970
box -8 -3 16 105
use FILL  FILL_284
timestamp 1710899220
transform 1 0 1768 0 1 1970
box -8 -3 16 105
use FILL  FILL_285
timestamp 1710899220
transform 1 0 1760 0 1 1970
box -8 -3 16 105
use FILL  FILL_286
timestamp 1710899220
transform 1 0 1752 0 1 1970
box -8 -3 16 105
use FILL  FILL_287
timestamp 1710899220
transform 1 0 1744 0 1 1970
box -8 -3 16 105
use FILL  FILL_288
timestamp 1710899220
transform 1 0 1736 0 1 1970
box -8 -3 16 105
use FILL  FILL_289
timestamp 1710899220
transform 1 0 1728 0 1 1970
box -8 -3 16 105
use FILL  FILL_290
timestamp 1710899220
transform 1 0 1720 0 1 1970
box -8 -3 16 105
use FILL  FILL_291
timestamp 1710899220
transform 1 0 1712 0 1 1970
box -8 -3 16 105
use FILL  FILL_292
timestamp 1710899220
transform 1 0 1704 0 1 1970
box -8 -3 16 105
use FILL  FILL_293
timestamp 1710899220
transform 1 0 1696 0 1 1970
box -8 -3 16 105
use FILL  FILL_294
timestamp 1710899220
transform 1 0 1688 0 1 1970
box -8 -3 16 105
use FILL  FILL_295
timestamp 1710899220
transform 1 0 1584 0 1 1970
box -8 -3 16 105
use FILL  FILL_296
timestamp 1710899220
transform 1 0 1576 0 1 1970
box -8 -3 16 105
use FILL  FILL_297
timestamp 1710899220
transform 1 0 1496 0 1 1970
box -8 -3 16 105
use FILL  FILL_298
timestamp 1710899220
transform 1 0 1392 0 1 1970
box -8 -3 16 105
use FILL  FILL_299
timestamp 1710899220
transform 1 0 1216 0 1 1970
box -8 -3 16 105
use FILL  FILL_300
timestamp 1710899220
transform 1 0 1208 0 1 1970
box -8 -3 16 105
use FILL  FILL_301
timestamp 1710899220
transform 1 0 1200 0 1 1970
box -8 -3 16 105
use FILL  FILL_302
timestamp 1710899220
transform 1 0 1024 0 1 1970
box -8 -3 16 105
use FILL  FILL_303
timestamp 1710899220
transform 1 0 952 0 1 1970
box -8 -3 16 105
use FILL  FILL_304
timestamp 1710899220
transform 1 0 944 0 1 1970
box -8 -3 16 105
use FILL  FILL_305
timestamp 1710899220
transform 1 0 824 0 1 1970
box -8 -3 16 105
use FILL  FILL_306
timestamp 1710899220
transform 1 0 296 0 1 1970
box -8 -3 16 105
use FILL  FILL_307
timestamp 1710899220
transform 1 0 288 0 1 1970
box -8 -3 16 105
use FILL  FILL_308
timestamp 1710899220
transform 1 0 224 0 1 1970
box -8 -3 16 105
use FILL  FILL_309
timestamp 1710899220
transform 1 0 216 0 1 1970
box -8 -3 16 105
use FILL  FILL_310
timestamp 1710899220
transform 1 0 208 0 1 1970
box -8 -3 16 105
use FILL  FILL_311
timestamp 1710899220
transform 1 0 200 0 1 1970
box -8 -3 16 105
use FILL  FILL_312
timestamp 1710899220
transform 1 0 192 0 1 1970
box -8 -3 16 105
use FILL  FILL_313
timestamp 1710899220
transform 1 0 184 0 1 1970
box -8 -3 16 105
use FILL  FILL_314
timestamp 1710899220
transform 1 0 176 0 1 1970
box -8 -3 16 105
use FILL  FILL_315
timestamp 1710899220
transform 1 0 168 0 1 1970
box -8 -3 16 105
use FILL  FILL_316
timestamp 1710899220
transform 1 0 160 0 1 1970
box -8 -3 16 105
use FILL  FILL_317
timestamp 1710899220
transform 1 0 152 0 1 1970
box -8 -3 16 105
use FILL  FILL_318
timestamp 1710899220
transform 1 0 144 0 1 1970
box -8 -3 16 105
use FILL  FILL_319
timestamp 1710899220
transform 1 0 136 0 1 1970
box -8 -3 16 105
use FILL  FILL_320
timestamp 1710899220
transform 1 0 128 0 1 1970
box -8 -3 16 105
use FILL  FILL_321
timestamp 1710899220
transform 1 0 120 0 1 1970
box -8 -3 16 105
use FILL  FILL_322
timestamp 1710899220
transform 1 0 112 0 1 1970
box -8 -3 16 105
use FILL  FILL_323
timestamp 1710899220
transform 1 0 104 0 1 1970
box -8 -3 16 105
use FILL  FILL_324
timestamp 1710899220
transform 1 0 96 0 1 1970
box -8 -3 16 105
use FILL  FILL_325
timestamp 1710899220
transform 1 0 88 0 1 1970
box -8 -3 16 105
use FILL  FILL_326
timestamp 1710899220
transform 1 0 80 0 1 1970
box -8 -3 16 105
use FILL  FILL_327
timestamp 1710899220
transform 1 0 72 0 1 1970
box -8 -3 16 105
use FILL  FILL_328
timestamp 1710899220
transform 1 0 2416 0 -1 1970
box -8 -3 16 105
use FILL  FILL_329
timestamp 1710899220
transform 1 0 2408 0 -1 1970
box -8 -3 16 105
use FILL  FILL_330
timestamp 1710899220
transform 1 0 2400 0 -1 1970
box -8 -3 16 105
use FILL  FILL_331
timestamp 1710899220
transform 1 0 2392 0 -1 1970
box -8 -3 16 105
use FILL  FILL_332
timestamp 1710899220
transform 1 0 2384 0 -1 1970
box -8 -3 16 105
use FILL  FILL_333
timestamp 1710899220
transform 1 0 2376 0 -1 1970
box -8 -3 16 105
use FILL  FILL_334
timestamp 1710899220
transform 1 0 2368 0 -1 1970
box -8 -3 16 105
use FILL  FILL_335
timestamp 1710899220
transform 1 0 2360 0 -1 1970
box -8 -3 16 105
use FILL  FILL_336
timestamp 1710899220
transform 1 0 2352 0 -1 1970
box -8 -3 16 105
use FILL  FILL_337
timestamp 1710899220
transform 1 0 2344 0 -1 1970
box -8 -3 16 105
use FILL  FILL_338
timestamp 1710899220
transform 1 0 2336 0 -1 1970
box -8 -3 16 105
use FILL  FILL_339
timestamp 1710899220
transform 1 0 2232 0 -1 1970
box -8 -3 16 105
use FILL  FILL_340
timestamp 1710899220
transform 1 0 2224 0 -1 1970
box -8 -3 16 105
use FILL  FILL_341
timestamp 1710899220
transform 1 0 2216 0 -1 1970
box -8 -3 16 105
use FILL  FILL_342
timestamp 1710899220
transform 1 0 2152 0 -1 1970
box -8 -3 16 105
use FILL  FILL_343
timestamp 1710899220
transform 1 0 2144 0 -1 1970
box -8 -3 16 105
use FILL  FILL_344
timestamp 1710899220
transform 1 0 2080 0 -1 1970
box -8 -3 16 105
use FILL  FILL_345
timestamp 1710899220
transform 1 0 1976 0 -1 1970
box -8 -3 16 105
use FILL  FILL_346
timestamp 1710899220
transform 1 0 1968 0 -1 1970
box -8 -3 16 105
use FILL  FILL_347
timestamp 1710899220
transform 1 0 1960 0 -1 1970
box -8 -3 16 105
use FILL  FILL_348
timestamp 1710899220
transform 1 0 1952 0 -1 1970
box -8 -3 16 105
use FILL  FILL_349
timestamp 1710899220
transform 1 0 1944 0 -1 1970
box -8 -3 16 105
use FILL  FILL_350
timestamp 1710899220
transform 1 0 1936 0 -1 1970
box -8 -3 16 105
use FILL  FILL_351
timestamp 1710899220
transform 1 0 1928 0 -1 1970
box -8 -3 16 105
use FILL  FILL_352
timestamp 1710899220
transform 1 0 1920 0 -1 1970
box -8 -3 16 105
use FILL  FILL_353
timestamp 1710899220
transform 1 0 1912 0 -1 1970
box -8 -3 16 105
use FILL  FILL_354
timestamp 1710899220
transform 1 0 1904 0 -1 1970
box -8 -3 16 105
use FILL  FILL_355
timestamp 1710899220
transform 1 0 1896 0 -1 1970
box -8 -3 16 105
use FILL  FILL_356
timestamp 1710899220
transform 1 0 1888 0 -1 1970
box -8 -3 16 105
use FILL  FILL_357
timestamp 1710899220
transform 1 0 1880 0 -1 1970
box -8 -3 16 105
use FILL  FILL_358
timestamp 1710899220
transform 1 0 1872 0 -1 1970
box -8 -3 16 105
use FILL  FILL_359
timestamp 1710899220
transform 1 0 1864 0 -1 1970
box -8 -3 16 105
use FILL  FILL_360
timestamp 1710899220
transform 1 0 1856 0 -1 1970
box -8 -3 16 105
use FILL  FILL_361
timestamp 1710899220
transform 1 0 1848 0 -1 1970
box -8 -3 16 105
use FILL  FILL_362
timestamp 1710899220
transform 1 0 1840 0 -1 1970
box -8 -3 16 105
use FILL  FILL_363
timestamp 1710899220
transform 1 0 1832 0 -1 1970
box -8 -3 16 105
use FILL  FILL_364
timestamp 1710899220
transform 1 0 1824 0 -1 1970
box -8 -3 16 105
use FILL  FILL_365
timestamp 1710899220
transform 1 0 1816 0 -1 1970
box -8 -3 16 105
use FILL  FILL_366
timestamp 1710899220
transform 1 0 1808 0 -1 1970
box -8 -3 16 105
use FILL  FILL_367
timestamp 1710899220
transform 1 0 1800 0 -1 1970
box -8 -3 16 105
use FILL  FILL_368
timestamp 1710899220
transform 1 0 1792 0 -1 1970
box -8 -3 16 105
use FILL  FILL_369
timestamp 1710899220
transform 1 0 1784 0 -1 1970
box -8 -3 16 105
use FILL  FILL_370
timestamp 1710899220
transform 1 0 1776 0 -1 1970
box -8 -3 16 105
use FILL  FILL_371
timestamp 1710899220
transform 1 0 1768 0 -1 1970
box -8 -3 16 105
use FILL  FILL_372
timestamp 1710899220
transform 1 0 1664 0 -1 1970
box -8 -3 16 105
use FILL  FILL_373
timestamp 1710899220
transform 1 0 1656 0 -1 1970
box -8 -3 16 105
use FILL  FILL_374
timestamp 1710899220
transform 1 0 1600 0 -1 1970
box -8 -3 16 105
use FILL  FILL_375
timestamp 1710899220
transform 1 0 1568 0 -1 1970
box -8 -3 16 105
use FILL  FILL_376
timestamp 1710899220
transform 1 0 1560 0 -1 1970
box -8 -3 16 105
use FILL  FILL_377
timestamp 1710899220
transform 1 0 1520 0 -1 1970
box -8 -3 16 105
use FILL  FILL_378
timestamp 1710899220
transform 1 0 1488 0 -1 1970
box -8 -3 16 105
use FILL  FILL_379
timestamp 1710899220
transform 1 0 1480 0 -1 1970
box -8 -3 16 105
use FILL  FILL_380
timestamp 1710899220
transform 1 0 1472 0 -1 1970
box -8 -3 16 105
use FILL  FILL_381
timestamp 1710899220
transform 1 0 1464 0 -1 1970
box -8 -3 16 105
use FILL  FILL_382
timestamp 1710899220
transform 1 0 1456 0 -1 1970
box -8 -3 16 105
use FILL  FILL_383
timestamp 1710899220
transform 1 0 1392 0 -1 1970
box -8 -3 16 105
use FILL  FILL_384
timestamp 1710899220
transform 1 0 1384 0 -1 1970
box -8 -3 16 105
use FILL  FILL_385
timestamp 1710899220
transform 1 0 1376 0 -1 1970
box -8 -3 16 105
use FILL  FILL_386
timestamp 1710899220
transform 1 0 1368 0 -1 1970
box -8 -3 16 105
use FILL  FILL_387
timestamp 1710899220
transform 1 0 1304 0 -1 1970
box -8 -3 16 105
use FILL  FILL_388
timestamp 1710899220
transform 1 0 1296 0 -1 1970
box -8 -3 16 105
use FILL  FILL_389
timestamp 1710899220
transform 1 0 1288 0 -1 1970
box -8 -3 16 105
use FILL  FILL_390
timestamp 1710899220
transform 1 0 1184 0 -1 1970
box -8 -3 16 105
use FILL  FILL_391
timestamp 1710899220
transform 1 0 1112 0 -1 1970
box -8 -3 16 105
use FILL  FILL_392
timestamp 1710899220
transform 1 0 1104 0 -1 1970
box -8 -3 16 105
use FILL  FILL_393
timestamp 1710899220
transform 1 0 1096 0 -1 1970
box -8 -3 16 105
use FILL  FILL_394
timestamp 1710899220
transform 1 0 1088 0 -1 1970
box -8 -3 16 105
use FILL  FILL_395
timestamp 1710899220
transform 1 0 928 0 -1 1970
box -8 -3 16 105
use FILL  FILL_396
timestamp 1710899220
transform 1 0 920 0 -1 1970
box -8 -3 16 105
use FILL  FILL_397
timestamp 1710899220
transform 1 0 760 0 -1 1970
box -8 -3 16 105
use FILL  FILL_398
timestamp 1710899220
transform 1 0 752 0 -1 1970
box -8 -3 16 105
use FILL  FILL_399
timestamp 1710899220
transform 1 0 744 0 -1 1970
box -8 -3 16 105
use FILL  FILL_400
timestamp 1710899220
transform 1 0 736 0 -1 1970
box -8 -3 16 105
use FILL  FILL_401
timestamp 1710899220
transform 1 0 728 0 -1 1970
box -8 -3 16 105
use FILL  FILL_402
timestamp 1710899220
transform 1 0 720 0 -1 1970
box -8 -3 16 105
use FILL  FILL_403
timestamp 1710899220
transform 1 0 696 0 -1 1970
box -8 -3 16 105
use FILL  FILL_404
timestamp 1710899220
transform 1 0 632 0 -1 1970
box -8 -3 16 105
use FILL  FILL_405
timestamp 1710899220
transform 1 0 624 0 -1 1970
box -8 -3 16 105
use FILL  FILL_406
timestamp 1710899220
transform 1 0 520 0 -1 1970
box -8 -3 16 105
use FILL  FILL_407
timestamp 1710899220
transform 1 0 512 0 -1 1970
box -8 -3 16 105
use FILL  FILL_408
timestamp 1710899220
transform 1 0 504 0 -1 1970
box -8 -3 16 105
use FILL  FILL_409
timestamp 1710899220
transform 1 0 448 0 -1 1970
box -8 -3 16 105
use FILL  FILL_410
timestamp 1710899220
transform 1 0 296 0 -1 1970
box -8 -3 16 105
use FILL  FILL_411
timestamp 1710899220
transform 1 0 120 0 -1 1970
box -8 -3 16 105
use FILL  FILL_412
timestamp 1710899220
transform 1 0 112 0 -1 1970
box -8 -3 16 105
use FILL  FILL_413
timestamp 1710899220
transform 1 0 104 0 -1 1970
box -8 -3 16 105
use FILL  FILL_414
timestamp 1710899220
transform 1 0 96 0 -1 1970
box -8 -3 16 105
use FILL  FILL_415
timestamp 1710899220
transform 1 0 88 0 -1 1970
box -8 -3 16 105
use FILL  FILL_416
timestamp 1710899220
transform 1 0 80 0 -1 1970
box -8 -3 16 105
use FILL  FILL_417
timestamp 1710899220
transform 1 0 72 0 -1 1970
box -8 -3 16 105
use FILL  FILL_418
timestamp 1710899220
transform 1 0 1992 0 1 1770
box -8 -3 16 105
use FILL  FILL_419
timestamp 1710899220
transform 1 0 1984 0 1 1770
box -8 -3 16 105
use FILL  FILL_420
timestamp 1710899220
transform 1 0 1976 0 1 1770
box -8 -3 16 105
use FILL  FILL_421
timestamp 1710899220
transform 1 0 1968 0 1 1770
box -8 -3 16 105
use FILL  FILL_422
timestamp 1710899220
transform 1 0 1960 0 1 1770
box -8 -3 16 105
use FILL  FILL_423
timestamp 1710899220
transform 1 0 1952 0 1 1770
box -8 -3 16 105
use FILL  FILL_424
timestamp 1710899220
transform 1 0 1864 0 1 1770
box -8 -3 16 105
use FILL  FILL_425
timestamp 1710899220
transform 1 0 1856 0 1 1770
box -8 -3 16 105
use FILL  FILL_426
timestamp 1710899220
transform 1 0 1752 0 1 1770
box -8 -3 16 105
use FILL  FILL_427
timestamp 1710899220
transform 1 0 1672 0 1 1770
box -8 -3 16 105
use FILL  FILL_428
timestamp 1710899220
transform 1 0 1592 0 1 1770
box -8 -3 16 105
use FILL  FILL_429
timestamp 1710899220
transform 1 0 1192 0 1 1770
box -8 -3 16 105
use FILL  FILL_430
timestamp 1710899220
transform 1 0 1056 0 1 1770
box -8 -3 16 105
use FILL  FILL_431
timestamp 1710899220
transform 1 0 1048 0 1 1770
box -8 -3 16 105
use FILL  FILL_432
timestamp 1710899220
transform 1 0 968 0 1 1770
box -8 -3 16 105
use FILL  FILL_433
timestamp 1710899220
transform 1 0 864 0 1 1770
box -8 -3 16 105
use FILL  FILL_434
timestamp 1710899220
transform 1 0 784 0 1 1770
box -8 -3 16 105
use FILL  FILL_435
timestamp 1710899220
transform 1 0 680 0 1 1770
box -8 -3 16 105
use FILL  FILL_436
timestamp 1710899220
transform 1 0 672 0 1 1770
box -8 -3 16 105
use FILL  FILL_437
timestamp 1710899220
transform 1 0 592 0 1 1770
box -8 -3 16 105
use FILL  FILL_438
timestamp 1710899220
transform 1 0 584 0 1 1770
box -8 -3 16 105
use FILL  FILL_439
timestamp 1710899220
transform 1 0 576 0 1 1770
box -8 -3 16 105
use FILL  FILL_440
timestamp 1710899220
transform 1 0 568 0 1 1770
box -8 -3 16 105
use FILL  FILL_441
timestamp 1710899220
transform 1 0 560 0 1 1770
box -8 -3 16 105
use FILL  FILL_442
timestamp 1710899220
transform 1 0 456 0 1 1770
box -8 -3 16 105
use FILL  FILL_443
timestamp 1710899220
transform 1 0 448 0 1 1770
box -8 -3 16 105
use FILL  FILL_444
timestamp 1710899220
transform 1 0 440 0 1 1770
box -8 -3 16 105
use FILL  FILL_445
timestamp 1710899220
transform 1 0 432 0 1 1770
box -8 -3 16 105
use FILL  FILL_446
timestamp 1710899220
transform 1 0 424 0 1 1770
box -8 -3 16 105
use FILL  FILL_447
timestamp 1710899220
transform 1 0 416 0 1 1770
box -8 -3 16 105
use FILL  FILL_448
timestamp 1710899220
transform 1 0 408 0 1 1770
box -8 -3 16 105
use FILL  FILL_449
timestamp 1710899220
transform 1 0 400 0 1 1770
box -8 -3 16 105
use FILL  FILL_450
timestamp 1710899220
transform 1 0 392 0 1 1770
box -8 -3 16 105
use FILL  FILL_451
timestamp 1710899220
transform 1 0 384 0 1 1770
box -8 -3 16 105
use FILL  FILL_452
timestamp 1710899220
transform 1 0 376 0 1 1770
box -8 -3 16 105
use FILL  FILL_453
timestamp 1710899220
transform 1 0 368 0 1 1770
box -8 -3 16 105
use FILL  FILL_454
timestamp 1710899220
transform 1 0 360 0 1 1770
box -8 -3 16 105
use FILL  FILL_455
timestamp 1710899220
transform 1 0 352 0 1 1770
box -8 -3 16 105
use FILL  FILL_456
timestamp 1710899220
transform 1 0 344 0 1 1770
box -8 -3 16 105
use FILL  FILL_457
timestamp 1710899220
transform 1 0 336 0 1 1770
box -8 -3 16 105
use FILL  FILL_458
timestamp 1710899220
transform 1 0 328 0 1 1770
box -8 -3 16 105
use FILL  FILL_459
timestamp 1710899220
transform 1 0 320 0 1 1770
box -8 -3 16 105
use FILL  FILL_460
timestamp 1710899220
transform 1 0 312 0 1 1770
box -8 -3 16 105
use FILL  FILL_461
timestamp 1710899220
transform 1 0 304 0 1 1770
box -8 -3 16 105
use FILL  FILL_462
timestamp 1710899220
transform 1 0 296 0 1 1770
box -8 -3 16 105
use FILL  FILL_463
timestamp 1710899220
transform 1 0 288 0 1 1770
box -8 -3 16 105
use FILL  FILL_464
timestamp 1710899220
transform 1 0 280 0 1 1770
box -8 -3 16 105
use FILL  FILL_465
timestamp 1710899220
transform 1 0 272 0 1 1770
box -8 -3 16 105
use FILL  FILL_466
timestamp 1710899220
transform 1 0 264 0 1 1770
box -8 -3 16 105
use FILL  FILL_467
timestamp 1710899220
transform 1 0 256 0 1 1770
box -8 -3 16 105
use FILL  FILL_468
timestamp 1710899220
transform 1 0 248 0 1 1770
box -8 -3 16 105
use FILL  FILL_469
timestamp 1710899220
transform 1 0 240 0 1 1770
box -8 -3 16 105
use FILL  FILL_470
timestamp 1710899220
transform 1 0 232 0 1 1770
box -8 -3 16 105
use FILL  FILL_471
timestamp 1710899220
transform 1 0 224 0 1 1770
box -8 -3 16 105
use FILL  FILL_472
timestamp 1710899220
transform 1 0 216 0 1 1770
box -8 -3 16 105
use FILL  FILL_473
timestamp 1710899220
transform 1 0 208 0 1 1770
box -8 -3 16 105
use FILL  FILL_474
timestamp 1710899220
transform 1 0 200 0 1 1770
box -8 -3 16 105
use FILL  FILL_475
timestamp 1710899220
transform 1 0 192 0 1 1770
box -8 -3 16 105
use FILL  FILL_476
timestamp 1710899220
transform 1 0 184 0 1 1770
box -8 -3 16 105
use FILL  FILL_477
timestamp 1710899220
transform 1 0 176 0 1 1770
box -8 -3 16 105
use FILL  FILL_478
timestamp 1710899220
transform 1 0 168 0 1 1770
box -8 -3 16 105
use FILL  FILL_479
timestamp 1710899220
transform 1 0 160 0 1 1770
box -8 -3 16 105
use FILL  FILL_480
timestamp 1710899220
transform 1 0 152 0 1 1770
box -8 -3 16 105
use FILL  FILL_481
timestamp 1710899220
transform 1 0 144 0 1 1770
box -8 -3 16 105
use FILL  FILL_482
timestamp 1710899220
transform 1 0 136 0 1 1770
box -8 -3 16 105
use FILL  FILL_483
timestamp 1710899220
transform 1 0 128 0 1 1770
box -8 -3 16 105
use FILL  FILL_484
timestamp 1710899220
transform 1 0 120 0 1 1770
box -8 -3 16 105
use FILL  FILL_485
timestamp 1710899220
transform 1 0 112 0 1 1770
box -8 -3 16 105
use FILL  FILL_486
timestamp 1710899220
transform 1 0 104 0 1 1770
box -8 -3 16 105
use FILL  FILL_487
timestamp 1710899220
transform 1 0 96 0 1 1770
box -8 -3 16 105
use FILL  FILL_488
timestamp 1710899220
transform 1 0 88 0 1 1770
box -8 -3 16 105
use FILL  FILL_489
timestamp 1710899220
transform 1 0 80 0 1 1770
box -8 -3 16 105
use FILL  FILL_490
timestamp 1710899220
transform 1 0 72 0 1 1770
box -8 -3 16 105
use FILL  FILL_491
timestamp 1710899220
transform 1 0 1784 0 -1 1770
box -8 -3 16 105
use FILL  FILL_492
timestamp 1710899220
transform 1 0 1680 0 -1 1770
box -8 -3 16 105
use FILL  FILL_493
timestamp 1710899220
transform 1 0 1672 0 -1 1770
box -8 -3 16 105
use FILL  FILL_494
timestamp 1710899220
transform 1 0 1616 0 -1 1770
box -8 -3 16 105
use FILL  FILL_495
timestamp 1710899220
transform 1 0 1544 0 -1 1770
box -8 -3 16 105
use FILL  FILL_496
timestamp 1710899220
transform 1 0 1472 0 -1 1770
box -8 -3 16 105
use FILL  FILL_497
timestamp 1710899220
transform 1 0 1464 0 -1 1770
box -8 -3 16 105
use FILL  FILL_498
timestamp 1710899220
transform 1 0 1432 0 -1 1770
box -8 -3 16 105
use FILL  FILL_499
timestamp 1710899220
transform 1 0 1424 0 -1 1770
box -8 -3 16 105
use FILL  FILL_500
timestamp 1710899220
transform 1 0 1352 0 -1 1770
box -8 -3 16 105
use FILL  FILL_501
timestamp 1710899220
transform 1 0 1344 0 -1 1770
box -8 -3 16 105
use FILL  FILL_502
timestamp 1710899220
transform 1 0 1288 0 -1 1770
box -8 -3 16 105
use FILL  FILL_503
timestamp 1710899220
transform 1 0 1248 0 -1 1770
box -8 -3 16 105
use FILL  FILL_504
timestamp 1710899220
transform 1 0 1208 0 -1 1770
box -8 -3 16 105
use FILL  FILL_505
timestamp 1710899220
transform 1 0 1184 0 -1 1770
box -8 -3 16 105
use FILL  FILL_506
timestamp 1710899220
transform 1 0 1112 0 -1 1770
box -8 -3 16 105
use FILL  FILL_507
timestamp 1710899220
transform 1 0 1104 0 -1 1770
box -8 -3 16 105
use FILL  FILL_508
timestamp 1710899220
transform 1 0 1032 0 -1 1770
box -8 -3 16 105
use FILL  FILL_509
timestamp 1710899220
transform 1 0 1024 0 -1 1770
box -8 -3 16 105
use FILL  FILL_510
timestamp 1710899220
transform 1 0 960 0 -1 1770
box -8 -3 16 105
use FILL  FILL_511
timestamp 1710899220
transform 1 0 800 0 -1 1770
box -8 -3 16 105
use FILL  FILL_512
timestamp 1710899220
transform 1 0 792 0 -1 1770
box -8 -3 16 105
use FILL  FILL_513
timestamp 1710899220
transform 1 0 784 0 -1 1770
box -8 -3 16 105
use FILL  FILL_514
timestamp 1710899220
transform 1 0 720 0 -1 1770
box -8 -3 16 105
use FILL  FILL_515
timestamp 1710899220
transform 1 0 712 0 -1 1770
box -8 -3 16 105
use FILL  FILL_516
timestamp 1710899220
transform 1 0 624 0 -1 1770
box -8 -3 16 105
use FILL  FILL_517
timestamp 1710899220
transform 1 0 544 0 -1 1770
box -8 -3 16 105
use FILL  FILL_518
timestamp 1710899220
transform 1 0 496 0 -1 1770
box -8 -3 16 105
use FILL  FILL_519
timestamp 1710899220
transform 1 0 488 0 -1 1770
box -8 -3 16 105
use FILL  FILL_520
timestamp 1710899220
transform 1 0 480 0 -1 1770
box -8 -3 16 105
use FILL  FILL_521
timestamp 1710899220
transform 1 0 392 0 -1 1770
box -8 -3 16 105
use FILL  FILL_522
timestamp 1710899220
transform 1 0 304 0 -1 1770
box -8 -3 16 105
use FILL  FILL_523
timestamp 1710899220
transform 1 0 248 0 -1 1770
box -8 -3 16 105
use FILL  FILL_524
timestamp 1710899220
transform 1 0 240 0 -1 1770
box -8 -3 16 105
use FILL  FILL_525
timestamp 1710899220
transform 1 0 176 0 -1 1770
box -8 -3 16 105
use FILL  FILL_526
timestamp 1710899220
transform 1 0 168 0 -1 1770
box -8 -3 16 105
use FILL  FILL_527
timestamp 1710899220
transform 1 0 160 0 -1 1770
box -8 -3 16 105
use FILL  FILL_528
timestamp 1710899220
transform 1 0 152 0 -1 1770
box -8 -3 16 105
use FILL  FILL_529
timestamp 1710899220
transform 1 0 144 0 -1 1770
box -8 -3 16 105
use FILL  FILL_530
timestamp 1710899220
transform 1 0 136 0 -1 1770
box -8 -3 16 105
use FILL  FILL_531
timestamp 1710899220
transform 1 0 128 0 -1 1770
box -8 -3 16 105
use FILL  FILL_532
timestamp 1710899220
transform 1 0 120 0 -1 1770
box -8 -3 16 105
use FILL  FILL_533
timestamp 1710899220
transform 1 0 112 0 -1 1770
box -8 -3 16 105
use FILL  FILL_534
timestamp 1710899220
transform 1 0 104 0 -1 1770
box -8 -3 16 105
use FILL  FILL_535
timestamp 1710899220
transform 1 0 96 0 -1 1770
box -8 -3 16 105
use FILL  FILL_536
timestamp 1710899220
transform 1 0 88 0 -1 1770
box -8 -3 16 105
use FILL  FILL_537
timestamp 1710899220
transform 1 0 80 0 -1 1770
box -8 -3 16 105
use FILL  FILL_538
timestamp 1710899220
transform 1 0 72 0 -1 1770
box -8 -3 16 105
use FILL  FILL_539
timestamp 1710899220
transform 1 0 2664 0 1 1570
box -8 -3 16 105
use FILL  FILL_540
timestamp 1710899220
transform 1 0 2656 0 1 1570
box -8 -3 16 105
use FILL  FILL_541
timestamp 1710899220
transform 1 0 2648 0 1 1570
box -8 -3 16 105
use FILL  FILL_542
timestamp 1710899220
transform 1 0 2640 0 1 1570
box -8 -3 16 105
use FILL  FILL_543
timestamp 1710899220
transform 1 0 2632 0 1 1570
box -8 -3 16 105
use FILL  FILL_544
timestamp 1710899220
transform 1 0 2624 0 1 1570
box -8 -3 16 105
use FILL  FILL_545
timestamp 1710899220
transform 1 0 2600 0 1 1570
box -8 -3 16 105
use FILL  FILL_546
timestamp 1710899220
transform 1 0 2592 0 1 1570
box -8 -3 16 105
use FILL  FILL_547
timestamp 1710899220
transform 1 0 2584 0 1 1570
box -8 -3 16 105
use FILL  FILL_548
timestamp 1710899220
transform 1 0 2576 0 1 1570
box -8 -3 16 105
use FILL  FILL_549
timestamp 1710899220
transform 1 0 2568 0 1 1570
box -8 -3 16 105
use FILL  FILL_550
timestamp 1710899220
transform 1 0 2560 0 1 1570
box -8 -3 16 105
use FILL  FILL_551
timestamp 1710899220
transform 1 0 2552 0 1 1570
box -8 -3 16 105
use FILL  FILL_552
timestamp 1710899220
transform 1 0 2544 0 1 1570
box -8 -3 16 105
use FILL  FILL_553
timestamp 1710899220
transform 1 0 2536 0 1 1570
box -8 -3 16 105
use FILL  FILL_554
timestamp 1710899220
transform 1 0 2528 0 1 1570
box -8 -3 16 105
use FILL  FILL_555
timestamp 1710899220
transform 1 0 2520 0 1 1570
box -8 -3 16 105
use FILL  FILL_556
timestamp 1710899220
transform 1 0 2512 0 1 1570
box -8 -3 16 105
use FILL  FILL_557
timestamp 1710899220
transform 1 0 2504 0 1 1570
box -8 -3 16 105
use FILL  FILL_558
timestamp 1710899220
transform 1 0 2496 0 1 1570
box -8 -3 16 105
use FILL  FILL_559
timestamp 1710899220
transform 1 0 2488 0 1 1570
box -8 -3 16 105
use FILL  FILL_560
timestamp 1710899220
transform 1 0 2480 0 1 1570
box -8 -3 16 105
use FILL  FILL_561
timestamp 1710899220
transform 1 0 2472 0 1 1570
box -8 -3 16 105
use FILL  FILL_562
timestamp 1710899220
transform 1 0 2464 0 1 1570
box -8 -3 16 105
use FILL  FILL_563
timestamp 1710899220
transform 1 0 2456 0 1 1570
box -8 -3 16 105
use FILL  FILL_564
timestamp 1710899220
transform 1 0 2448 0 1 1570
box -8 -3 16 105
use FILL  FILL_565
timestamp 1710899220
transform 1 0 2440 0 1 1570
box -8 -3 16 105
use FILL  FILL_566
timestamp 1710899220
transform 1 0 2432 0 1 1570
box -8 -3 16 105
use FILL  FILL_567
timestamp 1710899220
transform 1 0 2424 0 1 1570
box -8 -3 16 105
use FILL  FILL_568
timestamp 1710899220
transform 1 0 2416 0 1 1570
box -8 -3 16 105
use FILL  FILL_569
timestamp 1710899220
transform 1 0 2408 0 1 1570
box -8 -3 16 105
use FILL  FILL_570
timestamp 1710899220
transform 1 0 2400 0 1 1570
box -8 -3 16 105
use FILL  FILL_571
timestamp 1710899220
transform 1 0 2392 0 1 1570
box -8 -3 16 105
use FILL  FILL_572
timestamp 1710899220
transform 1 0 2384 0 1 1570
box -8 -3 16 105
use FILL  FILL_573
timestamp 1710899220
transform 1 0 2376 0 1 1570
box -8 -3 16 105
use FILL  FILL_574
timestamp 1710899220
transform 1 0 2368 0 1 1570
box -8 -3 16 105
use FILL  FILL_575
timestamp 1710899220
transform 1 0 2360 0 1 1570
box -8 -3 16 105
use FILL  FILL_576
timestamp 1710899220
transform 1 0 2352 0 1 1570
box -8 -3 16 105
use FILL  FILL_577
timestamp 1710899220
transform 1 0 2344 0 1 1570
box -8 -3 16 105
use FILL  FILL_578
timestamp 1710899220
transform 1 0 2336 0 1 1570
box -8 -3 16 105
use FILL  FILL_579
timestamp 1710899220
transform 1 0 2328 0 1 1570
box -8 -3 16 105
use FILL  FILL_580
timestamp 1710899220
transform 1 0 2264 0 1 1570
box -8 -3 16 105
use FILL  FILL_581
timestamp 1710899220
transform 1 0 2256 0 1 1570
box -8 -3 16 105
use FILL  FILL_582
timestamp 1710899220
transform 1 0 2168 0 1 1570
box -8 -3 16 105
use FILL  FILL_583
timestamp 1710899220
transform 1 0 2072 0 1 1570
box -8 -3 16 105
use FILL  FILL_584
timestamp 1710899220
transform 1 0 2064 0 1 1570
box -8 -3 16 105
use FILL  FILL_585
timestamp 1710899220
transform 1 0 2056 0 1 1570
box -8 -3 16 105
use FILL  FILL_586
timestamp 1710899220
transform 1 0 1992 0 1 1570
box -8 -3 16 105
use FILL  FILL_587
timestamp 1710899220
transform 1 0 1984 0 1 1570
box -8 -3 16 105
use FILL  FILL_588
timestamp 1710899220
transform 1 0 1976 0 1 1570
box -8 -3 16 105
use FILL  FILL_589
timestamp 1710899220
transform 1 0 1968 0 1 1570
box -8 -3 16 105
use FILL  FILL_590
timestamp 1710899220
transform 1 0 1864 0 1 1570
box -8 -3 16 105
use FILL  FILL_591
timestamp 1710899220
transform 1 0 1800 0 1 1570
box -8 -3 16 105
use FILL  FILL_592
timestamp 1710899220
transform 1 0 1760 0 1 1570
box -8 -3 16 105
use FILL  FILL_593
timestamp 1710899220
transform 1 0 1752 0 1 1570
box -8 -3 16 105
use FILL  FILL_594
timestamp 1710899220
transform 1 0 1648 0 1 1570
box -8 -3 16 105
use FILL  FILL_595
timestamp 1710899220
transform 1 0 1424 0 1 1570
box -8 -3 16 105
use FILL  FILL_596
timestamp 1710899220
transform 1 0 904 0 1 1570
box -8 -3 16 105
use FILL  FILL_597
timestamp 1710899220
transform 1 0 896 0 1 1570
box -8 -3 16 105
use FILL  FILL_598
timestamp 1710899220
transform 1 0 736 0 1 1570
box -8 -3 16 105
use FILL  FILL_599
timestamp 1710899220
transform 1 0 728 0 1 1570
box -8 -3 16 105
use FILL  FILL_600
timestamp 1710899220
transform 1 0 672 0 1 1570
box -8 -3 16 105
use FILL  FILL_601
timestamp 1710899220
transform 1 0 624 0 1 1570
box -8 -3 16 105
use FILL  FILL_602
timestamp 1710899220
transform 1 0 616 0 1 1570
box -8 -3 16 105
use FILL  FILL_603
timestamp 1710899220
transform 1 0 608 0 1 1570
box -8 -3 16 105
use FILL  FILL_604
timestamp 1710899220
transform 1 0 560 0 1 1570
box -8 -3 16 105
use FILL  FILL_605
timestamp 1710899220
transform 1 0 552 0 1 1570
box -8 -3 16 105
use FILL  FILL_606
timestamp 1710899220
transform 1 0 504 0 1 1570
box -8 -3 16 105
use FILL  FILL_607
timestamp 1710899220
transform 1 0 496 0 1 1570
box -8 -3 16 105
use FILL  FILL_608
timestamp 1710899220
transform 1 0 488 0 1 1570
box -8 -3 16 105
use FILL  FILL_609
timestamp 1710899220
transform 1 0 440 0 1 1570
box -8 -3 16 105
use FILL  FILL_610
timestamp 1710899220
transform 1 0 392 0 1 1570
box -8 -3 16 105
use FILL  FILL_611
timestamp 1710899220
transform 1 0 384 0 1 1570
box -8 -3 16 105
use FILL  FILL_612
timestamp 1710899220
transform 1 0 336 0 1 1570
box -8 -3 16 105
use FILL  FILL_613
timestamp 1710899220
transform 1 0 328 0 1 1570
box -8 -3 16 105
use FILL  FILL_614
timestamp 1710899220
transform 1 0 320 0 1 1570
box -8 -3 16 105
use FILL  FILL_615
timestamp 1710899220
transform 1 0 312 0 1 1570
box -8 -3 16 105
use FILL  FILL_616
timestamp 1710899220
transform 1 0 272 0 1 1570
box -8 -3 16 105
use FILL  FILL_617
timestamp 1710899220
transform 1 0 264 0 1 1570
box -8 -3 16 105
use FILL  FILL_618
timestamp 1710899220
transform 1 0 224 0 1 1570
box -8 -3 16 105
use FILL  FILL_619
timestamp 1710899220
transform 1 0 216 0 1 1570
box -8 -3 16 105
use FILL  FILL_620
timestamp 1710899220
transform 1 0 208 0 1 1570
box -8 -3 16 105
use FILL  FILL_621
timestamp 1710899220
transform 1 0 200 0 1 1570
box -8 -3 16 105
use FILL  FILL_622
timestamp 1710899220
transform 1 0 192 0 1 1570
box -8 -3 16 105
use FILL  FILL_623
timestamp 1710899220
transform 1 0 184 0 1 1570
box -8 -3 16 105
use FILL  FILL_624
timestamp 1710899220
transform 1 0 176 0 1 1570
box -8 -3 16 105
use FILL  FILL_625
timestamp 1710899220
transform 1 0 168 0 1 1570
box -8 -3 16 105
use FILL  FILL_626
timestamp 1710899220
transform 1 0 160 0 1 1570
box -8 -3 16 105
use FILL  FILL_627
timestamp 1710899220
transform 1 0 152 0 1 1570
box -8 -3 16 105
use FILL  FILL_628
timestamp 1710899220
transform 1 0 144 0 1 1570
box -8 -3 16 105
use FILL  FILL_629
timestamp 1710899220
transform 1 0 136 0 1 1570
box -8 -3 16 105
use FILL  FILL_630
timestamp 1710899220
transform 1 0 128 0 1 1570
box -8 -3 16 105
use FILL  FILL_631
timestamp 1710899220
transform 1 0 120 0 1 1570
box -8 -3 16 105
use FILL  FILL_632
timestamp 1710899220
transform 1 0 112 0 1 1570
box -8 -3 16 105
use FILL  FILL_633
timestamp 1710899220
transform 1 0 104 0 1 1570
box -8 -3 16 105
use FILL  FILL_634
timestamp 1710899220
transform 1 0 96 0 1 1570
box -8 -3 16 105
use FILL  FILL_635
timestamp 1710899220
transform 1 0 88 0 1 1570
box -8 -3 16 105
use FILL  FILL_636
timestamp 1710899220
transform 1 0 80 0 1 1570
box -8 -3 16 105
use FILL  FILL_637
timestamp 1710899220
transform 1 0 72 0 1 1570
box -8 -3 16 105
use FILL  FILL_638
timestamp 1710899220
transform 1 0 2664 0 -1 1570
box -8 -3 16 105
use FILL  FILL_639
timestamp 1710899220
transform 1 0 2256 0 -1 1570
box -8 -3 16 105
use FILL  FILL_640
timestamp 1710899220
transform 1 0 2248 0 -1 1570
box -8 -3 16 105
use FILL  FILL_641
timestamp 1710899220
transform 1 0 2208 0 -1 1570
box -8 -3 16 105
use FILL  FILL_642
timestamp 1710899220
transform 1 0 2200 0 -1 1570
box -8 -3 16 105
use FILL  FILL_643
timestamp 1710899220
transform 1 0 1904 0 -1 1570
box -8 -3 16 105
use FILL  FILL_644
timestamp 1710899220
transform 1 0 1672 0 -1 1570
box -8 -3 16 105
use FILL  FILL_645
timestamp 1710899220
transform 1 0 1568 0 -1 1570
box -8 -3 16 105
use FILL  FILL_646
timestamp 1710899220
transform 1 0 1560 0 -1 1570
box -8 -3 16 105
use FILL  FILL_647
timestamp 1710899220
transform 1 0 1480 0 -1 1570
box -8 -3 16 105
use FILL  FILL_648
timestamp 1710899220
transform 1 0 1304 0 -1 1570
box -8 -3 16 105
use FILL  FILL_649
timestamp 1710899220
transform 1 0 736 0 -1 1570
box -8 -3 16 105
use FILL  FILL_650
timestamp 1710899220
transform 1 0 728 0 -1 1570
box -8 -3 16 105
use FILL  FILL_651
timestamp 1710899220
transform 1 0 648 0 -1 1570
box -8 -3 16 105
use FILL  FILL_652
timestamp 1710899220
transform 1 0 640 0 -1 1570
box -8 -3 16 105
use FILL  FILL_653
timestamp 1710899220
transform 1 0 560 0 -1 1570
box -8 -3 16 105
use FILL  FILL_654
timestamp 1710899220
transform 1 0 552 0 -1 1570
box -8 -3 16 105
use FILL  FILL_655
timestamp 1710899220
transform 1 0 504 0 -1 1570
box -8 -3 16 105
use FILL  FILL_656
timestamp 1710899220
transform 1 0 496 0 -1 1570
box -8 -3 16 105
use FILL  FILL_657
timestamp 1710899220
transform 1 0 488 0 -1 1570
box -8 -3 16 105
use FILL  FILL_658
timestamp 1710899220
transform 1 0 440 0 -1 1570
box -8 -3 16 105
use FILL  FILL_659
timestamp 1710899220
transform 1 0 432 0 -1 1570
box -8 -3 16 105
use FILL  FILL_660
timestamp 1710899220
transform 1 0 384 0 -1 1570
box -8 -3 16 105
use FILL  FILL_661
timestamp 1710899220
transform 1 0 376 0 -1 1570
box -8 -3 16 105
use FILL  FILL_662
timestamp 1710899220
transform 1 0 368 0 -1 1570
box -8 -3 16 105
use FILL  FILL_663
timestamp 1710899220
transform 1 0 320 0 -1 1570
box -8 -3 16 105
use FILL  FILL_664
timestamp 1710899220
transform 1 0 312 0 -1 1570
box -8 -3 16 105
use FILL  FILL_665
timestamp 1710899220
transform 1 0 272 0 -1 1570
box -8 -3 16 105
use FILL  FILL_666
timestamp 1710899220
transform 1 0 264 0 -1 1570
box -8 -3 16 105
use FILL  FILL_667
timestamp 1710899220
transform 1 0 256 0 -1 1570
box -8 -3 16 105
use FILL  FILL_668
timestamp 1710899220
transform 1 0 216 0 -1 1570
box -8 -3 16 105
use FILL  FILL_669
timestamp 1710899220
transform 1 0 208 0 -1 1570
box -8 -3 16 105
use FILL  FILL_670
timestamp 1710899220
transform 1 0 200 0 -1 1570
box -8 -3 16 105
use FILL  FILL_671
timestamp 1710899220
transform 1 0 136 0 -1 1570
box -8 -3 16 105
use FILL  FILL_672
timestamp 1710899220
transform 1 0 128 0 -1 1570
box -8 -3 16 105
use FILL  FILL_673
timestamp 1710899220
transform 1 0 120 0 -1 1570
box -8 -3 16 105
use FILL  FILL_674
timestamp 1710899220
transform 1 0 112 0 -1 1570
box -8 -3 16 105
use FILL  FILL_675
timestamp 1710899220
transform 1 0 104 0 -1 1570
box -8 -3 16 105
use FILL  FILL_676
timestamp 1710899220
transform 1 0 96 0 -1 1570
box -8 -3 16 105
use FILL  FILL_677
timestamp 1710899220
transform 1 0 88 0 -1 1570
box -8 -3 16 105
use FILL  FILL_678
timestamp 1710899220
transform 1 0 80 0 -1 1570
box -8 -3 16 105
use FILL  FILL_679
timestamp 1710899220
transform 1 0 72 0 -1 1570
box -8 -3 16 105
use FILL  FILL_680
timestamp 1710899220
transform 1 0 2664 0 1 1370
box -8 -3 16 105
use FILL  FILL_681
timestamp 1710899220
transform 1 0 2656 0 1 1370
box -8 -3 16 105
use FILL  FILL_682
timestamp 1710899220
transform 1 0 2648 0 1 1370
box -8 -3 16 105
use FILL  FILL_683
timestamp 1710899220
transform 1 0 2640 0 1 1370
box -8 -3 16 105
use FILL  FILL_684
timestamp 1710899220
transform 1 0 2520 0 1 1370
box -8 -3 16 105
use FILL  FILL_685
timestamp 1710899220
transform 1 0 2400 0 1 1370
box -8 -3 16 105
use FILL  FILL_686
timestamp 1710899220
transform 1 0 2392 0 1 1370
box -8 -3 16 105
use FILL  FILL_687
timestamp 1710899220
transform 1 0 2384 0 1 1370
box -8 -3 16 105
use FILL  FILL_688
timestamp 1710899220
transform 1 0 2376 0 1 1370
box -8 -3 16 105
use FILL  FILL_689
timestamp 1710899220
transform 1 0 2368 0 1 1370
box -8 -3 16 105
use FILL  FILL_690
timestamp 1710899220
transform 1 0 2264 0 1 1370
box -8 -3 16 105
use FILL  FILL_691
timestamp 1710899220
transform 1 0 2160 0 1 1370
box -8 -3 16 105
use FILL  FILL_692
timestamp 1710899220
transform 1 0 2152 0 1 1370
box -8 -3 16 105
use FILL  FILL_693
timestamp 1710899220
transform 1 0 2144 0 1 1370
box -8 -3 16 105
use FILL  FILL_694
timestamp 1710899220
transform 1 0 2136 0 1 1370
box -8 -3 16 105
use FILL  FILL_695
timestamp 1710899220
transform 1 0 2128 0 1 1370
box -8 -3 16 105
use FILL  FILL_696
timestamp 1710899220
transform 1 0 2096 0 1 1370
box -8 -3 16 105
use FILL  FILL_697
timestamp 1710899220
transform 1 0 2088 0 1 1370
box -8 -3 16 105
use FILL  FILL_698
timestamp 1710899220
transform 1 0 2080 0 1 1370
box -8 -3 16 105
use FILL  FILL_699
timestamp 1710899220
transform 1 0 2072 0 1 1370
box -8 -3 16 105
use FILL  FILL_700
timestamp 1710899220
transform 1 0 2064 0 1 1370
box -8 -3 16 105
use FILL  FILL_701
timestamp 1710899220
transform 1 0 2056 0 1 1370
box -8 -3 16 105
use FILL  FILL_702
timestamp 1710899220
transform 1 0 2048 0 1 1370
box -8 -3 16 105
use FILL  FILL_703
timestamp 1710899220
transform 1 0 1944 0 1 1370
box -8 -3 16 105
use FILL  FILL_704
timestamp 1710899220
transform 1 0 1936 0 1 1370
box -8 -3 16 105
use FILL  FILL_705
timestamp 1710899220
transform 1 0 1832 0 1 1370
box -8 -3 16 105
use FILL  FILL_706
timestamp 1710899220
transform 1 0 1824 0 1 1370
box -8 -3 16 105
use FILL  FILL_707
timestamp 1710899220
transform 1 0 1768 0 1 1370
box -8 -3 16 105
use FILL  FILL_708
timestamp 1710899220
transform 1 0 1736 0 1 1370
box -8 -3 16 105
use FILL  FILL_709
timestamp 1710899220
transform 1 0 1728 0 1 1370
box -8 -3 16 105
use FILL  FILL_710
timestamp 1710899220
transform 1 0 1624 0 1 1370
box -8 -3 16 105
use FILL  FILL_711
timestamp 1710899220
transform 1 0 1616 0 1 1370
box -8 -3 16 105
use FILL  FILL_712
timestamp 1710899220
transform 1 0 1536 0 1 1370
box -8 -3 16 105
use FILL  FILL_713
timestamp 1710899220
transform 1 0 1528 0 1 1370
box -8 -3 16 105
use FILL  FILL_714
timestamp 1710899220
transform 1 0 1424 0 1 1370
box -8 -3 16 105
use FILL  FILL_715
timestamp 1710899220
transform 1 0 1416 0 1 1370
box -8 -3 16 105
use FILL  FILL_716
timestamp 1710899220
transform 1 0 1408 0 1 1370
box -8 -3 16 105
use FILL  FILL_717
timestamp 1710899220
transform 1 0 1400 0 1 1370
box -8 -3 16 105
use FILL  FILL_718
timestamp 1710899220
transform 1 0 1392 0 1 1370
box -8 -3 16 105
use FILL  FILL_719
timestamp 1710899220
transform 1 0 1384 0 1 1370
box -8 -3 16 105
use FILL  FILL_720
timestamp 1710899220
transform 1 0 1376 0 1 1370
box -8 -3 16 105
use FILL  FILL_721
timestamp 1710899220
transform 1 0 1312 0 1 1370
box -8 -3 16 105
use FILL  FILL_722
timestamp 1710899220
transform 1 0 1208 0 1 1370
box -8 -3 16 105
use FILL  FILL_723
timestamp 1710899220
transform 1 0 1200 0 1 1370
box -8 -3 16 105
use FILL  FILL_724
timestamp 1710899220
transform 1 0 1192 0 1 1370
box -8 -3 16 105
use FILL  FILL_725
timestamp 1710899220
transform 1 0 1184 0 1 1370
box -8 -3 16 105
use FILL  FILL_726
timestamp 1710899220
transform 1 0 1120 0 1 1370
box -8 -3 16 105
use FILL  FILL_727
timestamp 1710899220
transform 1 0 1016 0 1 1370
box -8 -3 16 105
use FILL  FILL_728
timestamp 1710899220
transform 1 0 1008 0 1 1370
box -8 -3 16 105
use FILL  FILL_729
timestamp 1710899220
transform 1 0 1000 0 1 1370
box -8 -3 16 105
use FILL  FILL_730
timestamp 1710899220
transform 1 0 992 0 1 1370
box -8 -3 16 105
use FILL  FILL_731
timestamp 1710899220
transform 1 0 984 0 1 1370
box -8 -3 16 105
use FILL  FILL_732
timestamp 1710899220
transform 1 0 976 0 1 1370
box -8 -3 16 105
use FILL  FILL_733
timestamp 1710899220
transform 1 0 968 0 1 1370
box -8 -3 16 105
use FILL  FILL_734
timestamp 1710899220
transform 1 0 960 0 1 1370
box -8 -3 16 105
use FILL  FILL_735
timestamp 1710899220
transform 1 0 952 0 1 1370
box -8 -3 16 105
use FILL  FILL_736
timestamp 1710899220
transform 1 0 944 0 1 1370
box -8 -3 16 105
use FILL  FILL_737
timestamp 1710899220
transform 1 0 936 0 1 1370
box -8 -3 16 105
use FILL  FILL_738
timestamp 1710899220
transform 1 0 928 0 1 1370
box -8 -3 16 105
use FILL  FILL_739
timestamp 1710899220
transform 1 0 920 0 1 1370
box -8 -3 16 105
use FILL  FILL_740
timestamp 1710899220
transform 1 0 912 0 1 1370
box -8 -3 16 105
use FILL  FILL_741
timestamp 1710899220
transform 1 0 872 0 1 1370
box -8 -3 16 105
use FILL  FILL_742
timestamp 1710899220
transform 1 0 864 0 1 1370
box -8 -3 16 105
use FILL  FILL_743
timestamp 1710899220
transform 1 0 856 0 1 1370
box -8 -3 16 105
use FILL  FILL_744
timestamp 1710899220
transform 1 0 816 0 1 1370
box -8 -3 16 105
use FILL  FILL_745
timestamp 1710899220
transform 1 0 808 0 1 1370
box -8 -3 16 105
use FILL  FILL_746
timestamp 1710899220
transform 1 0 768 0 1 1370
box -8 -3 16 105
use FILL  FILL_747
timestamp 1710899220
transform 1 0 760 0 1 1370
box -8 -3 16 105
use FILL  FILL_748
timestamp 1710899220
transform 1 0 720 0 1 1370
box -8 -3 16 105
use FILL  FILL_749
timestamp 1710899220
transform 1 0 672 0 1 1370
box -8 -3 16 105
use FILL  FILL_750
timestamp 1710899220
transform 1 0 624 0 1 1370
box -8 -3 16 105
use FILL  FILL_751
timestamp 1710899220
transform 1 0 568 0 1 1370
box -8 -3 16 105
use FILL  FILL_752
timestamp 1710899220
transform 1 0 496 0 1 1370
box -8 -3 16 105
use FILL  FILL_753
timestamp 1710899220
transform 1 0 488 0 1 1370
box -8 -3 16 105
use FILL  FILL_754
timestamp 1710899220
transform 1 0 440 0 1 1370
box -8 -3 16 105
use FILL  FILL_755
timestamp 1710899220
transform 1 0 408 0 1 1370
box -8 -3 16 105
use FILL  FILL_756
timestamp 1710899220
transform 1 0 400 0 1 1370
box -8 -3 16 105
use FILL  FILL_757
timestamp 1710899220
transform 1 0 328 0 1 1370
box -8 -3 16 105
use FILL  FILL_758
timestamp 1710899220
transform 1 0 320 0 1 1370
box -8 -3 16 105
use FILL  FILL_759
timestamp 1710899220
transform 1 0 312 0 1 1370
box -8 -3 16 105
use FILL  FILL_760
timestamp 1710899220
transform 1 0 272 0 1 1370
box -8 -3 16 105
use FILL  FILL_761
timestamp 1710899220
transform 1 0 232 0 1 1370
box -8 -3 16 105
use FILL  FILL_762
timestamp 1710899220
transform 1 0 224 0 1 1370
box -8 -3 16 105
use FILL  FILL_763
timestamp 1710899220
transform 1 0 216 0 1 1370
box -8 -3 16 105
use FILL  FILL_764
timestamp 1710899220
transform 1 0 176 0 1 1370
box -8 -3 16 105
use FILL  FILL_765
timestamp 1710899220
transform 1 0 136 0 1 1370
box -8 -3 16 105
use FILL  FILL_766
timestamp 1710899220
transform 1 0 128 0 1 1370
box -8 -3 16 105
use FILL  FILL_767
timestamp 1710899220
transform 1 0 120 0 1 1370
box -8 -3 16 105
use FILL  FILL_768
timestamp 1710899220
transform 1 0 112 0 1 1370
box -8 -3 16 105
use FILL  FILL_769
timestamp 1710899220
transform 1 0 104 0 1 1370
box -8 -3 16 105
use FILL  FILL_770
timestamp 1710899220
transform 1 0 96 0 1 1370
box -8 -3 16 105
use FILL  FILL_771
timestamp 1710899220
transform 1 0 88 0 1 1370
box -8 -3 16 105
use FILL  FILL_772
timestamp 1710899220
transform 1 0 80 0 1 1370
box -8 -3 16 105
use FILL  FILL_773
timestamp 1710899220
transform 1 0 72 0 1 1370
box -8 -3 16 105
use FILL  FILL_774
timestamp 1710899220
transform 1 0 2568 0 -1 1370
box -8 -3 16 105
use FILL  FILL_775
timestamp 1710899220
transform 1 0 2560 0 -1 1370
box -8 -3 16 105
use FILL  FILL_776
timestamp 1710899220
transform 1 0 2496 0 -1 1370
box -8 -3 16 105
use FILL  FILL_777
timestamp 1710899220
transform 1 0 2488 0 -1 1370
box -8 -3 16 105
use FILL  FILL_778
timestamp 1710899220
transform 1 0 2480 0 -1 1370
box -8 -3 16 105
use FILL  FILL_779
timestamp 1710899220
transform 1 0 2472 0 -1 1370
box -8 -3 16 105
use FILL  FILL_780
timestamp 1710899220
transform 1 0 2464 0 -1 1370
box -8 -3 16 105
use FILL  FILL_781
timestamp 1710899220
transform 1 0 2456 0 -1 1370
box -8 -3 16 105
use FILL  FILL_782
timestamp 1710899220
transform 1 0 2448 0 -1 1370
box -8 -3 16 105
use FILL  FILL_783
timestamp 1710899220
transform 1 0 2360 0 -1 1370
box -8 -3 16 105
use FILL  FILL_784
timestamp 1710899220
transform 1 0 2352 0 -1 1370
box -8 -3 16 105
use FILL  FILL_785
timestamp 1710899220
transform 1 0 2288 0 -1 1370
box -8 -3 16 105
use FILL  FILL_786
timestamp 1710899220
transform 1 0 2280 0 -1 1370
box -8 -3 16 105
use FILL  FILL_787
timestamp 1710899220
transform 1 0 2240 0 -1 1370
box -8 -3 16 105
use FILL  FILL_788
timestamp 1710899220
transform 1 0 2232 0 -1 1370
box -8 -3 16 105
use FILL  FILL_789
timestamp 1710899220
transform 1 0 2168 0 -1 1370
box -8 -3 16 105
use FILL  FILL_790
timestamp 1710899220
transform 1 0 2160 0 -1 1370
box -8 -3 16 105
use FILL  FILL_791
timestamp 1710899220
transform 1 0 2152 0 -1 1370
box -8 -3 16 105
use FILL  FILL_792
timestamp 1710899220
transform 1 0 2112 0 -1 1370
box -8 -3 16 105
use FILL  FILL_793
timestamp 1710899220
transform 1 0 2104 0 -1 1370
box -8 -3 16 105
use FILL  FILL_794
timestamp 1710899220
transform 1 0 2096 0 -1 1370
box -8 -3 16 105
use FILL  FILL_795
timestamp 1710899220
transform 1 0 2088 0 -1 1370
box -8 -3 16 105
use FILL  FILL_796
timestamp 1710899220
transform 1 0 2080 0 -1 1370
box -8 -3 16 105
use FILL  FILL_797
timestamp 1710899220
transform 1 0 2072 0 -1 1370
box -8 -3 16 105
use FILL  FILL_798
timestamp 1710899220
transform 1 0 2032 0 -1 1370
box -8 -3 16 105
use FILL  FILL_799
timestamp 1710899220
transform 1 0 2000 0 -1 1370
box -8 -3 16 105
use FILL  FILL_800
timestamp 1710899220
transform 1 0 1992 0 -1 1370
box -8 -3 16 105
use FILL  FILL_801
timestamp 1710899220
transform 1 0 1984 0 -1 1370
box -8 -3 16 105
use FILL  FILL_802
timestamp 1710899220
transform 1 0 1976 0 -1 1370
box -8 -3 16 105
use FILL  FILL_803
timestamp 1710899220
transform 1 0 1968 0 -1 1370
box -8 -3 16 105
use FILL  FILL_804
timestamp 1710899220
transform 1 0 1960 0 -1 1370
box -8 -3 16 105
use FILL  FILL_805
timestamp 1710899220
transform 1 0 1904 0 -1 1370
box -8 -3 16 105
use FILL  FILL_806
timestamp 1710899220
transform 1 0 1896 0 -1 1370
box -8 -3 16 105
use FILL  FILL_807
timestamp 1710899220
transform 1 0 1888 0 -1 1370
box -8 -3 16 105
use FILL  FILL_808
timestamp 1710899220
transform 1 0 1880 0 -1 1370
box -8 -3 16 105
use FILL  FILL_809
timestamp 1710899220
transform 1 0 1872 0 -1 1370
box -8 -3 16 105
use FILL  FILL_810
timestamp 1710899220
transform 1 0 1864 0 -1 1370
box -8 -3 16 105
use FILL  FILL_811
timestamp 1710899220
transform 1 0 1856 0 -1 1370
box -8 -3 16 105
use FILL  FILL_812
timestamp 1710899220
transform 1 0 1848 0 -1 1370
box -8 -3 16 105
use FILL  FILL_813
timestamp 1710899220
transform 1 0 1792 0 -1 1370
box -8 -3 16 105
use FILL  FILL_814
timestamp 1710899220
transform 1 0 1784 0 -1 1370
box -8 -3 16 105
use FILL  FILL_815
timestamp 1710899220
transform 1 0 1472 0 -1 1370
box -8 -3 16 105
use FILL  FILL_816
timestamp 1710899220
transform 1 0 1464 0 -1 1370
box -8 -3 16 105
use FILL  FILL_817
timestamp 1710899220
transform 1 0 1248 0 -1 1370
box -8 -3 16 105
use FILL  FILL_818
timestamp 1710899220
transform 1 0 1184 0 -1 1370
box -8 -3 16 105
use FILL  FILL_819
timestamp 1710899220
transform 1 0 1104 0 -1 1370
box -8 -3 16 105
use FILL  FILL_820
timestamp 1710899220
transform 1 0 1080 0 -1 1370
box -8 -3 16 105
use FILL  FILL_821
timestamp 1710899220
transform 1 0 1072 0 -1 1370
box -8 -3 16 105
use FILL  FILL_822
timestamp 1710899220
transform 1 0 1024 0 -1 1370
box -8 -3 16 105
use FILL  FILL_823
timestamp 1710899220
transform 1 0 992 0 -1 1370
box -8 -3 16 105
use FILL  FILL_824
timestamp 1710899220
transform 1 0 920 0 -1 1370
box -8 -3 16 105
use FILL  FILL_825
timestamp 1710899220
transform 1 0 832 0 -1 1370
box -8 -3 16 105
use FILL  FILL_826
timestamp 1710899220
transform 1 0 744 0 -1 1370
box -8 -3 16 105
use FILL  FILL_827
timestamp 1710899220
transform 1 0 736 0 -1 1370
box -8 -3 16 105
use FILL  FILL_828
timestamp 1710899220
transform 1 0 648 0 -1 1370
box -8 -3 16 105
use FILL  FILL_829
timestamp 1710899220
transform 1 0 568 0 -1 1370
box -8 -3 16 105
use FILL  FILL_830
timestamp 1710899220
transform 1 0 504 0 -1 1370
box -8 -3 16 105
use FILL  FILL_831
timestamp 1710899220
transform 1 0 496 0 -1 1370
box -8 -3 16 105
use FILL  FILL_832
timestamp 1710899220
transform 1 0 488 0 -1 1370
box -8 -3 16 105
use FILL  FILL_833
timestamp 1710899220
transform 1 0 416 0 -1 1370
box -8 -3 16 105
use FILL  FILL_834
timestamp 1710899220
transform 1 0 408 0 -1 1370
box -8 -3 16 105
use FILL  FILL_835
timestamp 1710899220
transform 1 0 400 0 -1 1370
box -8 -3 16 105
use FILL  FILL_836
timestamp 1710899220
transform 1 0 304 0 -1 1370
box -8 -3 16 105
use FILL  FILL_837
timestamp 1710899220
transform 1 0 1768 0 1 1170
box -8 -3 16 105
use FILL  FILL_838
timestamp 1710899220
transform 1 0 1704 0 1 1170
box -8 -3 16 105
use FILL  FILL_839
timestamp 1710899220
transform 1 0 1696 0 1 1170
box -8 -3 16 105
use FILL  FILL_840
timestamp 1710899220
transform 1 0 1688 0 1 1170
box -8 -3 16 105
use FILL  FILL_841
timestamp 1710899220
transform 1 0 1680 0 1 1170
box -8 -3 16 105
use FILL  FILL_842
timestamp 1710899220
transform 1 0 1656 0 1 1170
box -8 -3 16 105
use FILL  FILL_843
timestamp 1710899220
transform 1 0 1648 0 1 1170
box -8 -3 16 105
use FILL  FILL_844
timestamp 1710899220
transform 1 0 1512 0 1 1170
box -8 -3 16 105
use FILL  FILL_845
timestamp 1710899220
transform 1 0 1352 0 1 1170
box -8 -3 16 105
use FILL  FILL_846
timestamp 1710899220
transform 1 0 1248 0 1 1170
box -8 -3 16 105
use FILL  FILL_847
timestamp 1710899220
transform 1 0 1008 0 1 1170
box -8 -3 16 105
use FILL  FILL_848
timestamp 1710899220
transform 1 0 928 0 1 1170
box -8 -3 16 105
use FILL  FILL_849
timestamp 1710899220
transform 1 0 848 0 1 1170
box -8 -3 16 105
use FILL  FILL_850
timestamp 1710899220
transform 1 0 776 0 1 1170
box -8 -3 16 105
use FILL  FILL_851
timestamp 1710899220
transform 1 0 664 0 1 1170
box -8 -3 16 105
use FILL  FILL_852
timestamp 1710899220
transform 1 0 656 0 1 1170
box -8 -3 16 105
use FILL  FILL_853
timestamp 1710899220
transform 1 0 576 0 1 1170
box -8 -3 16 105
use FILL  FILL_854
timestamp 1710899220
transform 1 0 568 0 1 1170
box -8 -3 16 105
use FILL  FILL_855
timestamp 1710899220
transform 1 0 488 0 1 1170
box -8 -3 16 105
use FILL  FILL_856
timestamp 1710899220
transform 1 0 400 0 1 1170
box -8 -3 16 105
use FILL  FILL_857
timestamp 1710899220
transform 1 0 328 0 1 1170
box -8 -3 16 105
use FILL  FILL_858
timestamp 1710899220
transform 1 0 320 0 1 1170
box -8 -3 16 105
use FILL  FILL_859
timestamp 1710899220
transform 1 0 248 0 1 1170
box -8 -3 16 105
use FILL  FILL_860
timestamp 1710899220
transform 1 0 240 0 1 1170
box -8 -3 16 105
use FILL  FILL_861
timestamp 1710899220
transform 1 0 168 0 1 1170
box -8 -3 16 105
use FILL  FILL_862
timestamp 1710899220
transform 1 0 160 0 1 1170
box -8 -3 16 105
use FILL  FILL_863
timestamp 1710899220
transform 1 0 152 0 1 1170
box -8 -3 16 105
use FILL  FILL_864
timestamp 1710899220
transform 1 0 144 0 1 1170
box -8 -3 16 105
use FILL  FILL_865
timestamp 1710899220
transform 1 0 80 0 1 1170
box -8 -3 16 105
use FILL  FILL_866
timestamp 1710899220
transform 1 0 72 0 1 1170
box -8 -3 16 105
use FILL  FILL_867
timestamp 1710899220
transform 1 0 2440 0 -1 1170
box -8 -3 16 105
use FILL  FILL_868
timestamp 1710899220
transform 1 0 2432 0 -1 1170
box -8 -3 16 105
use FILL  FILL_869
timestamp 1710899220
transform 1 0 2424 0 -1 1170
box -8 -3 16 105
use FILL  FILL_870
timestamp 1710899220
transform 1 0 2320 0 -1 1170
box -8 -3 16 105
use FILL  FILL_871
timestamp 1710899220
transform 1 0 2312 0 -1 1170
box -8 -3 16 105
use FILL  FILL_872
timestamp 1710899220
transform 1 0 2304 0 -1 1170
box -8 -3 16 105
use FILL  FILL_873
timestamp 1710899220
transform 1 0 2240 0 -1 1170
box -8 -3 16 105
use FILL  FILL_874
timestamp 1710899220
transform 1 0 2136 0 -1 1170
box -8 -3 16 105
use FILL  FILL_875
timestamp 1710899220
transform 1 0 2128 0 -1 1170
box -8 -3 16 105
use FILL  FILL_876
timestamp 1710899220
transform 1 0 2120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_877
timestamp 1710899220
transform 1 0 2112 0 -1 1170
box -8 -3 16 105
use FILL  FILL_878
timestamp 1710899220
transform 1 0 2104 0 -1 1170
box -8 -3 16 105
use FILL  FILL_879
timestamp 1710899220
transform 1 0 2096 0 -1 1170
box -8 -3 16 105
use FILL  FILL_880
timestamp 1710899220
transform 1 0 2088 0 -1 1170
box -8 -3 16 105
use FILL  FILL_881
timestamp 1710899220
transform 1 0 2080 0 -1 1170
box -8 -3 16 105
use FILL  FILL_882
timestamp 1710899220
transform 1 0 2072 0 -1 1170
box -8 -3 16 105
use FILL  FILL_883
timestamp 1710899220
transform 1 0 2064 0 -1 1170
box -8 -3 16 105
use FILL  FILL_884
timestamp 1710899220
transform 1 0 2032 0 -1 1170
box -8 -3 16 105
use FILL  FILL_885
timestamp 1710899220
transform 1 0 2024 0 -1 1170
box -8 -3 16 105
use FILL  FILL_886
timestamp 1710899220
transform 1 0 2016 0 -1 1170
box -8 -3 16 105
use FILL  FILL_887
timestamp 1710899220
transform 1 0 2008 0 -1 1170
box -8 -3 16 105
use FILL  FILL_888
timestamp 1710899220
transform 1 0 2000 0 -1 1170
box -8 -3 16 105
use FILL  FILL_889
timestamp 1710899220
transform 1 0 1992 0 -1 1170
box -8 -3 16 105
use FILL  FILL_890
timestamp 1710899220
transform 1 0 1984 0 -1 1170
box -8 -3 16 105
use FILL  FILL_891
timestamp 1710899220
transform 1 0 1976 0 -1 1170
box -8 -3 16 105
use FILL  FILL_892
timestamp 1710899220
transform 1 0 1872 0 -1 1170
box -8 -3 16 105
use FILL  FILL_893
timestamp 1710899220
transform 1 0 1864 0 -1 1170
box -8 -3 16 105
use FILL  FILL_894
timestamp 1710899220
transform 1 0 1856 0 -1 1170
box -8 -3 16 105
use FILL  FILL_895
timestamp 1710899220
transform 1 0 1792 0 -1 1170
box -8 -3 16 105
use FILL  FILL_896
timestamp 1710899220
transform 1 0 1784 0 -1 1170
box -8 -3 16 105
use FILL  FILL_897
timestamp 1710899220
transform 1 0 1776 0 -1 1170
box -8 -3 16 105
use FILL  FILL_898
timestamp 1710899220
transform 1 0 1744 0 -1 1170
box -8 -3 16 105
use FILL  FILL_899
timestamp 1710899220
transform 1 0 1720 0 -1 1170
box -8 -3 16 105
use FILL  FILL_900
timestamp 1710899220
transform 1 0 1712 0 -1 1170
box -8 -3 16 105
use FILL  FILL_901
timestamp 1710899220
transform 1 0 1616 0 -1 1170
box -8 -3 16 105
use FILL  FILL_902
timestamp 1710899220
transform 1 0 1608 0 -1 1170
box -8 -3 16 105
use FILL  FILL_903
timestamp 1710899220
transform 1 0 1600 0 -1 1170
box -8 -3 16 105
use FILL  FILL_904
timestamp 1710899220
transform 1 0 1456 0 -1 1170
box -8 -3 16 105
use FILL  FILL_905
timestamp 1710899220
transform 1 0 1296 0 -1 1170
box -8 -3 16 105
use FILL  FILL_906
timestamp 1710899220
transform 1 0 1192 0 -1 1170
box -8 -3 16 105
use FILL  FILL_907
timestamp 1710899220
transform 1 0 1088 0 -1 1170
box -8 -3 16 105
use FILL  FILL_908
timestamp 1710899220
transform 1 0 1080 0 -1 1170
box -8 -3 16 105
use FILL  FILL_909
timestamp 1710899220
transform 1 0 1072 0 -1 1170
box -8 -3 16 105
use FILL  FILL_910
timestamp 1710899220
transform 1 0 1064 0 -1 1170
box -8 -3 16 105
use FILL  FILL_911
timestamp 1710899220
transform 1 0 1056 0 -1 1170
box -8 -3 16 105
use FILL  FILL_912
timestamp 1710899220
transform 1 0 1008 0 -1 1170
box -8 -3 16 105
use FILL  FILL_913
timestamp 1710899220
transform 1 0 1000 0 -1 1170
box -8 -3 16 105
use FILL  FILL_914
timestamp 1710899220
transform 1 0 944 0 -1 1170
box -8 -3 16 105
use FILL  FILL_915
timestamp 1710899220
transform 1 0 936 0 -1 1170
box -8 -3 16 105
use FILL  FILL_916
timestamp 1710899220
transform 1 0 928 0 -1 1170
box -8 -3 16 105
use FILL  FILL_917
timestamp 1710899220
transform 1 0 896 0 -1 1170
box -8 -3 16 105
use FILL  FILL_918
timestamp 1710899220
transform 1 0 888 0 -1 1170
box -8 -3 16 105
use FILL  FILL_919
timestamp 1710899220
transform 1 0 840 0 -1 1170
box -8 -3 16 105
use FILL  FILL_920
timestamp 1710899220
transform 1 0 832 0 -1 1170
box -8 -3 16 105
use FILL  FILL_921
timestamp 1710899220
transform 1 0 824 0 -1 1170
box -8 -3 16 105
use FILL  FILL_922
timestamp 1710899220
transform 1 0 792 0 -1 1170
box -8 -3 16 105
use FILL  FILL_923
timestamp 1710899220
transform 1 0 784 0 -1 1170
box -8 -3 16 105
use FILL  FILL_924
timestamp 1710899220
transform 1 0 776 0 -1 1170
box -8 -3 16 105
use FILL  FILL_925
timestamp 1710899220
transform 1 0 768 0 -1 1170
box -8 -3 16 105
use FILL  FILL_926
timestamp 1710899220
transform 1 0 728 0 -1 1170
box -8 -3 16 105
use FILL  FILL_927
timestamp 1710899220
transform 1 0 720 0 -1 1170
box -8 -3 16 105
use FILL  FILL_928
timestamp 1710899220
transform 1 0 672 0 -1 1170
box -8 -3 16 105
use FILL  FILL_929
timestamp 1710899220
transform 1 0 664 0 -1 1170
box -8 -3 16 105
use FILL  FILL_930
timestamp 1710899220
transform 1 0 656 0 -1 1170
box -8 -3 16 105
use FILL  FILL_931
timestamp 1710899220
transform 1 0 648 0 -1 1170
box -8 -3 16 105
use FILL  FILL_932
timestamp 1710899220
transform 1 0 640 0 -1 1170
box -8 -3 16 105
use FILL  FILL_933
timestamp 1710899220
transform 1 0 592 0 -1 1170
box -8 -3 16 105
use FILL  FILL_934
timestamp 1710899220
transform 1 0 584 0 -1 1170
box -8 -3 16 105
use FILL  FILL_935
timestamp 1710899220
transform 1 0 536 0 -1 1170
box -8 -3 16 105
use FILL  FILL_936
timestamp 1710899220
transform 1 0 528 0 -1 1170
box -8 -3 16 105
use FILL  FILL_937
timestamp 1710899220
transform 1 0 520 0 -1 1170
box -8 -3 16 105
use FILL  FILL_938
timestamp 1710899220
transform 1 0 512 0 -1 1170
box -8 -3 16 105
use FILL  FILL_939
timestamp 1710899220
transform 1 0 464 0 -1 1170
box -8 -3 16 105
use FILL  FILL_940
timestamp 1710899220
transform 1 0 456 0 -1 1170
box -8 -3 16 105
use FILL  FILL_941
timestamp 1710899220
transform 1 0 448 0 -1 1170
box -8 -3 16 105
use FILL  FILL_942
timestamp 1710899220
transform 1 0 440 0 -1 1170
box -8 -3 16 105
use FILL  FILL_943
timestamp 1710899220
transform 1 0 432 0 -1 1170
box -8 -3 16 105
use FILL  FILL_944
timestamp 1710899220
transform 1 0 384 0 -1 1170
box -8 -3 16 105
use FILL  FILL_945
timestamp 1710899220
transform 1 0 376 0 -1 1170
box -8 -3 16 105
use FILL  FILL_946
timestamp 1710899220
transform 1 0 328 0 -1 1170
box -8 -3 16 105
use FILL  FILL_947
timestamp 1710899220
transform 1 0 320 0 -1 1170
box -8 -3 16 105
use FILL  FILL_948
timestamp 1710899220
transform 1 0 312 0 -1 1170
box -8 -3 16 105
use FILL  FILL_949
timestamp 1710899220
transform 1 0 304 0 -1 1170
box -8 -3 16 105
use FILL  FILL_950
timestamp 1710899220
transform 1 0 296 0 -1 1170
box -8 -3 16 105
use FILL  FILL_951
timestamp 1710899220
transform 1 0 288 0 -1 1170
box -8 -3 16 105
use FILL  FILL_952
timestamp 1710899220
transform 1 0 280 0 -1 1170
box -8 -3 16 105
use FILL  FILL_953
timestamp 1710899220
transform 1 0 216 0 -1 1170
box -8 -3 16 105
use FILL  FILL_954
timestamp 1710899220
transform 1 0 208 0 -1 1170
box -8 -3 16 105
use FILL  FILL_955
timestamp 1710899220
transform 1 0 200 0 -1 1170
box -8 -3 16 105
use FILL  FILL_956
timestamp 1710899220
transform 1 0 192 0 -1 1170
box -8 -3 16 105
use FILL  FILL_957
timestamp 1710899220
transform 1 0 96 0 -1 1170
box -8 -3 16 105
use FILL  FILL_958
timestamp 1710899220
transform 1 0 88 0 -1 1170
box -8 -3 16 105
use FILL  FILL_959
timestamp 1710899220
transform 1 0 80 0 -1 1170
box -8 -3 16 105
use FILL  FILL_960
timestamp 1710899220
transform 1 0 72 0 -1 1170
box -8 -3 16 105
use FILL  FILL_961
timestamp 1710899220
transform 1 0 2664 0 1 970
box -8 -3 16 105
use FILL  FILL_962
timestamp 1710899220
transform 1 0 2656 0 1 970
box -8 -3 16 105
use FILL  FILL_963
timestamp 1710899220
transform 1 0 2648 0 1 970
box -8 -3 16 105
use FILL  FILL_964
timestamp 1710899220
transform 1 0 2640 0 1 970
box -8 -3 16 105
use FILL  FILL_965
timestamp 1710899220
transform 1 0 2632 0 1 970
box -8 -3 16 105
use FILL  FILL_966
timestamp 1710899220
transform 1 0 2624 0 1 970
box -8 -3 16 105
use FILL  FILL_967
timestamp 1710899220
transform 1 0 2592 0 1 970
box -8 -3 16 105
use FILL  FILL_968
timestamp 1710899220
transform 1 0 2584 0 1 970
box -8 -3 16 105
use FILL  FILL_969
timestamp 1710899220
transform 1 0 2544 0 1 970
box -8 -3 16 105
use FILL  FILL_970
timestamp 1710899220
transform 1 0 2536 0 1 970
box -8 -3 16 105
use FILL  FILL_971
timestamp 1710899220
transform 1 0 2528 0 1 970
box -8 -3 16 105
use FILL  FILL_972
timestamp 1710899220
transform 1 0 2520 0 1 970
box -8 -3 16 105
use FILL  FILL_973
timestamp 1710899220
transform 1 0 2512 0 1 970
box -8 -3 16 105
use FILL  FILL_974
timestamp 1710899220
transform 1 0 2504 0 1 970
box -8 -3 16 105
use FILL  FILL_975
timestamp 1710899220
transform 1 0 2432 0 1 970
box -8 -3 16 105
use FILL  FILL_976
timestamp 1710899220
transform 1 0 2424 0 1 970
box -8 -3 16 105
use FILL  FILL_977
timestamp 1710899220
transform 1 0 2416 0 1 970
box -8 -3 16 105
use FILL  FILL_978
timestamp 1710899220
transform 1 0 2408 0 1 970
box -8 -3 16 105
use FILL  FILL_979
timestamp 1710899220
transform 1 0 2400 0 1 970
box -8 -3 16 105
use FILL  FILL_980
timestamp 1710899220
transform 1 0 2392 0 1 970
box -8 -3 16 105
use FILL  FILL_981
timestamp 1710899220
transform 1 0 2384 0 1 970
box -8 -3 16 105
use FILL  FILL_982
timestamp 1710899220
transform 1 0 2376 0 1 970
box -8 -3 16 105
use FILL  FILL_983
timestamp 1710899220
transform 1 0 2368 0 1 970
box -8 -3 16 105
use FILL  FILL_984
timestamp 1710899220
transform 1 0 2360 0 1 970
box -8 -3 16 105
use FILL  FILL_985
timestamp 1710899220
transform 1 0 2352 0 1 970
box -8 -3 16 105
use FILL  FILL_986
timestamp 1710899220
transform 1 0 2344 0 1 970
box -8 -3 16 105
use FILL  FILL_987
timestamp 1710899220
transform 1 0 2336 0 1 970
box -8 -3 16 105
use FILL  FILL_988
timestamp 1710899220
transform 1 0 2328 0 1 970
box -8 -3 16 105
use FILL  FILL_989
timestamp 1710899220
transform 1 0 2296 0 1 970
box -8 -3 16 105
use FILL  FILL_990
timestamp 1710899220
transform 1 0 1944 0 1 970
box -8 -3 16 105
use FILL  FILL_991
timestamp 1710899220
transform 1 0 1880 0 1 970
box -8 -3 16 105
use FILL  FILL_992
timestamp 1710899220
transform 1 0 1872 0 1 970
box -8 -3 16 105
use FILL  FILL_993
timestamp 1710899220
transform 1 0 1776 0 1 970
box -8 -3 16 105
use FILL  FILL_994
timestamp 1710899220
transform 1 0 1656 0 1 970
box -8 -3 16 105
use FILL  FILL_995
timestamp 1710899220
transform 1 0 1472 0 1 970
box -8 -3 16 105
use FILL  FILL_996
timestamp 1710899220
transform 1 0 1464 0 1 970
box -8 -3 16 105
use FILL  FILL_997
timestamp 1710899220
transform 1 0 1400 0 1 970
box -8 -3 16 105
use FILL  FILL_998
timestamp 1710899220
transform 1 0 1392 0 1 970
box -8 -3 16 105
use FILL  FILL_999
timestamp 1710899220
transform 1 0 1384 0 1 970
box -8 -3 16 105
use FILL  FILL_1000
timestamp 1710899220
transform 1 0 1376 0 1 970
box -8 -3 16 105
use FILL  FILL_1001
timestamp 1710899220
transform 1 0 1312 0 1 970
box -8 -3 16 105
use FILL  FILL_1002
timestamp 1710899220
transform 1 0 1208 0 1 970
box -8 -3 16 105
use FILL  FILL_1003
timestamp 1710899220
transform 1 0 1200 0 1 970
box -8 -3 16 105
use FILL  FILL_1004
timestamp 1710899220
transform 1 0 1136 0 1 970
box -8 -3 16 105
use FILL  FILL_1005
timestamp 1710899220
transform 1 0 1032 0 1 970
box -8 -3 16 105
use FILL  FILL_1006
timestamp 1710899220
transform 1 0 776 0 1 970
box -8 -3 16 105
use FILL  FILL_1007
timestamp 1710899220
transform 1 0 768 0 1 970
box -8 -3 16 105
use FILL  FILL_1008
timestamp 1710899220
transform 1 0 688 0 1 970
box -8 -3 16 105
use FILL  FILL_1009
timestamp 1710899220
transform 1 0 664 0 1 970
box -8 -3 16 105
use FILL  FILL_1010
timestamp 1710899220
transform 1 0 608 0 1 970
box -8 -3 16 105
use FILL  FILL_1011
timestamp 1710899220
transform 1 0 600 0 1 970
box -8 -3 16 105
use FILL  FILL_1012
timestamp 1710899220
transform 1 0 544 0 1 970
box -8 -3 16 105
use FILL  FILL_1013
timestamp 1710899220
transform 1 0 536 0 1 970
box -8 -3 16 105
use FILL  FILL_1014
timestamp 1710899220
transform 1 0 528 0 1 970
box -8 -3 16 105
use FILL  FILL_1015
timestamp 1710899220
transform 1 0 448 0 1 970
box -8 -3 16 105
use FILL  FILL_1016
timestamp 1710899220
transform 1 0 400 0 1 970
box -8 -3 16 105
use FILL  FILL_1017
timestamp 1710899220
transform 1 0 392 0 1 970
box -8 -3 16 105
use FILL  FILL_1018
timestamp 1710899220
transform 1 0 344 0 1 970
box -8 -3 16 105
use FILL  FILL_1019
timestamp 1710899220
transform 1 0 336 0 1 970
box -8 -3 16 105
use FILL  FILL_1020
timestamp 1710899220
transform 1 0 328 0 1 970
box -8 -3 16 105
use FILL  FILL_1021
timestamp 1710899220
transform 1 0 264 0 1 970
box -8 -3 16 105
use FILL  FILL_1022
timestamp 1710899220
transform 1 0 256 0 1 970
box -8 -3 16 105
use FILL  FILL_1023
timestamp 1710899220
transform 1 0 248 0 1 970
box -8 -3 16 105
use FILL  FILL_1024
timestamp 1710899220
transform 1 0 240 0 1 970
box -8 -3 16 105
use FILL  FILL_1025
timestamp 1710899220
transform 1 0 232 0 1 970
box -8 -3 16 105
use FILL  FILL_1026
timestamp 1710899220
transform 1 0 160 0 1 970
box -8 -3 16 105
use FILL  FILL_1027
timestamp 1710899220
transform 1 0 152 0 1 970
box -8 -3 16 105
use FILL  FILL_1028
timestamp 1710899220
transform 1 0 144 0 1 970
box -8 -3 16 105
use FILL  FILL_1029
timestamp 1710899220
transform 1 0 80 0 1 970
box -8 -3 16 105
use FILL  FILL_1030
timestamp 1710899220
transform 1 0 72 0 1 970
box -8 -3 16 105
use FILL  FILL_1031
timestamp 1710899220
transform 1 0 2664 0 -1 970
box -8 -3 16 105
use FILL  FILL_1032
timestamp 1710899220
transform 1 0 2656 0 -1 970
box -8 -3 16 105
use FILL  FILL_1033
timestamp 1710899220
transform 1 0 2648 0 -1 970
box -8 -3 16 105
use FILL  FILL_1034
timestamp 1710899220
transform 1 0 2640 0 -1 970
box -8 -3 16 105
use FILL  FILL_1035
timestamp 1710899220
transform 1 0 2536 0 -1 970
box -8 -3 16 105
use FILL  FILL_1036
timestamp 1710899220
transform 1 0 2456 0 -1 970
box -8 -3 16 105
use FILL  FILL_1037
timestamp 1710899220
transform 1 0 2448 0 -1 970
box -8 -3 16 105
use FILL  FILL_1038
timestamp 1710899220
transform 1 0 2440 0 -1 970
box -8 -3 16 105
use FILL  FILL_1039
timestamp 1710899220
transform 1 0 2360 0 -1 970
box -8 -3 16 105
use FILL  FILL_1040
timestamp 1710899220
transform 1 0 2320 0 -1 970
box -8 -3 16 105
use FILL  FILL_1041
timestamp 1710899220
transform 1 0 2240 0 -1 970
box -8 -3 16 105
use FILL  FILL_1042
timestamp 1710899220
transform 1 0 2232 0 -1 970
box -8 -3 16 105
use FILL  FILL_1043
timestamp 1710899220
transform 1 0 2224 0 -1 970
box -8 -3 16 105
use FILL  FILL_1044
timestamp 1710899220
transform 1 0 2216 0 -1 970
box -8 -3 16 105
use FILL  FILL_1045
timestamp 1710899220
transform 1 0 2208 0 -1 970
box -8 -3 16 105
use FILL  FILL_1046
timestamp 1710899220
transform 1 0 2200 0 -1 970
box -8 -3 16 105
use FILL  FILL_1047
timestamp 1710899220
transform 1 0 2192 0 -1 970
box -8 -3 16 105
use FILL  FILL_1048
timestamp 1710899220
transform 1 0 2184 0 -1 970
box -8 -3 16 105
use FILL  FILL_1049
timestamp 1710899220
transform 1 0 2176 0 -1 970
box -8 -3 16 105
use FILL  FILL_1050
timestamp 1710899220
transform 1 0 2664 0 1 770
box -8 -3 16 105
use FILL  FILL_1051
timestamp 1710899220
transform 1 0 2576 0 1 770
box -8 -3 16 105
use FILL  FILL_1052
timestamp 1710899220
transform 1 0 2568 0 1 770
box -8 -3 16 105
use FILL  FILL_1053
timestamp 1710899220
transform 1 0 2496 0 1 770
box -8 -3 16 105
use FILL  FILL_1054
timestamp 1710899220
transform 1 0 2488 0 1 770
box -8 -3 16 105
use FILL  FILL_1055
timestamp 1710899220
transform 1 0 2400 0 1 770
box -8 -3 16 105
use FILL  FILL_1056
timestamp 1710899220
transform 1 0 2392 0 1 770
box -8 -3 16 105
use FILL  FILL_1057
timestamp 1710899220
transform 1 0 2384 0 1 770
box -8 -3 16 105
use FILL  FILL_1058
timestamp 1710899220
transform 1 0 2312 0 1 770
box -8 -3 16 105
use FILL  FILL_1059
timestamp 1710899220
transform 1 0 2304 0 1 770
box -8 -3 16 105
use FILL  FILL_1060
timestamp 1710899220
transform 1 0 2296 0 1 770
box -8 -3 16 105
use FILL  FILL_1061
timestamp 1710899220
transform 1 0 2256 0 1 770
box -8 -3 16 105
use FILL  FILL_1062
timestamp 1710899220
transform 1 0 2248 0 1 770
box -8 -3 16 105
use FILL  FILL_1063
timestamp 1710899220
transform 1 0 2240 0 1 770
box -8 -3 16 105
use FILL  FILL_1064
timestamp 1710899220
transform 1 0 2232 0 1 770
box -8 -3 16 105
use FILL  FILL_1065
timestamp 1710899220
transform 1 0 2224 0 1 770
box -8 -3 16 105
use FILL  FILL_1066
timestamp 1710899220
transform 1 0 2216 0 1 770
box -8 -3 16 105
use FILL  FILL_1067
timestamp 1710899220
transform 1 0 2152 0 1 770
box -8 -3 16 105
use FILL  FILL_1068
timestamp 1710899220
transform 1 0 2144 0 1 770
box -8 -3 16 105
use FILL  FILL_1069
timestamp 1710899220
transform 1 0 2024 0 1 770
box -8 -3 16 105
use FILL  FILL_1070
timestamp 1710899220
transform 1 0 2016 0 1 770
box -8 -3 16 105
use FILL  FILL_1071
timestamp 1710899220
transform 1 0 1952 0 1 770
box -8 -3 16 105
use FILL  FILL_1072
timestamp 1710899220
transform 1 0 1840 0 1 770
box -8 -3 16 105
use FILL  FILL_1073
timestamp 1710899220
transform 1 0 1760 0 1 770
box -8 -3 16 105
use FILL  FILL_1074
timestamp 1710899220
transform 1 0 1752 0 1 770
box -8 -3 16 105
use FILL  FILL_1075
timestamp 1710899220
transform 1 0 1360 0 1 770
box -8 -3 16 105
use FILL  FILL_1076
timestamp 1710899220
transform 1 0 1352 0 1 770
box -8 -3 16 105
use FILL  FILL_1077
timestamp 1710899220
transform 1 0 1248 0 1 770
box -8 -3 16 105
use FILL  FILL_1078
timestamp 1710899220
transform 1 0 1160 0 1 770
box -8 -3 16 105
use FILL  FILL_1079
timestamp 1710899220
transform 1 0 1152 0 1 770
box -8 -3 16 105
use FILL  FILL_1080
timestamp 1710899220
transform 1 0 1064 0 1 770
box -8 -3 16 105
use FILL  FILL_1081
timestamp 1710899220
transform 1 0 944 0 1 770
box -8 -3 16 105
use FILL  FILL_1082
timestamp 1710899220
transform 1 0 864 0 1 770
box -8 -3 16 105
use FILL  FILL_1083
timestamp 1710899220
transform 1 0 856 0 1 770
box -8 -3 16 105
use FILL  FILL_1084
timestamp 1710899220
transform 1 0 832 0 1 770
box -8 -3 16 105
use FILL  FILL_1085
timestamp 1710899220
transform 1 0 760 0 1 770
box -8 -3 16 105
use FILL  FILL_1086
timestamp 1710899220
transform 1 0 656 0 1 770
box -8 -3 16 105
use FILL  FILL_1087
timestamp 1710899220
transform 1 0 648 0 1 770
box -8 -3 16 105
use FILL  FILL_1088
timestamp 1710899220
transform 1 0 576 0 1 770
box -8 -3 16 105
use FILL  FILL_1089
timestamp 1710899220
transform 1 0 568 0 1 770
box -8 -3 16 105
use FILL  FILL_1090
timestamp 1710899220
transform 1 0 488 0 1 770
box -8 -3 16 105
use FILL  FILL_1091
timestamp 1710899220
transform 1 0 480 0 1 770
box -8 -3 16 105
use FILL  FILL_1092
timestamp 1710899220
transform 1 0 312 0 1 770
box -8 -3 16 105
use FILL  FILL_1093
timestamp 1710899220
transform 1 0 224 0 1 770
box -8 -3 16 105
use FILL  FILL_1094
timestamp 1710899220
transform 1 0 192 0 1 770
box -8 -3 16 105
use FILL  FILL_1095
timestamp 1710899220
transform 1 0 128 0 1 770
box -8 -3 16 105
use FILL  FILL_1096
timestamp 1710899220
transform 1 0 88 0 1 770
box -8 -3 16 105
use FILL  FILL_1097
timestamp 1710899220
transform 1 0 80 0 1 770
box -8 -3 16 105
use FILL  FILL_1098
timestamp 1710899220
transform 1 0 72 0 1 770
box -8 -3 16 105
use FILL  FILL_1099
timestamp 1710899220
transform 1 0 2664 0 -1 770
box -8 -3 16 105
use FILL  FILL_1100
timestamp 1710899220
transform 1 0 2656 0 -1 770
box -8 -3 16 105
use FILL  FILL_1101
timestamp 1710899220
transform 1 0 2648 0 -1 770
box -8 -3 16 105
use FILL  FILL_1102
timestamp 1710899220
transform 1 0 2640 0 -1 770
box -8 -3 16 105
use FILL  FILL_1103
timestamp 1710899220
transform 1 0 2584 0 -1 770
box -8 -3 16 105
use FILL  FILL_1104
timestamp 1710899220
transform 1 0 2552 0 -1 770
box -8 -3 16 105
use FILL  FILL_1105
timestamp 1710899220
transform 1 0 2512 0 -1 770
box -8 -3 16 105
use FILL  FILL_1106
timestamp 1710899220
transform 1 0 2504 0 -1 770
box -8 -3 16 105
use FILL  FILL_1107
timestamp 1710899220
transform 1 0 2496 0 -1 770
box -8 -3 16 105
use FILL  FILL_1108
timestamp 1710899220
transform 1 0 2440 0 -1 770
box -8 -3 16 105
use FILL  FILL_1109
timestamp 1710899220
transform 1 0 2432 0 -1 770
box -8 -3 16 105
use FILL  FILL_1110
timestamp 1710899220
transform 1 0 2424 0 -1 770
box -8 -3 16 105
use FILL  FILL_1111
timestamp 1710899220
transform 1 0 2352 0 -1 770
box -8 -3 16 105
use FILL  FILL_1112
timestamp 1710899220
transform 1 0 2344 0 -1 770
box -8 -3 16 105
use FILL  FILL_1113
timestamp 1710899220
transform 1 0 2336 0 -1 770
box -8 -3 16 105
use FILL  FILL_1114
timestamp 1710899220
transform 1 0 2136 0 -1 770
box -8 -3 16 105
use FILL  FILL_1115
timestamp 1710899220
transform 1 0 2104 0 -1 770
box -8 -3 16 105
use FILL  FILL_1116
timestamp 1710899220
transform 1 0 2096 0 -1 770
box -8 -3 16 105
use FILL  FILL_1117
timestamp 1710899220
transform 1 0 2088 0 -1 770
box -8 -3 16 105
use FILL  FILL_1118
timestamp 1710899220
transform 1 0 2080 0 -1 770
box -8 -3 16 105
use FILL  FILL_1119
timestamp 1710899220
transform 1 0 2072 0 -1 770
box -8 -3 16 105
use FILL  FILL_1120
timestamp 1710899220
transform 1 0 2064 0 -1 770
box -8 -3 16 105
use FILL  FILL_1121
timestamp 1710899220
transform 1 0 2056 0 -1 770
box -8 -3 16 105
use FILL  FILL_1122
timestamp 1710899220
transform 1 0 1936 0 -1 770
box -8 -3 16 105
use FILL  FILL_1123
timestamp 1710899220
transform 1 0 1872 0 -1 770
box -8 -3 16 105
use FILL  FILL_1124
timestamp 1710899220
transform 1 0 1864 0 -1 770
box -8 -3 16 105
use FILL  FILL_1125
timestamp 1710899220
transform 1 0 1832 0 -1 770
box -8 -3 16 105
use FILL  FILL_1126
timestamp 1710899220
transform 1 0 1824 0 -1 770
box -8 -3 16 105
use FILL  FILL_1127
timestamp 1710899220
transform 1 0 1752 0 -1 770
box -8 -3 16 105
use FILL  FILL_1128
timestamp 1710899220
transform 1 0 1744 0 -1 770
box -8 -3 16 105
use FILL  FILL_1129
timestamp 1710899220
transform 1 0 1648 0 -1 770
box -8 -3 16 105
use FILL  FILL_1130
timestamp 1710899220
transform 1 0 1264 0 -1 770
box -8 -3 16 105
use FILL  FILL_1131
timestamp 1710899220
transform 1 0 1208 0 -1 770
box -8 -3 16 105
use FILL  FILL_1132
timestamp 1710899220
transform 1 0 1200 0 -1 770
box -8 -3 16 105
use FILL  FILL_1133
timestamp 1710899220
transform 1 0 856 0 -1 770
box -8 -3 16 105
use FILL  FILL_1134
timestamp 1710899220
transform 1 0 768 0 -1 770
box -8 -3 16 105
use FILL  FILL_1135
timestamp 1710899220
transform 1 0 712 0 -1 770
box -8 -3 16 105
use FILL  FILL_1136
timestamp 1710899220
transform 1 0 704 0 -1 770
box -8 -3 16 105
use FILL  FILL_1137
timestamp 1710899220
transform 1 0 680 0 -1 770
box -8 -3 16 105
use FILL  FILL_1138
timestamp 1710899220
transform 1 0 672 0 -1 770
box -8 -3 16 105
use FILL  FILL_1139
timestamp 1710899220
transform 1 0 664 0 -1 770
box -8 -3 16 105
use FILL  FILL_1140
timestamp 1710899220
transform 1 0 576 0 -1 770
box -8 -3 16 105
use FILL  FILL_1141
timestamp 1710899220
transform 1 0 512 0 -1 770
box -8 -3 16 105
use FILL  FILL_1142
timestamp 1710899220
transform 1 0 504 0 -1 770
box -8 -3 16 105
use FILL  FILL_1143
timestamp 1710899220
transform 1 0 496 0 -1 770
box -8 -3 16 105
use FILL  FILL_1144
timestamp 1710899220
transform 1 0 488 0 -1 770
box -8 -3 16 105
use FILL  FILL_1145
timestamp 1710899220
transform 1 0 480 0 -1 770
box -8 -3 16 105
use FILL  FILL_1146
timestamp 1710899220
transform 1 0 456 0 -1 770
box -8 -3 16 105
use FILL  FILL_1147
timestamp 1710899220
transform 1 0 448 0 -1 770
box -8 -3 16 105
use FILL  FILL_1148
timestamp 1710899220
transform 1 0 440 0 -1 770
box -8 -3 16 105
use FILL  FILL_1149
timestamp 1710899220
transform 1 0 432 0 -1 770
box -8 -3 16 105
use FILL  FILL_1150
timestamp 1710899220
transform 1 0 424 0 -1 770
box -8 -3 16 105
use FILL  FILL_1151
timestamp 1710899220
transform 1 0 416 0 -1 770
box -8 -3 16 105
use FILL  FILL_1152
timestamp 1710899220
transform 1 0 408 0 -1 770
box -8 -3 16 105
use FILL  FILL_1153
timestamp 1710899220
transform 1 0 400 0 -1 770
box -8 -3 16 105
use FILL  FILL_1154
timestamp 1710899220
transform 1 0 392 0 -1 770
box -8 -3 16 105
use FILL  FILL_1155
timestamp 1710899220
transform 1 0 384 0 -1 770
box -8 -3 16 105
use FILL  FILL_1156
timestamp 1710899220
transform 1 0 376 0 -1 770
box -8 -3 16 105
use FILL  FILL_1157
timestamp 1710899220
transform 1 0 368 0 -1 770
box -8 -3 16 105
use FILL  FILL_1158
timestamp 1710899220
transform 1 0 360 0 -1 770
box -8 -3 16 105
use FILL  FILL_1159
timestamp 1710899220
transform 1 0 352 0 -1 770
box -8 -3 16 105
use FILL  FILL_1160
timestamp 1710899220
transform 1 0 344 0 -1 770
box -8 -3 16 105
use FILL  FILL_1161
timestamp 1710899220
transform 1 0 336 0 -1 770
box -8 -3 16 105
use FILL  FILL_1162
timestamp 1710899220
transform 1 0 328 0 -1 770
box -8 -3 16 105
use FILL  FILL_1163
timestamp 1710899220
transform 1 0 320 0 -1 770
box -8 -3 16 105
use FILL  FILL_1164
timestamp 1710899220
transform 1 0 312 0 -1 770
box -8 -3 16 105
use FILL  FILL_1165
timestamp 1710899220
transform 1 0 304 0 -1 770
box -8 -3 16 105
use FILL  FILL_1166
timestamp 1710899220
transform 1 0 296 0 -1 770
box -8 -3 16 105
use FILL  FILL_1167
timestamp 1710899220
transform 1 0 288 0 -1 770
box -8 -3 16 105
use FILL  FILL_1168
timestamp 1710899220
transform 1 0 280 0 -1 770
box -8 -3 16 105
use FILL  FILL_1169
timestamp 1710899220
transform 1 0 272 0 -1 770
box -8 -3 16 105
use FILL  FILL_1170
timestamp 1710899220
transform 1 0 264 0 -1 770
box -8 -3 16 105
use FILL  FILL_1171
timestamp 1710899220
transform 1 0 256 0 -1 770
box -8 -3 16 105
use FILL  FILL_1172
timestamp 1710899220
transform 1 0 248 0 -1 770
box -8 -3 16 105
use FILL  FILL_1173
timestamp 1710899220
transform 1 0 240 0 -1 770
box -8 -3 16 105
use FILL  FILL_1174
timestamp 1710899220
transform 1 0 232 0 -1 770
box -8 -3 16 105
use FILL  FILL_1175
timestamp 1710899220
transform 1 0 224 0 -1 770
box -8 -3 16 105
use FILL  FILL_1176
timestamp 1710899220
transform 1 0 216 0 -1 770
box -8 -3 16 105
use FILL  FILL_1177
timestamp 1710899220
transform 1 0 208 0 -1 770
box -8 -3 16 105
use FILL  FILL_1178
timestamp 1710899220
transform 1 0 200 0 -1 770
box -8 -3 16 105
use FILL  FILL_1179
timestamp 1710899220
transform 1 0 192 0 -1 770
box -8 -3 16 105
use FILL  FILL_1180
timestamp 1710899220
transform 1 0 184 0 -1 770
box -8 -3 16 105
use FILL  FILL_1181
timestamp 1710899220
transform 1 0 176 0 -1 770
box -8 -3 16 105
use FILL  FILL_1182
timestamp 1710899220
transform 1 0 168 0 -1 770
box -8 -3 16 105
use FILL  FILL_1183
timestamp 1710899220
transform 1 0 160 0 -1 770
box -8 -3 16 105
use FILL  FILL_1184
timestamp 1710899220
transform 1 0 152 0 -1 770
box -8 -3 16 105
use FILL  FILL_1185
timestamp 1710899220
transform 1 0 144 0 -1 770
box -8 -3 16 105
use FILL  FILL_1186
timestamp 1710899220
transform 1 0 136 0 -1 770
box -8 -3 16 105
use FILL  FILL_1187
timestamp 1710899220
transform 1 0 128 0 -1 770
box -8 -3 16 105
use FILL  FILL_1188
timestamp 1710899220
transform 1 0 120 0 -1 770
box -8 -3 16 105
use FILL  FILL_1189
timestamp 1710899220
transform 1 0 112 0 -1 770
box -8 -3 16 105
use FILL  FILL_1190
timestamp 1710899220
transform 1 0 104 0 -1 770
box -8 -3 16 105
use FILL  FILL_1191
timestamp 1710899220
transform 1 0 96 0 -1 770
box -8 -3 16 105
use FILL  FILL_1192
timestamp 1710899220
transform 1 0 88 0 -1 770
box -8 -3 16 105
use FILL  FILL_1193
timestamp 1710899220
transform 1 0 80 0 -1 770
box -8 -3 16 105
use FILL  FILL_1194
timestamp 1710899220
transform 1 0 72 0 -1 770
box -8 -3 16 105
use FILL  FILL_1195
timestamp 1710899220
transform 1 0 168 0 1 570
box -8 -3 16 105
use FILL  FILL_1196
timestamp 1710899220
transform 1 0 160 0 1 570
box -8 -3 16 105
use FILL  FILL_1197
timestamp 1710899220
transform 1 0 152 0 1 570
box -8 -3 16 105
use FILL  FILL_1198
timestamp 1710899220
transform 1 0 144 0 1 570
box -8 -3 16 105
use FILL  FILL_1199
timestamp 1710899220
transform 1 0 136 0 1 570
box -8 -3 16 105
use FILL  FILL_1200
timestamp 1710899220
transform 1 0 128 0 1 570
box -8 -3 16 105
use FILL  FILL_1201
timestamp 1710899220
transform 1 0 120 0 1 570
box -8 -3 16 105
use FILL  FILL_1202
timestamp 1710899220
transform 1 0 112 0 1 570
box -8 -3 16 105
use FILL  FILL_1203
timestamp 1710899220
transform 1 0 104 0 1 570
box -8 -3 16 105
use FILL  FILL_1204
timestamp 1710899220
transform 1 0 96 0 1 570
box -8 -3 16 105
use FILL  FILL_1205
timestamp 1710899220
transform 1 0 88 0 1 570
box -8 -3 16 105
use FILL  FILL_1206
timestamp 1710899220
transform 1 0 80 0 1 570
box -8 -3 16 105
use FILL  FILL_1207
timestamp 1710899220
transform 1 0 72 0 1 570
box -8 -3 16 105
use FILL  FILL_1208
timestamp 1710899220
transform 1 0 2664 0 -1 570
box -8 -3 16 105
use FILL  FILL_1209
timestamp 1710899220
transform 1 0 2656 0 -1 570
box -8 -3 16 105
use FILL  FILL_1210
timestamp 1710899220
transform 1 0 2648 0 -1 570
box -8 -3 16 105
use FILL  FILL_1211
timestamp 1710899220
transform 1 0 2640 0 -1 570
box -8 -3 16 105
use FILL  FILL_1212
timestamp 1710899220
transform 1 0 2632 0 -1 570
box -8 -3 16 105
use FILL  FILL_1213
timestamp 1710899220
transform 1 0 2624 0 -1 570
box -8 -3 16 105
use FILL  FILL_1214
timestamp 1710899220
transform 1 0 2424 0 -1 570
box -8 -3 16 105
use FILL  FILL_1215
timestamp 1710899220
transform 1 0 2320 0 -1 570
box -8 -3 16 105
use FILL  FILL_1216
timestamp 1710899220
transform 1 0 2312 0 -1 570
box -8 -3 16 105
use FILL  FILL_1217
timestamp 1710899220
transform 1 0 2304 0 -1 570
box -8 -3 16 105
use FILL  FILL_1218
timestamp 1710899220
transform 1 0 2296 0 -1 570
box -8 -3 16 105
use FILL  FILL_1219
timestamp 1710899220
transform 1 0 2288 0 -1 570
box -8 -3 16 105
use FILL  FILL_1220
timestamp 1710899220
transform 1 0 2256 0 -1 570
box -8 -3 16 105
use FILL  FILL_1221
timestamp 1710899220
transform 1 0 2248 0 -1 570
box -8 -3 16 105
use FILL  FILL_1222
timestamp 1710899220
transform 1 0 2240 0 -1 570
box -8 -3 16 105
use FILL  FILL_1223
timestamp 1710899220
transform 1 0 2232 0 -1 570
box -8 -3 16 105
use FILL  FILL_1224
timestamp 1710899220
transform 1 0 2224 0 -1 570
box -8 -3 16 105
use FILL  FILL_1225
timestamp 1710899220
transform 1 0 2216 0 -1 570
box -8 -3 16 105
use FILL  FILL_1226
timestamp 1710899220
transform 1 0 2208 0 -1 570
box -8 -3 16 105
use FILL  FILL_1227
timestamp 1710899220
transform 1 0 2200 0 -1 570
box -8 -3 16 105
use FILL  FILL_1228
timestamp 1710899220
transform 1 0 2192 0 -1 570
box -8 -3 16 105
use FILL  FILL_1229
timestamp 1710899220
transform 1 0 2184 0 -1 570
box -8 -3 16 105
use FILL  FILL_1230
timestamp 1710899220
transform 1 0 2176 0 -1 570
box -8 -3 16 105
use FILL  FILL_1231
timestamp 1710899220
transform 1 0 2168 0 -1 570
box -8 -3 16 105
use FILL  FILL_1232
timestamp 1710899220
transform 1 0 2160 0 -1 570
box -8 -3 16 105
use FILL  FILL_1233
timestamp 1710899220
transform 1 0 2152 0 -1 570
box -8 -3 16 105
use FILL  FILL_1234
timestamp 1710899220
transform 1 0 2144 0 -1 570
box -8 -3 16 105
use FILL  FILL_1235
timestamp 1710899220
transform 1 0 2136 0 -1 570
box -8 -3 16 105
use FILL  FILL_1236
timestamp 1710899220
transform 1 0 1944 0 -1 570
box -8 -3 16 105
use FILL  FILL_1237
timestamp 1710899220
transform 1 0 1936 0 -1 570
box -8 -3 16 105
use FILL  FILL_1238
timestamp 1710899220
transform 1 0 1872 0 -1 570
box -8 -3 16 105
use FILL  FILL_1239
timestamp 1710899220
transform 1 0 1816 0 -1 570
box -8 -3 16 105
use FILL  FILL_1240
timestamp 1710899220
transform 1 0 1640 0 -1 570
box -8 -3 16 105
use FILL  FILL_1241
timestamp 1710899220
transform 1 0 1632 0 -1 570
box -8 -3 16 105
use FILL  FILL_1242
timestamp 1710899220
transform 1 0 1520 0 -1 570
box -8 -3 16 105
use FILL  FILL_1243
timestamp 1710899220
transform 1 0 432 0 -1 570
box -8 -3 16 105
use FILL  FILL_1244
timestamp 1710899220
transform 1 0 408 0 -1 570
box -8 -3 16 105
use FILL  FILL_1245
timestamp 1710899220
transform 1 0 400 0 -1 570
box -8 -3 16 105
use FILL  FILL_1246
timestamp 1710899220
transform 1 0 368 0 -1 570
box -8 -3 16 105
use FILL  FILL_1247
timestamp 1710899220
transform 1 0 360 0 -1 570
box -8 -3 16 105
use FILL  FILL_1248
timestamp 1710899220
transform 1 0 296 0 -1 570
box -8 -3 16 105
use FILL  FILL_1249
timestamp 1710899220
transform 1 0 288 0 -1 570
box -8 -3 16 105
use FILL  FILL_1250
timestamp 1710899220
transform 1 0 280 0 -1 570
box -8 -3 16 105
use FILL  FILL_1251
timestamp 1710899220
transform 1 0 272 0 -1 570
box -8 -3 16 105
use FILL  FILL_1252
timestamp 1710899220
transform 1 0 264 0 -1 570
box -8 -3 16 105
use FILL  FILL_1253
timestamp 1710899220
transform 1 0 160 0 -1 570
box -8 -3 16 105
use FILL  FILL_1254
timestamp 1710899220
transform 1 0 152 0 -1 570
box -8 -3 16 105
use FILL  FILL_1255
timestamp 1710899220
transform 1 0 144 0 -1 570
box -8 -3 16 105
use FILL  FILL_1256
timestamp 1710899220
transform 1 0 136 0 -1 570
box -8 -3 16 105
use FILL  FILL_1257
timestamp 1710899220
transform 1 0 128 0 -1 570
box -8 -3 16 105
use FILL  FILL_1258
timestamp 1710899220
transform 1 0 120 0 -1 570
box -8 -3 16 105
use FILL  FILL_1259
timestamp 1710899220
transform 1 0 112 0 -1 570
box -8 -3 16 105
use FILL  FILL_1260
timestamp 1710899220
transform 1 0 104 0 -1 570
box -8 -3 16 105
use FILL  FILL_1261
timestamp 1710899220
transform 1 0 96 0 -1 570
box -8 -3 16 105
use FILL  FILL_1262
timestamp 1710899220
transform 1 0 88 0 -1 570
box -8 -3 16 105
use FILL  FILL_1263
timestamp 1710899220
transform 1 0 80 0 -1 570
box -8 -3 16 105
use FILL  FILL_1264
timestamp 1710899220
transform 1 0 72 0 -1 570
box -8 -3 16 105
use FILL  FILL_1265
timestamp 1710899220
transform 1 0 2568 0 1 370
box -8 -3 16 105
use FILL  FILL_1266
timestamp 1710899220
transform 1 0 2560 0 1 370
box -8 -3 16 105
use FILL  FILL_1267
timestamp 1710899220
transform 1 0 2552 0 1 370
box -8 -3 16 105
use FILL  FILL_1268
timestamp 1710899220
transform 1 0 2544 0 1 370
box -8 -3 16 105
use FILL  FILL_1269
timestamp 1710899220
transform 1 0 2536 0 1 370
box -8 -3 16 105
use FILL  FILL_1270
timestamp 1710899220
transform 1 0 2528 0 1 370
box -8 -3 16 105
use FILL  FILL_1271
timestamp 1710899220
transform 1 0 2520 0 1 370
box -8 -3 16 105
use FILL  FILL_1272
timestamp 1710899220
transform 1 0 2496 0 1 370
box -8 -3 16 105
use FILL  FILL_1273
timestamp 1710899220
transform 1 0 2488 0 1 370
box -8 -3 16 105
use FILL  FILL_1274
timestamp 1710899220
transform 1 0 2480 0 1 370
box -8 -3 16 105
use FILL  FILL_1275
timestamp 1710899220
transform 1 0 2472 0 1 370
box -8 -3 16 105
use FILL  FILL_1276
timestamp 1710899220
transform 1 0 2464 0 1 370
box -8 -3 16 105
use FILL  FILL_1277
timestamp 1710899220
transform 1 0 2456 0 1 370
box -8 -3 16 105
use FILL  FILL_1278
timestamp 1710899220
transform 1 0 2424 0 1 370
box -8 -3 16 105
use FILL  FILL_1279
timestamp 1710899220
transform 1 0 2416 0 1 370
box -8 -3 16 105
use FILL  FILL_1280
timestamp 1710899220
transform 1 0 2408 0 1 370
box -8 -3 16 105
use FILL  FILL_1281
timestamp 1710899220
transform 1 0 2400 0 1 370
box -8 -3 16 105
use FILL  FILL_1282
timestamp 1710899220
transform 1 0 2392 0 1 370
box -8 -3 16 105
use FILL  FILL_1283
timestamp 1710899220
transform 1 0 2384 0 1 370
box -8 -3 16 105
use FILL  FILL_1284
timestamp 1710899220
transform 1 0 2344 0 1 370
box -8 -3 16 105
use FILL  FILL_1285
timestamp 1710899220
transform 1 0 2336 0 1 370
box -8 -3 16 105
use FILL  FILL_1286
timestamp 1710899220
transform 1 0 2296 0 1 370
box -8 -3 16 105
use FILL  FILL_1287
timestamp 1710899220
transform 1 0 2288 0 1 370
box -8 -3 16 105
use FILL  FILL_1288
timestamp 1710899220
transform 1 0 2184 0 1 370
box -8 -3 16 105
use FILL  FILL_1289
timestamp 1710899220
transform 1 0 2080 0 1 370
box -8 -3 16 105
use FILL  FILL_1290
timestamp 1710899220
transform 1 0 2072 0 1 370
box -8 -3 16 105
use FILL  FILL_1291
timestamp 1710899220
transform 1 0 2064 0 1 370
box -8 -3 16 105
use FILL  FILL_1292
timestamp 1710899220
transform 1 0 2056 0 1 370
box -8 -3 16 105
use FILL  FILL_1293
timestamp 1710899220
transform 1 0 2048 0 1 370
box -8 -3 16 105
use FILL  FILL_1294
timestamp 1710899220
transform 1 0 2040 0 1 370
box -8 -3 16 105
use FILL  FILL_1295
timestamp 1710899220
transform 1 0 2032 0 1 370
box -8 -3 16 105
use FILL  FILL_1296
timestamp 1710899220
transform 1 0 1960 0 1 370
box -8 -3 16 105
use FILL  FILL_1297
timestamp 1710899220
transform 1 0 1824 0 1 370
box -8 -3 16 105
use FILL  FILL_1298
timestamp 1710899220
transform 1 0 1816 0 1 370
box -8 -3 16 105
use FILL  FILL_1299
timestamp 1710899220
transform 1 0 1744 0 1 370
box -8 -3 16 105
use FILL  FILL_1300
timestamp 1710899220
transform 1 0 1736 0 1 370
box -8 -3 16 105
use FILL  FILL_1301
timestamp 1710899220
transform 1 0 1544 0 1 370
box -8 -3 16 105
use FILL  FILL_1302
timestamp 1710899220
transform 1 0 1464 0 1 370
box -8 -3 16 105
use FILL  FILL_1303
timestamp 1710899220
transform 1 0 1456 0 1 370
box -8 -3 16 105
use FILL  FILL_1304
timestamp 1710899220
transform 1 0 1368 0 1 370
box -8 -3 16 105
use FILL  FILL_1305
timestamp 1710899220
transform 1 0 1312 0 1 370
box -8 -3 16 105
use FILL  FILL_1306
timestamp 1710899220
transform 1 0 1304 0 1 370
box -8 -3 16 105
use FILL  FILL_1307
timestamp 1710899220
transform 1 0 1296 0 1 370
box -8 -3 16 105
use FILL  FILL_1308
timestamp 1710899220
transform 1 0 1288 0 1 370
box -8 -3 16 105
use FILL  FILL_1309
timestamp 1710899220
transform 1 0 1224 0 1 370
box -8 -3 16 105
use FILL  FILL_1310
timestamp 1710899220
transform 1 0 1216 0 1 370
box -8 -3 16 105
use FILL  FILL_1311
timestamp 1710899220
transform 1 0 1208 0 1 370
box -8 -3 16 105
use FILL  FILL_1312
timestamp 1710899220
transform 1 0 1200 0 1 370
box -8 -3 16 105
use FILL  FILL_1313
timestamp 1710899220
transform 1 0 1176 0 1 370
box -8 -3 16 105
use FILL  FILL_1314
timestamp 1710899220
transform 1 0 1168 0 1 370
box -8 -3 16 105
use FILL  FILL_1315
timestamp 1710899220
transform 1 0 1160 0 1 370
box -8 -3 16 105
use FILL  FILL_1316
timestamp 1710899220
transform 1 0 1152 0 1 370
box -8 -3 16 105
use FILL  FILL_1317
timestamp 1710899220
transform 1 0 1144 0 1 370
box -8 -3 16 105
use FILL  FILL_1318
timestamp 1710899220
transform 1 0 1136 0 1 370
box -8 -3 16 105
use FILL  FILL_1319
timestamp 1710899220
transform 1 0 1128 0 1 370
box -8 -3 16 105
use FILL  FILL_1320
timestamp 1710899220
transform 1 0 1072 0 1 370
box -8 -3 16 105
use FILL  FILL_1321
timestamp 1710899220
transform 1 0 1032 0 1 370
box -8 -3 16 105
use FILL  FILL_1322
timestamp 1710899220
transform 1 0 1024 0 1 370
box -8 -3 16 105
use FILL  FILL_1323
timestamp 1710899220
transform 1 0 1016 0 1 370
box -8 -3 16 105
use FILL  FILL_1324
timestamp 1710899220
transform 1 0 1008 0 1 370
box -8 -3 16 105
use FILL  FILL_1325
timestamp 1710899220
transform 1 0 936 0 1 370
box -8 -3 16 105
use FILL  FILL_1326
timestamp 1710899220
transform 1 0 928 0 1 370
box -8 -3 16 105
use FILL  FILL_1327
timestamp 1710899220
transform 1 0 920 0 1 370
box -8 -3 16 105
use FILL  FILL_1328
timestamp 1710899220
transform 1 0 912 0 1 370
box -8 -3 16 105
use FILL  FILL_1329
timestamp 1710899220
transform 1 0 904 0 1 370
box -8 -3 16 105
use FILL  FILL_1330
timestamp 1710899220
transform 1 0 816 0 1 370
box -8 -3 16 105
use FILL  FILL_1331
timestamp 1710899220
transform 1 0 808 0 1 370
box -8 -3 16 105
use FILL  FILL_1332
timestamp 1710899220
transform 1 0 728 0 1 370
box -8 -3 16 105
use FILL  FILL_1333
timestamp 1710899220
transform 1 0 648 0 1 370
box -8 -3 16 105
use FILL  FILL_1334
timestamp 1710899220
transform 1 0 640 0 1 370
box -8 -3 16 105
use FILL  FILL_1335
timestamp 1710899220
transform 1 0 632 0 1 370
box -8 -3 16 105
use FILL  FILL_1336
timestamp 1710899220
transform 1 0 576 0 1 370
box -8 -3 16 105
use FILL  FILL_1337
timestamp 1710899220
transform 1 0 504 0 1 370
box -8 -3 16 105
use FILL  FILL_1338
timestamp 1710899220
transform 1 0 496 0 1 370
box -8 -3 16 105
use FILL  FILL_1339
timestamp 1710899220
transform 1 0 392 0 1 370
box -8 -3 16 105
use FILL  FILL_1340
timestamp 1710899220
transform 1 0 328 0 1 370
box -8 -3 16 105
use FILL  FILL_1341
timestamp 1710899220
transform 1 0 224 0 1 370
box -8 -3 16 105
use FILL  FILL_1342
timestamp 1710899220
transform 1 0 216 0 1 370
box -8 -3 16 105
use FILL  FILL_1343
timestamp 1710899220
transform 1 0 208 0 1 370
box -8 -3 16 105
use FILL  FILL_1344
timestamp 1710899220
transform 1 0 200 0 1 370
box -8 -3 16 105
use FILL  FILL_1345
timestamp 1710899220
transform 1 0 192 0 1 370
box -8 -3 16 105
use FILL  FILL_1346
timestamp 1710899220
transform 1 0 184 0 1 370
box -8 -3 16 105
use FILL  FILL_1347
timestamp 1710899220
transform 1 0 176 0 1 370
box -8 -3 16 105
use FILL  FILL_1348
timestamp 1710899220
transform 1 0 168 0 1 370
box -8 -3 16 105
use FILL  FILL_1349
timestamp 1710899220
transform 1 0 160 0 1 370
box -8 -3 16 105
use FILL  FILL_1350
timestamp 1710899220
transform 1 0 152 0 1 370
box -8 -3 16 105
use FILL  FILL_1351
timestamp 1710899220
transform 1 0 144 0 1 370
box -8 -3 16 105
use FILL  FILL_1352
timestamp 1710899220
transform 1 0 136 0 1 370
box -8 -3 16 105
use FILL  FILL_1353
timestamp 1710899220
transform 1 0 128 0 1 370
box -8 -3 16 105
use FILL  FILL_1354
timestamp 1710899220
transform 1 0 120 0 1 370
box -8 -3 16 105
use FILL  FILL_1355
timestamp 1710899220
transform 1 0 112 0 1 370
box -8 -3 16 105
use FILL  FILL_1356
timestamp 1710899220
transform 1 0 104 0 1 370
box -8 -3 16 105
use FILL  FILL_1357
timestamp 1710899220
transform 1 0 96 0 1 370
box -8 -3 16 105
use FILL  FILL_1358
timestamp 1710899220
transform 1 0 88 0 1 370
box -8 -3 16 105
use FILL  FILL_1359
timestamp 1710899220
transform 1 0 80 0 1 370
box -8 -3 16 105
use FILL  FILL_1360
timestamp 1710899220
transform 1 0 72 0 1 370
box -8 -3 16 105
use FILL  FILL_1361
timestamp 1710899220
transform 1 0 2664 0 -1 370
box -8 -3 16 105
use FILL  FILL_1362
timestamp 1710899220
transform 1 0 2656 0 -1 370
box -8 -3 16 105
use FILL  FILL_1363
timestamp 1710899220
transform 1 0 2648 0 -1 370
box -8 -3 16 105
use FILL  FILL_1364
timestamp 1710899220
transform 1 0 2640 0 -1 370
box -8 -3 16 105
use FILL  FILL_1365
timestamp 1710899220
transform 1 0 2576 0 -1 370
box -8 -3 16 105
use FILL  FILL_1366
timestamp 1710899220
transform 1 0 2568 0 -1 370
box -8 -3 16 105
use FILL  FILL_1367
timestamp 1710899220
transform 1 0 2456 0 -1 370
box -8 -3 16 105
use FILL  FILL_1368
timestamp 1710899220
transform 1 0 2448 0 -1 370
box -8 -3 16 105
use FILL  FILL_1369
timestamp 1710899220
transform 1 0 2408 0 -1 370
box -8 -3 16 105
use FILL  FILL_1370
timestamp 1710899220
transform 1 0 2400 0 -1 370
box -8 -3 16 105
use FILL  FILL_1371
timestamp 1710899220
transform 1 0 2392 0 -1 370
box -8 -3 16 105
use FILL  FILL_1372
timestamp 1710899220
transform 1 0 2328 0 -1 370
box -8 -3 16 105
use FILL  FILL_1373
timestamp 1710899220
transform 1 0 2320 0 -1 370
box -8 -3 16 105
use FILL  FILL_1374
timestamp 1710899220
transform 1 0 2312 0 -1 370
box -8 -3 16 105
use FILL  FILL_1375
timestamp 1710899220
transform 1 0 2304 0 -1 370
box -8 -3 16 105
use FILL  FILL_1376
timestamp 1710899220
transform 1 0 2232 0 -1 370
box -8 -3 16 105
use FILL  FILL_1377
timestamp 1710899220
transform 1 0 2224 0 -1 370
box -8 -3 16 105
use FILL  FILL_1378
timestamp 1710899220
transform 1 0 448 0 -1 370
box -8 -3 16 105
use FILL  FILL_1379
timestamp 1710899220
transform 1 0 384 0 -1 370
box -8 -3 16 105
use FILL  FILL_1380
timestamp 1710899220
transform 1 0 376 0 -1 370
box -8 -3 16 105
use FILL  FILL_1381
timestamp 1710899220
transform 1 0 288 0 -1 370
box -8 -3 16 105
use FILL  FILL_1382
timestamp 1710899220
transform 1 0 280 0 -1 370
box -8 -3 16 105
use FILL  FILL_1383
timestamp 1710899220
transform 1 0 272 0 -1 370
box -8 -3 16 105
use FILL  FILL_1384
timestamp 1710899220
transform 1 0 264 0 -1 370
box -8 -3 16 105
use FILL  FILL_1385
timestamp 1710899220
transform 1 0 160 0 -1 370
box -8 -3 16 105
use FILL  FILL_1386
timestamp 1710899220
transform 1 0 152 0 -1 370
box -8 -3 16 105
use FILL  FILL_1387
timestamp 1710899220
transform 1 0 144 0 -1 370
box -8 -3 16 105
use FILL  FILL_1388
timestamp 1710899220
transform 1 0 136 0 -1 370
box -8 -3 16 105
use FILL  FILL_1389
timestamp 1710899220
transform 1 0 128 0 -1 370
box -8 -3 16 105
use FILL  FILL_1390
timestamp 1710899220
transform 1 0 120 0 -1 370
box -8 -3 16 105
use FILL  FILL_1391
timestamp 1710899220
transform 1 0 112 0 -1 370
box -8 -3 16 105
use FILL  FILL_1392
timestamp 1710899220
transform 1 0 104 0 -1 370
box -8 -3 16 105
use FILL  FILL_1393
timestamp 1710899220
transform 1 0 96 0 -1 370
box -8 -3 16 105
use FILL  FILL_1394
timestamp 1710899220
transform 1 0 88 0 -1 370
box -8 -3 16 105
use FILL  FILL_1395
timestamp 1710899220
transform 1 0 80 0 -1 370
box -8 -3 16 105
use FILL  FILL_1396
timestamp 1710899220
transform 1 0 72 0 -1 370
box -8 -3 16 105
use FILL  FILL_1397
timestamp 1710899220
transform 1 0 2488 0 1 170
box -8 -3 16 105
use FILL  FILL_1398
timestamp 1710899220
transform 1 0 2400 0 1 170
box -8 -3 16 105
use FILL  FILL_1399
timestamp 1710899220
transform 1 0 2344 0 1 170
box -8 -3 16 105
use FILL  FILL_1400
timestamp 1710899220
transform 1 0 2336 0 1 170
box -8 -3 16 105
use FILL  FILL_1401
timestamp 1710899220
transform 1 0 2240 0 1 170
box -8 -3 16 105
use FILL  FILL_1402
timestamp 1710899220
transform 1 0 2176 0 1 170
box -8 -3 16 105
use FILL  FILL_1403
timestamp 1710899220
transform 1 0 2168 0 1 170
box -8 -3 16 105
use FILL  FILL_1404
timestamp 1710899220
transform 1 0 2064 0 1 170
box -8 -3 16 105
use FILL  FILL_1405
timestamp 1710899220
transform 1 0 2056 0 1 170
box -8 -3 16 105
use FILL  FILL_1406
timestamp 1710899220
transform 1 0 2048 0 1 170
box -8 -3 16 105
use FILL  FILL_1407
timestamp 1710899220
transform 1 0 2040 0 1 170
box -8 -3 16 105
use FILL  FILL_1408
timestamp 1710899220
transform 1 0 2032 0 1 170
box -8 -3 16 105
use FILL  FILL_1409
timestamp 1710899220
transform 1 0 2024 0 1 170
box -8 -3 16 105
use FILL  FILL_1410
timestamp 1710899220
transform 1 0 2016 0 1 170
box -8 -3 16 105
use FILL  FILL_1411
timestamp 1710899220
transform 1 0 2008 0 1 170
box -8 -3 16 105
use FILL  FILL_1412
timestamp 1710899220
transform 1 0 1944 0 1 170
box -8 -3 16 105
use FILL  FILL_1413
timestamp 1710899220
transform 1 0 1840 0 1 170
box -8 -3 16 105
use FILL  FILL_1414
timestamp 1710899220
transform 1 0 1832 0 1 170
box -8 -3 16 105
use FILL  FILL_1415
timestamp 1710899220
transform 1 0 1824 0 1 170
box -8 -3 16 105
use FILL  FILL_1416
timestamp 1710899220
transform 1 0 1816 0 1 170
box -8 -3 16 105
use FILL  FILL_1417
timestamp 1710899220
transform 1 0 1808 0 1 170
box -8 -3 16 105
use FILL  FILL_1418
timestamp 1710899220
transform 1 0 1752 0 1 170
box -8 -3 16 105
use FILL  FILL_1419
timestamp 1710899220
transform 1 0 1744 0 1 170
box -8 -3 16 105
use FILL  FILL_1420
timestamp 1710899220
transform 1 0 1736 0 1 170
box -8 -3 16 105
use FILL  FILL_1421
timestamp 1710899220
transform 1 0 1728 0 1 170
box -8 -3 16 105
use FILL  FILL_1422
timestamp 1710899220
transform 1 0 1720 0 1 170
box -8 -3 16 105
use FILL  FILL_1423
timestamp 1710899220
transform 1 0 1712 0 1 170
box -8 -3 16 105
use FILL  FILL_1424
timestamp 1710899220
transform 1 0 1648 0 1 170
box -8 -3 16 105
use FILL  FILL_1425
timestamp 1710899220
transform 1 0 1640 0 1 170
box -8 -3 16 105
use FILL  FILL_1426
timestamp 1710899220
transform 1 0 1632 0 1 170
box -8 -3 16 105
use FILL  FILL_1427
timestamp 1710899220
transform 1 0 1568 0 1 170
box -8 -3 16 105
use FILL  FILL_1428
timestamp 1710899220
transform 1 0 1416 0 1 170
box -8 -3 16 105
use FILL  FILL_1429
timestamp 1710899220
transform 1 0 1408 0 1 170
box -8 -3 16 105
use FILL  FILL_1430
timestamp 1710899220
transform 1 0 1352 0 1 170
box -8 -3 16 105
use FILL  FILL_1431
timestamp 1710899220
transform 1 0 1344 0 1 170
box -8 -3 16 105
use FILL  FILL_1432
timestamp 1710899220
transform 1 0 1336 0 1 170
box -8 -3 16 105
use FILL  FILL_1433
timestamp 1710899220
transform 1 0 1296 0 1 170
box -8 -3 16 105
use FILL  FILL_1434
timestamp 1710899220
transform 1 0 1216 0 1 170
box -8 -3 16 105
use FILL  FILL_1435
timestamp 1710899220
transform 1 0 1208 0 1 170
box -8 -3 16 105
use FILL  FILL_1436
timestamp 1710899220
transform 1 0 1200 0 1 170
box -8 -3 16 105
use FILL  FILL_1437
timestamp 1710899220
transform 1 0 960 0 1 170
box -8 -3 16 105
use FILL  FILL_1438
timestamp 1710899220
transform 1 0 880 0 1 170
box -8 -3 16 105
use FILL  FILL_1439
timestamp 1710899220
transform 1 0 872 0 1 170
box -8 -3 16 105
use FILL  FILL_1440
timestamp 1710899220
transform 1 0 864 0 1 170
box -8 -3 16 105
use FILL  FILL_1441
timestamp 1710899220
transform 1 0 792 0 1 170
box -8 -3 16 105
use FILL  FILL_1442
timestamp 1710899220
transform 1 0 696 0 1 170
box -8 -3 16 105
use FILL  FILL_1443
timestamp 1710899220
transform 1 0 640 0 1 170
box -8 -3 16 105
use FILL  FILL_1444
timestamp 1710899220
transform 1 0 584 0 1 170
box -8 -3 16 105
use FILL  FILL_1445
timestamp 1710899220
transform 1 0 576 0 1 170
box -8 -3 16 105
use FILL  FILL_1446
timestamp 1710899220
transform 1 0 480 0 1 170
box -8 -3 16 105
use FILL  FILL_1447
timestamp 1710899220
transform 1 0 472 0 1 170
box -8 -3 16 105
use FILL  FILL_1448
timestamp 1710899220
transform 1 0 464 0 1 170
box -8 -3 16 105
use FILL  FILL_1449
timestamp 1710899220
transform 1 0 224 0 1 170
box -8 -3 16 105
use FILL  FILL_1450
timestamp 1710899220
transform 1 0 216 0 1 170
box -8 -3 16 105
use FILL  FILL_1451
timestamp 1710899220
transform 1 0 208 0 1 170
box -8 -3 16 105
use FILL  FILL_1452
timestamp 1710899220
transform 1 0 200 0 1 170
box -8 -3 16 105
use FILL  FILL_1453
timestamp 1710899220
transform 1 0 192 0 1 170
box -8 -3 16 105
use FILL  FILL_1454
timestamp 1710899220
transform 1 0 184 0 1 170
box -8 -3 16 105
use FILL  FILL_1455
timestamp 1710899220
transform 1 0 176 0 1 170
box -8 -3 16 105
use FILL  FILL_1456
timestamp 1710899220
transform 1 0 168 0 1 170
box -8 -3 16 105
use FILL  FILL_1457
timestamp 1710899220
transform 1 0 160 0 1 170
box -8 -3 16 105
use FILL  FILL_1458
timestamp 1710899220
transform 1 0 152 0 1 170
box -8 -3 16 105
use FILL  FILL_1459
timestamp 1710899220
transform 1 0 144 0 1 170
box -8 -3 16 105
use FILL  FILL_1460
timestamp 1710899220
transform 1 0 136 0 1 170
box -8 -3 16 105
use FILL  FILL_1461
timestamp 1710899220
transform 1 0 128 0 1 170
box -8 -3 16 105
use FILL  FILL_1462
timestamp 1710899220
transform 1 0 120 0 1 170
box -8 -3 16 105
use FILL  FILL_1463
timestamp 1710899220
transform 1 0 112 0 1 170
box -8 -3 16 105
use FILL  FILL_1464
timestamp 1710899220
transform 1 0 104 0 1 170
box -8 -3 16 105
use FILL  FILL_1465
timestamp 1710899220
transform 1 0 96 0 1 170
box -8 -3 16 105
use FILL  FILL_1466
timestamp 1710899220
transform 1 0 88 0 1 170
box -8 -3 16 105
use FILL  FILL_1467
timestamp 1710899220
transform 1 0 80 0 1 170
box -8 -3 16 105
use FILL  FILL_1468
timestamp 1710899220
transform 1 0 72 0 1 170
box -8 -3 16 105
use FILL  FILL_1469
timestamp 1710899220
transform 1 0 2664 0 -1 170
box -8 -3 16 105
use FILL  FILL_1470
timestamp 1710899220
transform 1 0 2656 0 -1 170
box -8 -3 16 105
use FILL  FILL_1471
timestamp 1710899220
transform 1 0 2648 0 -1 170
box -8 -3 16 105
use FILL  FILL_1472
timestamp 1710899220
transform 1 0 2640 0 -1 170
box -8 -3 16 105
use FILL  FILL_1473
timestamp 1710899220
transform 1 0 2632 0 -1 170
box -8 -3 16 105
use FILL  FILL_1474
timestamp 1710899220
transform 1 0 2624 0 -1 170
box -8 -3 16 105
use FILL  FILL_1475
timestamp 1710899220
transform 1 0 2616 0 -1 170
box -8 -3 16 105
use FILL  FILL_1476
timestamp 1710899220
transform 1 0 2608 0 -1 170
box -8 -3 16 105
use FILL  FILL_1477
timestamp 1710899220
transform 1 0 2600 0 -1 170
box -8 -3 16 105
use FILL  FILL_1478
timestamp 1710899220
transform 1 0 2592 0 -1 170
box -8 -3 16 105
use FILL  FILL_1479
timestamp 1710899220
transform 1 0 2584 0 -1 170
box -8 -3 16 105
use FILL  FILL_1480
timestamp 1710899220
transform 1 0 2576 0 -1 170
box -8 -3 16 105
use FILL  FILL_1481
timestamp 1710899220
transform 1 0 2568 0 -1 170
box -8 -3 16 105
use FILL  FILL_1482
timestamp 1710899220
transform 1 0 2560 0 -1 170
box -8 -3 16 105
use FILL  FILL_1483
timestamp 1710899220
transform 1 0 2552 0 -1 170
box -8 -3 16 105
use FILL  FILL_1484
timestamp 1710899220
transform 1 0 2544 0 -1 170
box -8 -3 16 105
use FILL  FILL_1485
timestamp 1710899220
transform 1 0 2536 0 -1 170
box -8 -3 16 105
use FILL  FILL_1486
timestamp 1710899220
transform 1 0 2528 0 -1 170
box -8 -3 16 105
use FILL  FILL_1487
timestamp 1710899220
transform 1 0 2520 0 -1 170
box -8 -3 16 105
use FILL  FILL_1488
timestamp 1710899220
transform 1 0 2512 0 -1 170
box -8 -3 16 105
use FILL  FILL_1489
timestamp 1710899220
transform 1 0 2504 0 -1 170
box -8 -3 16 105
use FILL  FILL_1490
timestamp 1710899220
transform 1 0 2496 0 -1 170
box -8 -3 16 105
use FILL  FILL_1491
timestamp 1710899220
transform 1 0 2488 0 -1 170
box -8 -3 16 105
use FILL  FILL_1492
timestamp 1710899220
transform 1 0 2480 0 -1 170
box -8 -3 16 105
use FILL  FILL_1493
timestamp 1710899220
transform 1 0 2472 0 -1 170
box -8 -3 16 105
use FILL  FILL_1494
timestamp 1710899220
transform 1 0 2464 0 -1 170
box -8 -3 16 105
use FILL  FILL_1495
timestamp 1710899220
transform 1 0 2456 0 -1 170
box -8 -3 16 105
use FILL  FILL_1496
timestamp 1710899220
transform 1 0 2448 0 -1 170
box -8 -3 16 105
use FILL  FILL_1497
timestamp 1710899220
transform 1 0 2440 0 -1 170
box -8 -3 16 105
use FILL  FILL_1498
timestamp 1710899220
transform 1 0 2432 0 -1 170
box -8 -3 16 105
use FILL  FILL_1499
timestamp 1710899220
transform 1 0 2424 0 -1 170
box -8 -3 16 105
use FILL  FILL_1500
timestamp 1710899220
transform 1 0 2416 0 -1 170
box -8 -3 16 105
use FILL  FILL_1501
timestamp 1710899220
transform 1 0 2408 0 -1 170
box -8 -3 16 105
use FILL  FILL_1502
timestamp 1710899220
transform 1 0 2400 0 -1 170
box -8 -3 16 105
use FILL  FILL_1503
timestamp 1710899220
transform 1 0 2392 0 -1 170
box -8 -3 16 105
use FILL  FILL_1504
timestamp 1710899220
transform 1 0 2384 0 -1 170
box -8 -3 16 105
use FILL  FILL_1505
timestamp 1710899220
transform 1 0 2376 0 -1 170
box -8 -3 16 105
use FILL  FILL_1506
timestamp 1710899220
transform 1 0 2368 0 -1 170
box -8 -3 16 105
use FILL  FILL_1507
timestamp 1710899220
transform 1 0 2360 0 -1 170
box -8 -3 16 105
use FILL  FILL_1508
timestamp 1710899220
transform 1 0 2352 0 -1 170
box -8 -3 16 105
use FILL  FILL_1509
timestamp 1710899220
transform 1 0 2344 0 -1 170
box -8 -3 16 105
use FILL  FILL_1510
timestamp 1710899220
transform 1 0 2336 0 -1 170
box -8 -3 16 105
use FILL  FILL_1511
timestamp 1710899220
transform 1 0 2328 0 -1 170
box -8 -3 16 105
use FILL  FILL_1512
timestamp 1710899220
transform 1 0 2320 0 -1 170
box -8 -3 16 105
use FILL  FILL_1513
timestamp 1710899220
transform 1 0 2312 0 -1 170
box -8 -3 16 105
use FILL  FILL_1514
timestamp 1710899220
transform 1 0 2304 0 -1 170
box -8 -3 16 105
use FILL  FILL_1515
timestamp 1710899220
transform 1 0 2296 0 -1 170
box -8 -3 16 105
use FILL  FILL_1516
timestamp 1710899220
transform 1 0 2288 0 -1 170
box -8 -3 16 105
use FILL  FILL_1517
timestamp 1710899220
transform 1 0 2280 0 -1 170
box -8 -3 16 105
use FILL  FILL_1518
timestamp 1710899220
transform 1 0 2272 0 -1 170
box -8 -3 16 105
use FILL  FILL_1519
timestamp 1710899220
transform 1 0 2264 0 -1 170
box -8 -3 16 105
use FILL  FILL_1520
timestamp 1710899220
transform 1 0 2256 0 -1 170
box -8 -3 16 105
use FILL  FILL_1521
timestamp 1710899220
transform 1 0 2248 0 -1 170
box -8 -3 16 105
use FILL  FILL_1522
timestamp 1710899220
transform 1 0 2240 0 -1 170
box -8 -3 16 105
use FILL  FILL_1523
timestamp 1710899220
transform 1 0 2232 0 -1 170
box -8 -3 16 105
use FILL  FILL_1524
timestamp 1710899220
transform 1 0 2224 0 -1 170
box -8 -3 16 105
use FILL  FILL_1525
timestamp 1710899220
transform 1 0 2216 0 -1 170
box -8 -3 16 105
use FILL  FILL_1526
timestamp 1710899220
transform 1 0 2208 0 -1 170
box -8 -3 16 105
use FILL  FILL_1527
timestamp 1710899220
transform 1 0 2200 0 -1 170
box -8 -3 16 105
use FILL  FILL_1528
timestamp 1710899220
transform 1 0 2192 0 -1 170
box -8 -3 16 105
use FILL  FILL_1529
timestamp 1710899220
transform 1 0 2184 0 -1 170
box -8 -3 16 105
use FILL  FILL_1530
timestamp 1710899220
transform 1 0 2176 0 -1 170
box -8 -3 16 105
use FILL  FILL_1531
timestamp 1710899220
transform 1 0 2168 0 -1 170
box -8 -3 16 105
use FILL  FILL_1532
timestamp 1710899220
transform 1 0 2160 0 -1 170
box -8 -3 16 105
use FILL  FILL_1533
timestamp 1710899220
transform 1 0 2152 0 -1 170
box -8 -3 16 105
use FILL  FILL_1534
timestamp 1710899220
transform 1 0 2144 0 -1 170
box -8 -3 16 105
use FILL  FILL_1535
timestamp 1710899220
transform 1 0 2136 0 -1 170
box -8 -3 16 105
use FILL  FILL_1536
timestamp 1710899220
transform 1 0 2128 0 -1 170
box -8 -3 16 105
use FILL  FILL_1537
timestamp 1710899220
transform 1 0 2120 0 -1 170
box -8 -3 16 105
use FILL  FILL_1538
timestamp 1710899220
transform 1 0 2112 0 -1 170
box -8 -3 16 105
use FILL  FILL_1539
timestamp 1710899220
transform 1 0 2104 0 -1 170
box -8 -3 16 105
use FILL  FILL_1540
timestamp 1710899220
transform 1 0 2096 0 -1 170
box -8 -3 16 105
use FILL  FILL_1541
timestamp 1710899220
transform 1 0 2088 0 -1 170
box -8 -3 16 105
use FILL  FILL_1542
timestamp 1710899220
transform 1 0 2080 0 -1 170
box -8 -3 16 105
use FILL  FILL_1543
timestamp 1710899220
transform 1 0 2072 0 -1 170
box -8 -3 16 105
use FILL  FILL_1544
timestamp 1710899220
transform 1 0 2064 0 -1 170
box -8 -3 16 105
use FILL  FILL_1545
timestamp 1710899220
transform 1 0 2056 0 -1 170
box -8 -3 16 105
use FILL  FILL_1546
timestamp 1710899220
transform 1 0 2048 0 -1 170
box -8 -3 16 105
use FILL  FILL_1547
timestamp 1710899220
transform 1 0 2040 0 -1 170
box -8 -3 16 105
use FILL  FILL_1548
timestamp 1710899220
transform 1 0 1936 0 -1 170
box -8 -3 16 105
use FILL  FILL_1549
timestamp 1710899220
transform 1 0 1928 0 -1 170
box -8 -3 16 105
use FILL  FILL_1550
timestamp 1710899220
transform 1 0 1920 0 -1 170
box -8 -3 16 105
use FILL  FILL_1551
timestamp 1710899220
transform 1 0 1912 0 -1 170
box -8 -3 16 105
use FILL  FILL_1552
timestamp 1710899220
transform 1 0 1904 0 -1 170
box -8 -3 16 105
use FILL  FILL_1553
timestamp 1710899220
transform 1 0 1896 0 -1 170
box -8 -3 16 105
use FILL  FILL_1554
timestamp 1710899220
transform 1 0 1888 0 -1 170
box -8 -3 16 105
use FILL  FILL_1555
timestamp 1710899220
transform 1 0 1880 0 -1 170
box -8 -3 16 105
use FILL  FILL_1556
timestamp 1710899220
transform 1 0 1872 0 -1 170
box -8 -3 16 105
use FILL  FILL_1557
timestamp 1710899220
transform 1 0 1864 0 -1 170
box -8 -3 16 105
use FILL  FILL_1558
timestamp 1710899220
transform 1 0 1856 0 -1 170
box -8 -3 16 105
use FILL  FILL_1559
timestamp 1710899220
transform 1 0 1656 0 -1 170
box -8 -3 16 105
use FILL  FILL_1560
timestamp 1710899220
transform 1 0 1648 0 -1 170
box -8 -3 16 105
use FILL  FILL_1561
timestamp 1710899220
transform 1 0 1544 0 -1 170
box -8 -3 16 105
use FILL  FILL_1562
timestamp 1710899220
transform 1 0 1536 0 -1 170
box -8 -3 16 105
use FILL  FILL_1563
timestamp 1710899220
transform 1 0 1528 0 -1 170
box -8 -3 16 105
use FILL  FILL_1564
timestamp 1710899220
transform 1 0 1520 0 -1 170
box -8 -3 16 105
use FILL  FILL_1565
timestamp 1710899220
transform 1 0 1512 0 -1 170
box -8 -3 16 105
use FILL  FILL_1566
timestamp 1710899220
transform 1 0 1504 0 -1 170
box -8 -3 16 105
use FILL  FILL_1567
timestamp 1710899220
transform 1 0 1496 0 -1 170
box -8 -3 16 105
use FILL  FILL_1568
timestamp 1710899220
transform 1 0 1488 0 -1 170
box -8 -3 16 105
use FILL  FILL_1569
timestamp 1710899220
transform 1 0 1480 0 -1 170
box -8 -3 16 105
use FILL  FILL_1570
timestamp 1710899220
transform 1 0 1472 0 -1 170
box -8 -3 16 105
use FILL  FILL_1571
timestamp 1710899220
transform 1 0 1464 0 -1 170
box -8 -3 16 105
use FILL  FILL_1572
timestamp 1710899220
transform 1 0 1456 0 -1 170
box -8 -3 16 105
use FILL  FILL_1573
timestamp 1710899220
transform 1 0 1448 0 -1 170
box -8 -3 16 105
use FILL  FILL_1574
timestamp 1710899220
transform 1 0 1248 0 -1 170
box -8 -3 16 105
use FILL  FILL_1575
timestamp 1710899220
transform 1 0 1240 0 -1 170
box -8 -3 16 105
use FILL  FILL_1576
timestamp 1710899220
transform 1 0 848 0 -1 170
box -8 -3 16 105
use FILL  FILL_1577
timestamp 1710899220
transform 1 0 648 0 -1 170
box -8 -3 16 105
use FILL  FILL_1578
timestamp 1710899220
transform 1 0 544 0 -1 170
box -8 -3 16 105
use FILL  FILL_1579
timestamp 1710899220
transform 1 0 536 0 -1 170
box -8 -3 16 105
use FILL  FILL_1580
timestamp 1710899220
transform 1 0 432 0 -1 170
box -8 -3 16 105
use FILL  FILL_1581
timestamp 1710899220
transform 1 0 424 0 -1 170
box -8 -3 16 105
use FILL  FILL_1582
timestamp 1710899220
transform 1 0 416 0 -1 170
box -8 -3 16 105
use FILL  FILL_1583
timestamp 1710899220
transform 1 0 408 0 -1 170
box -8 -3 16 105
use FILL  FILL_1584
timestamp 1710899220
transform 1 0 400 0 -1 170
box -8 -3 16 105
use FILL  FILL_1585
timestamp 1710899220
transform 1 0 392 0 -1 170
box -8 -3 16 105
use FILL  FILL_1586
timestamp 1710899220
transform 1 0 384 0 -1 170
box -8 -3 16 105
use FILL  FILL_1587
timestamp 1710899220
transform 1 0 376 0 -1 170
box -8 -3 16 105
use FILL  FILL_1588
timestamp 1710899220
transform 1 0 368 0 -1 170
box -8 -3 16 105
use FILL  FILL_1589
timestamp 1710899220
transform 1 0 360 0 -1 170
box -8 -3 16 105
use FILL  FILL_1590
timestamp 1710899220
transform 1 0 352 0 -1 170
box -8 -3 16 105
use FILL  FILL_1591
timestamp 1710899220
transform 1 0 344 0 -1 170
box -8 -3 16 105
use FILL  FILL_1592
timestamp 1710899220
transform 1 0 336 0 -1 170
box -8 -3 16 105
use FILL  FILL_1593
timestamp 1710899220
transform 1 0 328 0 -1 170
box -8 -3 16 105
use FILL  FILL_1594
timestamp 1710899220
transform 1 0 320 0 -1 170
box -8 -3 16 105
use FILL  FILL_1595
timestamp 1710899220
transform 1 0 312 0 -1 170
box -8 -3 16 105
use FILL  FILL_1596
timestamp 1710899220
transform 1 0 304 0 -1 170
box -8 -3 16 105
use FILL  FILL_1597
timestamp 1710899220
transform 1 0 296 0 -1 170
box -8 -3 16 105
use FILL  FILL_1598
timestamp 1710899220
transform 1 0 288 0 -1 170
box -8 -3 16 105
use FILL  FILL_1599
timestamp 1710899220
transform 1 0 280 0 -1 170
box -8 -3 16 105
use FILL  FILL_1600
timestamp 1710899220
transform 1 0 272 0 -1 170
box -8 -3 16 105
use FILL  FILL_1601
timestamp 1710899220
transform 1 0 264 0 -1 170
box -8 -3 16 105
use FILL  FILL_1602
timestamp 1710899220
transform 1 0 256 0 -1 170
box -8 -3 16 105
use FILL  FILL_1603
timestamp 1710899220
transform 1 0 248 0 -1 170
box -8 -3 16 105
use FILL  FILL_1604
timestamp 1710899220
transform 1 0 240 0 -1 170
box -8 -3 16 105
use FILL  FILL_1605
timestamp 1710899220
transform 1 0 232 0 -1 170
box -8 -3 16 105
use FILL  FILL_1606
timestamp 1710899220
transform 1 0 224 0 -1 170
box -8 -3 16 105
use FILL  FILL_1607
timestamp 1710899220
transform 1 0 216 0 -1 170
box -8 -3 16 105
use FILL  FILL_1608
timestamp 1710899220
transform 1 0 208 0 -1 170
box -8 -3 16 105
use FILL  FILL_1609
timestamp 1710899220
transform 1 0 200 0 -1 170
box -8 -3 16 105
use FILL  FILL_1610
timestamp 1710899220
transform 1 0 192 0 -1 170
box -8 -3 16 105
use FILL  FILL_1611
timestamp 1710899220
transform 1 0 184 0 -1 170
box -8 -3 16 105
use FILL  FILL_1612
timestamp 1710899220
transform 1 0 176 0 -1 170
box -8 -3 16 105
use FILL  FILL_1613
timestamp 1710899220
transform 1 0 168 0 -1 170
box -8 -3 16 105
use FILL  FILL_1614
timestamp 1710899220
transform 1 0 160 0 -1 170
box -8 -3 16 105
use FILL  FILL_1615
timestamp 1710899220
transform 1 0 152 0 -1 170
box -8 -3 16 105
use FILL  FILL_1616
timestamp 1710899220
transform 1 0 144 0 -1 170
box -8 -3 16 105
use FILL  FILL_1617
timestamp 1710899220
transform 1 0 136 0 -1 170
box -8 -3 16 105
use FILL  FILL_1618
timestamp 1710899220
transform 1 0 128 0 -1 170
box -8 -3 16 105
use FILL  FILL_1619
timestamp 1710899220
transform 1 0 120 0 -1 170
box -8 -3 16 105
use FILL  FILL_1620
timestamp 1710899220
transform 1 0 112 0 -1 170
box -8 -3 16 105
use FILL  FILL_1621
timestamp 1710899220
transform 1 0 104 0 -1 170
box -8 -3 16 105
use FILL  FILL_1622
timestamp 1710899220
transform 1 0 96 0 -1 170
box -8 -3 16 105
use FILL  FILL_1623
timestamp 1710899220
transform 1 0 88 0 -1 170
box -8 -3 16 105
use FILL  FILL_1624
timestamp 1710899220
transform 1 0 80 0 -1 170
box -8 -3 16 105
use FILL  FILL_1625
timestamp 1710899220
transform 1 0 72 0 -1 170
box -8 -3 16 105
use HAX1  HAX1_0
timestamp 1710899220
transform 1 0 2496 0 1 1170
box -5 -3 84 105
use HAX1  HAX1_1
timestamp 1710899220
transform 1 0 2376 0 1 1170
box -5 -3 84 105
use HAX1  HAX1_2
timestamp 1710899220
transform 1 0 2368 0 -1 1370
box -5 -3 84 105
use HAX1  HAX1_3
timestamp 1710899220
transform 1 0 2344 0 -1 1570
box -5 -3 84 105
use HAX1  HAX1_4
timestamp 1710899220
transform 1 0 2424 0 -1 1570
box -5 -3 84 105
use HAX1  HAX1_5
timestamp 1710899220
transform 1 0 2544 0 -1 1570
box -5 -3 84 105
use HAX1  HAX1_6
timestamp 1710899220
transform 1 0 2456 0 -1 1770
box -5 -3 84 105
use HAX1  HAX1_7
timestamp 1710899220
transform 1 0 2376 0 -1 1770
box -5 -3 84 105
use HAX1  HAX1_8
timestamp 1710899220
transform 1 0 2376 0 1 1770
box -5 -3 84 105
use HAX1  HAX1_9
timestamp 1710899220
transform 1 0 2456 0 1 1770
box -5 -3 84 105
use HAX1  HAX1_10
timestamp 1710899220
transform 1 0 2424 0 -1 1970
box -5 -3 84 105
use HAX1  HAX1_11
timestamp 1710899220
transform 1 0 2440 0 1 1970
box -5 -3 84 105
use HAX1  HAX1_12
timestamp 1710899220
transform 1 0 2440 0 1 2170
box -5 -3 84 105
use HAX1  HAX1_13
timestamp 1710899220
transform 1 0 2360 0 1 2170
box -5 -3 84 105
use HAX1  HAX1_14
timestamp 1710899220
transform 1 0 2440 0 -1 2370
box -5 -3 84 105
use HAX1  HAX1_15
timestamp 1710899220
transform 1 0 2480 0 1 2370
box -5 -3 84 105
use HAX1  HAX1_16
timestamp 1710899220
transform 1 0 2400 0 1 2370
box -5 -3 84 105
use HAX1  HAX1_17
timestamp 1710899220
transform 1 0 2200 0 1 2370
box -5 -3 84 105
use HAX1  HAX1_18
timestamp 1710899220
transform 1 0 2152 0 -1 2370
box -5 -3 84 105
use HAX1  HAX1_19
timestamp 1710899220
transform 1 0 2064 0 -1 2370
box -5 -3 84 105
use HAX1  HAX1_20
timestamp 1710899220
transform 1 0 2064 0 -1 2570
box -5 -3 84 105
use HAX1  HAX1_21
timestamp 1710899220
transform 1 0 1984 0 -1 2570
box -5 -3 84 105
use HAX1  HAX1_22
timestamp 1710899220
transform 1 0 1968 0 1 2370
box -5 -3 84 105
use HAX1  HAX1_23
timestamp 1710899220
transform 1 0 1968 0 1 2170
box -5 -3 84 105
use HAX1  HAX1_24
timestamp 1710899220
transform 1 0 1936 0 -1 2170
box -5 -3 84 105
use HAX1  HAX1_25
timestamp 1710899220
transform 1 0 1968 0 1 1970
box -5 -3 84 105
use HAX1  HAX1_26
timestamp 1710899220
transform 1 0 2080 0 1 1970
box -5 -3 84 105
use HAX1  HAX1_27
timestamp 1710899220
transform 1 0 2168 0 1 1970
box -5 -3 84 105
use HAX1  HAX1_28
timestamp 1710899220
transform 1 0 2176 0 -1 2170
box -5 -3 84 105
use HAX1  HAX1_29
timestamp 1710899220
transform 1 0 2272 0 -1 2170
box -5 -3 84 105
use HAX1  HAX1_30
timestamp 1710899220
transform 1 0 1120 0 -1 2170
box -5 -3 84 105
use HAX1  HAX1_31
timestamp 1710899220
transform 1 0 424 0 1 1970
box -5 -3 84 105
use HAX1  HAX1_32
timestamp 1710899220
transform 1 0 744 0 1 1970
box -5 -3 84 105
use HAX1  HAX1_33
timestamp 1710899220
transform 1 0 648 0 1 2170
box -5 -3 84 105
use HAX1  HAX1_34
timestamp 1710899220
transform 1 0 1056 0 1 1970
box -5 -3 84 105
use HAX1  HAX1_35
timestamp 1710899220
transform 1 0 2120 0 -1 1570
box -5 -3 84 105
use HAX1  HAX1_36
timestamp 1710899220
transform 1 0 2112 0 -1 1770
box -5 -3 84 105
use HAX1  HAX1_37
timestamp 1710899220
transform 1 0 2032 0 -1 1770
box -5 -3 84 105
use HAX1  HAX1_38
timestamp 1710899220
transform 1 0 392 0 -1 2570
box -5 -3 84 105
use HAX1  HAX1_39
timestamp 1710899220
transform 1 0 264 0 -1 2570
box -5 -3 84 105
use HAX1  HAX1_40
timestamp 1710899220
transform 1 0 696 0 -1 2570
box -5 -3 84 105
use HAX1  HAX1_41
timestamp 1710899220
transform 1 0 568 0 -1 2570
box -5 -3 84 105
use HAX1  HAX1_42
timestamp 1710899220
transform 1 0 1016 0 -1 2570
box -5 -3 84 105
use HAX1  HAX1_43
timestamp 1710899220
transform 1 0 888 0 -1 2570
box -5 -3 84 105
use HAX1  HAX1_44
timestamp 1710899220
transform 1 0 1496 0 -1 2570
box -5 -3 84 105
use HAX1  HAX1_45
timestamp 1710899220
transform 1 0 1368 0 -1 2570
box -5 -3 84 105
use HAX1  HAX1_46
timestamp 1710899220
transform 1 0 1592 0 1 2370
box -5 -3 84 105
use HAX1  HAX1_47
timestamp 1710899220
transform 1 0 1688 0 -1 2570
box -5 -3 84 105
use HAX1  HAX1_48
timestamp 1710899220
transform 1 0 1720 0 1 2170
box -5 -3 84 105
use HAX1  HAX1_49
timestamp 1710899220
transform 1 0 1752 0 -1 2370
box -5 -3 84 105
use INVX1  INVX1_0
timestamp 1710899220
transform 1 0 2264 0 1 970
box -9 -3 26 105
use INVX2  INVX2_0
timestamp 1710899220
transform 1 0 2080 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_1
timestamp 1710899220
transform 1 0 1376 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_2
timestamp 1710899220
transform 1 0 1504 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_3
timestamp 1710899220
transform 1 0 1152 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_4
timestamp 1710899220
transform 1 0 1008 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_5
timestamp 1710899220
transform 1 0 1920 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_6
timestamp 1710899220
transform 1 0 1528 0 1 970
box -9 -3 26 105
use INVX2  INVX2_7
timestamp 1710899220
transform 1 0 1888 0 1 370
box -9 -3 26 105
use INVX2  INVX2_8
timestamp 1710899220
transform 1 0 1536 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_9
timestamp 1710899220
transform 1 0 1824 0 1 770
box -9 -3 26 105
use INVX2  INVX2_10
timestamp 1710899220
transform 1 0 1784 0 1 970
box -9 -3 26 105
use INVX2  INVX2_11
timestamp 1710899220
transform 1 0 448 0 1 170
box -9 -3 26 105
use INVX2  INVX2_12
timestamp 1710899220
transform 1 0 968 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_13
timestamp 1710899220
transform 1 0 944 0 1 370
box -9 -3 26 105
use INVX2  INVX2_14
timestamp 1710899220
transform 1 0 984 0 1 770
box -9 -3 26 105
use INVX2  INVX2_15
timestamp 1710899220
transform 1 0 1600 0 1 770
box -9 -3 26 105
use INVX2  INVX2_16
timestamp 1710899220
transform 1 0 840 0 1 770
box -9 -3 26 105
use INVX2  INVX2_17
timestamp 1710899220
transform 1 0 1136 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_18
timestamp 1710899220
transform 1 0 560 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_19
timestamp 1710899220
transform 1 0 464 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_20
timestamp 1710899220
transform 1 0 672 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_21
timestamp 1710899220
transform 1 0 968 0 1 770
box -9 -3 26 105
use INVX2  INVX2_22
timestamp 1710899220
transform 1 0 528 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_23
timestamp 1710899220
transform 1 0 760 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_24
timestamp 1710899220
transform 1 0 824 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_25
timestamp 1710899220
transform 1 0 808 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_26
timestamp 1710899220
transform 1 0 1184 0 1 370
box -9 -3 26 105
use INVX2  INVX2_27
timestamp 1710899220
transform 1 0 1552 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_28
timestamp 1710899220
transform 1 0 1664 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_29
timestamp 1710899220
transform 1 0 2016 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_30
timestamp 1710899220
transform 1 0 1168 0 1 770
box -9 -3 26 105
use INVX2  INVX2_31
timestamp 1710899220
transform 1 0 952 0 1 770
box -9 -3 26 105
use INVX2  INVX2_32
timestamp 1710899220
transform 1 0 984 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_33
timestamp 1710899220
transform 1 0 944 0 1 970
box -9 -3 26 105
use INVX2  INVX2_34
timestamp 1710899220
transform 1 0 264 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_35
timestamp 1710899220
transform 1 0 264 0 1 770
box -9 -3 26 105
use INVX2  INVX2_36
timestamp 1710899220
transform 1 0 160 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_37
timestamp 1710899220
transform 1 0 424 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_38
timestamp 1710899220
transform 1 0 256 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_39
timestamp 1710899220
transform 1 0 184 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_40
timestamp 1710899220
transform 1 0 1232 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_41
timestamp 1710899220
transform 1 0 880 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_42
timestamp 1710899220
transform 1 0 888 0 1 970
box -9 -3 26 105
use INVX2  INVX2_43
timestamp 1710899220
transform 1 0 1040 0 1 970
box -9 -3 26 105
use INVX2  INVX2_44
timestamp 1710899220
transform 1 0 1664 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_45
timestamp 1710899220
transform 1 0 1392 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_46
timestamp 1710899220
transform 1 0 1032 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_47
timestamp 1710899220
transform 1 0 1016 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_48
timestamp 1710899220
transform 1 0 1576 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_49
timestamp 1710899220
transform 1 0 1616 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_50
timestamp 1710899220
transform 1 0 1168 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_51
timestamp 1710899220
transform 1 0 816 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_52
timestamp 1710899220
transform 1 0 712 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_53
timestamp 1710899220
transform 1 0 552 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_54
timestamp 1710899220
transform 1 0 720 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_55
timestamp 1710899220
transform 1 0 720 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_56
timestamp 1710899220
transform 1 0 584 0 1 370
box -9 -3 26 105
use INVX2  INVX2_57
timestamp 1710899220
transform 1 0 416 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_58
timestamp 1710899220
transform 1 0 1688 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_59
timestamp 1710899220
transform 1 0 472 0 1 570
box -9 -3 26 105
use INVX2  INVX2_60
timestamp 1710899220
transform 1 0 1136 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_61
timestamp 1710899220
transform 1 0 944 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_62
timestamp 1710899220
transform 1 0 1592 0 1 570
box -9 -3 26 105
use INVX2  INVX2_63
timestamp 1710899220
transform 1 0 832 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_64
timestamp 1710899220
transform 1 0 592 0 1 170
box -9 -3 26 105
use INVX2  INVX2_65
timestamp 1710899220
transform 1 0 680 0 1 170
box -9 -3 26 105
use INVX2  INVX2_66
timestamp 1710899220
transform 1 0 776 0 1 170
box -9 -3 26 105
use INVX2  INVX2_67
timestamp 1710899220
transform 1 0 920 0 1 170
box -9 -3 26 105
use INVX2  INVX2_68
timestamp 1710899220
transform 1 0 1128 0 1 170
box -9 -3 26 105
use INVX2  INVX2_69
timestamp 1710899220
transform 1 0 1224 0 1 170
box -9 -3 26 105
use INVX2  INVX2_70
timestamp 1710899220
transform 1 0 1552 0 1 170
box -9 -3 26 105
use INVX2  INVX2_71
timestamp 1710899220
transform 1 0 1608 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_72
timestamp 1710899220
transform 1 0 1392 0 1 170
box -9 -3 26 105
use INVX2  INVX2_73
timestamp 1710899220
transform 1 0 1672 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_74
timestamp 1710899220
transform 1 0 1792 0 1 170
box -9 -3 26 105
use INVX2  INVX2_75
timestamp 1710899220
transform 1 0 1936 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_76
timestamp 1710899220
transform 1 0 1824 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_77
timestamp 1710899220
transform 1 0 1832 0 1 370
box -9 -3 26 105
use INVX2  INVX2_78
timestamp 1710899220
transform 1 0 1544 0 1 770
box -9 -3 26 105
use INVX2  INVX2_79
timestamp 1710899220
transform 1 0 1448 0 1 770
box -9 -3 26 105
use INVX2  INVX2_80
timestamp 1710899220
transform 1 0 1664 0 1 770
box -9 -3 26 105
use INVX2  INVX2_81
timestamp 1710899220
transform 1 0 1616 0 1 770
box -9 -3 26 105
use INVX2  INVX2_82
timestamp 1710899220
transform 1 0 1816 0 1 570
box -9 -3 26 105
use INVX2  INVX2_83
timestamp 1710899220
transform 1 0 1944 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_84
timestamp 1710899220
transform 1 0 1736 0 1 770
box -9 -3 26 105
use INVX2  INVX2_85
timestamp 1710899220
transform 1 0 1552 0 1 570
box -9 -3 26 105
use INVX2  INVX2_86
timestamp 1710899220
transform 1 0 1544 0 1 970
box -9 -3 26 105
use INVX2  INVX2_87
timestamp 1710899220
transform 1 0 1480 0 1 970
box -9 -3 26 105
use INVX2  INVX2_88
timestamp 1710899220
transform 1 0 1728 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_89
timestamp 1710899220
transform 1 0 688 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_90
timestamp 1710899220
transform 1 0 376 0 1 370
box -9 -3 26 105
use INVX2  INVX2_91
timestamp 1710899220
transform 1 0 344 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_92
timestamp 1710899220
transform 1 0 312 0 1 570
box -9 -3 26 105
use INVX2  INVX2_93
timestamp 1710899220
transform 1 0 1120 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_94
timestamp 1710899220
transform 1 0 1008 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_95
timestamp 1710899220
transform 1 0 840 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_96
timestamp 1710899220
transform 1 0 488 0 1 170
box -9 -3 26 105
use INVX2  INVX2_97
timestamp 1710899220
transform 1 0 336 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_98
timestamp 1710899220
transform 1 0 328 0 1 170
box -9 -3 26 105
use INVX2  INVX2_99
timestamp 1710899220
transform 1 0 1008 0 1 170
box -9 -3 26 105
use INVX2  INVX2_100
timestamp 1710899220
transform 1 0 1072 0 1 170
box -9 -3 26 105
use INVX2  INVX2_101
timestamp 1710899220
transform 1 0 1184 0 1 170
box -9 -3 26 105
use INVX2  INVX2_102
timestamp 1710899220
transform 1 0 1696 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_103
timestamp 1710899220
transform 1 0 1616 0 1 170
box -9 -3 26 105
use INVX2  INVX2_104
timestamp 1710899220
transform 1 0 1696 0 1 170
box -9 -3 26 105
use INVX2  INVX2_105
timestamp 1710899220
transform 1 0 2024 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_106
timestamp 1710899220
transform 1 0 2016 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_107
timestamp 1710899220
transform 1 0 1992 0 1 170
box -9 -3 26 105
use INVX2  INVX2_108
timestamp 1710899220
transform 1 0 1552 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_109
timestamp 1710899220
transform 1 0 1760 0 1 970
box -9 -3 26 105
use INVX2  INVX2_110
timestamp 1710899220
transform 1 0 1888 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_111
timestamp 1710899220
transform 1 0 1992 0 1 570
box -9 -3 26 105
use INVX2  INVX2_112
timestamp 1710899220
transform 1 0 2000 0 1 770
box -9 -3 26 105
use INVX2  INVX2_113
timestamp 1710899220
transform 1 0 2040 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_114
timestamp 1710899220
transform 1 0 2304 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_115
timestamp 1710899220
transform 1 0 2248 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_116
timestamp 1710899220
transform 1 0 2552 0 1 770
box -9 -3 26 105
use INVX2  INVX2_117
timestamp 1710899220
transform 1 0 2504 0 1 370
box -9 -3 26 105
use INVX2  INVX2_118
timestamp 1710899220
transform 1 0 2496 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_119
timestamp 1710899220
transform 1 0 2472 0 1 170
box -9 -3 26 105
use INVX2  INVX2_120
timestamp 1710899220
transform 1 0 2520 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_121
timestamp 1710899220
transform 1 0 2560 0 1 170
box -9 -3 26 105
use INVX2  INVX2_122
timestamp 1710899220
transform 1 0 2440 0 1 770
box -9 -3 26 105
use INVX2  INVX2_123
timestamp 1710899220
transform 1 0 2536 0 1 770
box -9 -3 26 105
use INVX2  INVX2_124
timestamp 1710899220
transform 1 0 2384 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_125
timestamp 1710899220
transform 1 0 2624 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_126
timestamp 1710899220
transform 1 0 2624 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_127
timestamp 1710899220
transform 1 0 2456 0 1 170
box -9 -3 26 105
use INVX2  INVX2_128
timestamp 1710899220
transform 1 0 2440 0 1 170
box -9 -3 26 105
use INVX2  INVX2_129
timestamp 1710899220
transform 1 0 2128 0 1 770
box -9 -3 26 105
use INVX2  INVX2_130
timestamp 1710899220
transform 1 0 2248 0 1 970
box -9 -3 26 105
use INVX2  INVX2_131
timestamp 1710899220
transform 1 0 2176 0 1 570
box -9 -3 26 105
use INVX2  INVX2_132
timestamp 1710899220
transform 1 0 2160 0 1 570
box -9 -3 26 105
use INVX2  INVX2_133
timestamp 1710899220
transform 1 0 2480 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_134
timestamp 1710899220
transform 1 0 1232 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_135
timestamp 1710899220
transform 1 0 1432 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_136
timestamp 1710899220
transform 1 0 1184 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_137
timestamp 1710899220
transform 1 0 1512 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_138
timestamp 1710899220
transform 1 0 928 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_139
timestamp 1710899220
transform 1 0 1440 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_140
timestamp 1710899220
transform 1 0 272 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_141
timestamp 1710899220
transform 1 0 1256 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_142
timestamp 1710899220
transform 1 0 256 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_143
timestamp 1710899220
transform 1 0 992 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_144
timestamp 1710899220
transform 1 0 696 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_145
timestamp 1710899220
transform 1 0 424 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_146
timestamp 1710899220
transform 1 0 216 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_147
timestamp 1710899220
transform 1 0 216 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_148
timestamp 1710899220
transform 1 0 248 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_149
timestamp 1710899220
transform 1 0 272 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_150
timestamp 1710899220
transform 1 0 512 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_151
timestamp 1710899220
transform 1 0 456 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_152
timestamp 1710899220
transform 1 0 496 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_153
timestamp 1710899220
transform 1 0 520 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_154
timestamp 1710899220
transform 1 0 744 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_155
timestamp 1710899220
transform 1 0 640 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_156
timestamp 1710899220
transform 1 0 760 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_157
timestamp 1710899220
transform 1 0 824 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_158
timestamp 1710899220
transform 1 0 840 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_159
timestamp 1710899220
transform 1 0 1224 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_160
timestamp 1710899220
transform 1 0 1040 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_161
timestamp 1710899220
transform 1 0 832 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_162
timestamp 1710899220
transform 1 0 1288 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_163
timestamp 1710899220
transform 1 0 1304 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_164
timestamp 1710899220
transform 1 0 1320 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_165
timestamp 1710899220
transform 1 0 1472 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_166
timestamp 1710899220
transform 1 0 1296 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_167
timestamp 1710899220
transform 1 0 1624 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_168
timestamp 1710899220
transform 1 0 1640 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_169
timestamp 1710899220
transform 1 0 1424 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_170
timestamp 1710899220
transform 1 0 1552 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_171
timestamp 1710899220
transform 1 0 1576 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_172
timestamp 1710899220
transform 1 0 1816 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_173
timestamp 1710899220
transform 1 0 1728 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_174
timestamp 1710899220
transform 1 0 1648 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_175
timestamp 1710899220
transform 1 0 1528 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_176
timestamp 1710899220
transform 1 0 1632 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_177
timestamp 1710899220
transform 1 0 1440 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_178
timestamp 1710899220
transform 1 0 1456 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_179
timestamp 1710899220
transform 1 0 1528 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_180
timestamp 1710899220
transform 1 0 1264 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_181
timestamp 1710899220
transform 1 0 1360 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_182
timestamp 1710899220
transform 1 0 1600 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_183
timestamp 1710899220
transform 1 0 1496 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_184
timestamp 1710899220
transform 1 0 2168 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_185
timestamp 1710899220
transform 1 0 2656 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_186
timestamp 1710899220
transform 1 0 2544 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_187
timestamp 1710899220
transform 1 0 2448 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_188
timestamp 1710899220
transform 1 0 2296 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_189
timestamp 1710899220
transform 1 0 2328 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_190
timestamp 1710899220
transform 1 0 2504 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_191
timestamp 1710899220
transform 1 0 2624 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_192
timestamp 1710899220
transform 1 0 2608 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_193
timestamp 1710899220
transform 1 0 2320 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_194
timestamp 1710899220
transform 1 0 2320 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_195
timestamp 1710899220
transform 1 0 2656 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_196
timestamp 1710899220
transform 1 0 2544 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_197
timestamp 1710899220
transform 1 0 2560 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_198
timestamp 1710899220
transform 1 0 2656 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_199
timestamp 1710899220
transform 1 0 2384 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_200
timestamp 1710899220
transform 1 0 2560 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_201
timestamp 1710899220
transform 1 0 2600 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_202
timestamp 1710899220
transform 1 0 2392 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_203
timestamp 1710899220
transform 1 0 2320 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_204
timestamp 1710899220
transform 1 0 2288 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_205
timestamp 1710899220
transform 1 0 2040 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_206
timestamp 1710899220
transform 1 0 2184 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_207
timestamp 1710899220
transform 1 0 1928 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_208
timestamp 1710899220
transform 1 0 1912 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_209
timestamp 1710899220
transform 1 0 1912 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_210
timestamp 1710899220
transform 1 0 1872 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_211
timestamp 1710899220
transform 1 0 1912 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_212
timestamp 1710899220
transform 1 0 2088 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_213
timestamp 1710899220
transform 1 0 2200 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_214
timestamp 1710899220
transform 1 0 2120 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_215
timestamp 1710899220
transform 1 0 2312 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_216
timestamp 1710899220
transform 1 0 2248 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_217
timestamp 1710899220
transform 1 0 1768 0 1 770
box -9 -3 26 105
use INVX2  INVX2_218
timestamp 1710899220
transform 1 0 2040 0 1 970
box -9 -3 26 105
use INVX2  INVX2_219
timestamp 1710899220
transform 1 0 2264 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_220
timestamp 1710899220
transform 1 0 1168 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_221
timestamp 1710899220
transform 1 0 1088 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_222
timestamp 1710899220
transform 1 0 1680 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_223
timestamp 1710899220
transform 1 0 1040 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_224
timestamp 1710899220
transform 1 0 848 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_225
timestamp 1710899220
transform 1 0 1408 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_226
timestamp 1710899220
transform 1 0 1712 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_227
timestamp 1710899220
transform 1 0 704 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_228
timestamp 1710899220
transform 1 0 1072 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_229
timestamp 1710899220
transform 1 0 1176 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_230
timestamp 1710899220
transform 1 0 1160 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_231
timestamp 1710899220
transform 1 0 1784 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_232
timestamp 1710899220
transform 1 0 1680 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_233
timestamp 1710899220
transform 1 0 656 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_234
timestamp 1710899220
transform 1 0 1120 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_235
timestamp 1710899220
transform 1 0 1288 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_236
timestamp 1710899220
transform 1 0 1192 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_237
timestamp 1710899220
transform 1 0 1544 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_238
timestamp 1710899220
transform 1 0 1544 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_239
timestamp 1710899220
transform 1 0 1032 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_240
timestamp 1710899220
transform 1 0 1056 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_241
timestamp 1710899220
transform 1 0 1312 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_242
timestamp 1710899220
transform 1 0 1352 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_243
timestamp 1710899220
transform 1 0 1624 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_244
timestamp 1710899220
transform 1 0 1768 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_245
timestamp 1710899220
transform 1 0 1640 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_246
timestamp 1710899220
transform 1 0 128 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_247
timestamp 1710899220
transform 1 0 1072 0 1 770
box -9 -3 26 105
use INVX2  INVX2_248
timestamp 1710899220
transform 1 0 1888 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_249
timestamp 1710899220
transform 1 0 1912 0 1 970
box -9 -3 26 105
use INVX2  INVX2_250
timestamp 1710899220
transform 1 0 1928 0 1 970
box -9 -3 26 105
use INVX2  INVX2_251
timestamp 1710899220
transform 1 0 576 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_252
timestamp 1710899220
transform 1 0 672 0 1 970
box -9 -3 26 105
use INVX2  INVX2_253
timestamp 1710899220
transform 1 0 1872 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_254
timestamp 1710899220
transform 1 0 1088 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_255
timestamp 1710899220
transform 1 0 2040 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_256
timestamp 1710899220
transform 1 0 2056 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_257
timestamp 1710899220
transform 1 0 2264 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_258
timestamp 1710899220
transform 1 0 2248 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_259
timestamp 1710899220
transform 1 0 2280 0 1 970
box -9 -3 26 105
use M2_M1  M2_M1_0
timestamp 1710899220
transform 1 0 2300 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1
timestamp 1710899220
transform 1 0 2188 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2
timestamp 1710899220
transform 1 0 2204 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_3
timestamp 1710899220
transform 1 0 2180 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4
timestamp 1710899220
transform 1 0 2196 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5
timestamp 1710899220
transform 1 0 2092 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_6
timestamp 1710899220
transform 1 0 2108 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_7
timestamp 1710899220
transform 1 0 1980 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_8
timestamp 1710899220
transform 1 0 1996 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_9
timestamp 1710899220
transform 1 0 1948 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_10
timestamp 1710899220
transform 1 0 1972 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_11
timestamp 1710899220
transform 1 0 1972 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_12
timestamp 1710899220
transform 1 0 1996 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_13
timestamp 1710899220
transform 1 0 1980 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_14
timestamp 1710899220
transform 1 0 1996 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_15
timestamp 1710899220
transform 1 0 1996 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_16
timestamp 1710899220
transform 1 0 2060 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_17
timestamp 1710899220
transform 1 0 2020 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_18
timestamp 1710899220
transform 1 0 2092 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_19
timestamp 1710899220
transform 1 0 2076 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_20
timestamp 1710899220
transform 1 0 2140 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_21
timestamp 1710899220
transform 1 0 2100 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_22
timestamp 1710899220
transform 1 0 2188 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_23
timestamp 1710899220
transform 1 0 2188 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_24
timestamp 1710899220
transform 1 0 2412 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_25
timestamp 1710899220
transform 1 0 2236 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_26
timestamp 1710899220
transform 1 0 2476 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_27
timestamp 1710899220
transform 1 0 2428 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_28
timestamp 1710899220
transform 1 0 2508 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_29
timestamp 1710899220
transform 1 0 2452 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_30
timestamp 1710899220
transform 1 0 2468 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_31
timestamp 1710899220
transform 1 0 2372 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_32
timestamp 1710899220
transform 1 0 2444 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_33
timestamp 1710899220
transform 1 0 2396 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_34
timestamp 1710899220
transform 1 0 2476 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_35
timestamp 1710899220
transform 1 0 2452 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_36
timestamp 1710899220
transform 1 0 2468 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_37
timestamp 1710899220
transform 1 0 2436 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_38
timestamp 1710899220
transform 1 0 2460 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_39
timestamp 1710899220
transform 1 0 2460 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_40
timestamp 1710899220
transform 1 0 2484 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_41
timestamp 1710899220
transform 1 0 2388 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_42
timestamp 1710899220
transform 1 0 2412 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_43
timestamp 1710899220
transform 1 0 2388 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_44
timestamp 1710899220
transform 1 0 2452 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_45
timestamp 1710899220
transform 1 0 2412 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_46
timestamp 1710899220
transform 1 0 2556 0 1 1585
box -2 -2 2 2
use M2_M1  M2_M1_47
timestamp 1710899220
transform 1 0 2556 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_48
timestamp 1710899220
transform 1 0 2484 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_49
timestamp 1710899220
transform 1 0 2484 0 1 1585
box -2 -2 2 2
use M2_M1  M2_M1_50
timestamp 1710899220
transform 1 0 2572 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_51
timestamp 1710899220
transform 1 0 2436 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_52
timestamp 1710899220
transform 1 0 2452 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_53
timestamp 1710899220
transform 1 0 2356 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_54
timestamp 1710899220
transform 1 0 2380 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_55
timestamp 1710899220
transform 1 0 2372 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_56
timestamp 1710899220
transform 1 0 2396 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_57
timestamp 1710899220
transform 1 0 2388 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_58
timestamp 1710899220
transform 1 0 2500 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_59
timestamp 1710899220
transform 1 0 2412 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_60
timestamp 1710899220
transform 1 0 2620 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_61
timestamp 1710899220
transform 1 0 2532 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_62
timestamp 1710899220
transform 1 0 1348 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_63
timestamp 1710899220
transform 1 0 1164 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_64
timestamp 1710899220
transform 1 0 1260 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_65
timestamp 1710899220
transform 1 0 1012 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_66
timestamp 1710899220
transform 1 0 1108 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_67
timestamp 1710899220
transform 1 0 804 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_68
timestamp 1710899220
transform 1 0 900 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_69
timestamp 1710899220
transform 1 0 500 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_70
timestamp 1710899220
transform 1 0 492 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_71
timestamp 1710899220
transform 1 0 2108 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_72
timestamp 1710899220
transform 1 0 2068 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_73
timestamp 1710899220
transform 1 0 2140 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_74
timestamp 1710899220
transform 1 0 2132 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_75
timestamp 1710899220
transform 1 0 2156 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_76
timestamp 1710899220
transform 1 0 2068 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_77
timestamp 1710899220
transform 1 0 1732 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_78
timestamp 1710899220
transform 1 0 1652 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_79
timestamp 1710899220
transform 1 0 1652 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_80
timestamp 1710899220
transform 1 0 1604 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_81
timestamp 1710899220
transform 1 0 1524 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_82
timestamp 1710899220
transform 1 0 1388 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_83
timestamp 1710899220
transform 1 0 1764 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_84
timestamp 1710899220
transform 1 0 1684 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_85
timestamp 1710899220
transform 1 0 1668 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_86
timestamp 1710899220
transform 1 0 1596 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_87
timestamp 1710899220
transform 1 0 1572 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_88
timestamp 1710899220
transform 1 0 1548 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_89
timestamp 1710899220
transform 1 0 1468 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_90
timestamp 1710899220
transform 1 0 1572 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_91
timestamp 1710899220
transform 1 0 1492 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_92
timestamp 1710899220
transform 1 0 1444 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_93
timestamp 1710899220
transform 1 0 1380 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_94
timestamp 1710899220
transform 1 0 1364 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_95
timestamp 1710899220
transform 1 0 1340 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_96
timestamp 1710899220
transform 1 0 1244 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_97
timestamp 1710899220
transform 1 0 1196 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_98
timestamp 1710899220
transform 1 0 1156 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_99
timestamp 1710899220
transform 1 0 1092 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_100
timestamp 1710899220
transform 1 0 964 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_101
timestamp 1710899220
transform 1 0 892 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_102
timestamp 1710899220
transform 1 0 948 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_103
timestamp 1710899220
transform 1 0 892 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_104
timestamp 1710899220
transform 1 0 788 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_105
timestamp 1710899220
transform 1 0 772 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_106
timestamp 1710899220
transform 1 0 644 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_107
timestamp 1710899220
transform 1 0 564 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_108
timestamp 1710899220
transform 1 0 652 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_109
timestamp 1710899220
transform 1 0 572 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_110
timestamp 1710899220
transform 1 0 532 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_111
timestamp 1710899220
transform 1 0 468 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_112
timestamp 1710899220
transform 1 0 340 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_113
timestamp 1710899220
transform 1 0 260 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_114
timestamp 1710899220
transform 1 0 380 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_115
timestamp 1710899220
transform 1 0 300 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_116
timestamp 1710899220
transform 1 0 236 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_117
timestamp 1710899220
transform 1 0 180 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_118
timestamp 1710899220
transform 1 0 172 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_119
timestamp 1710899220
transform 1 0 164 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_120
timestamp 1710899220
transform 1 0 2516 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_121
timestamp 1710899220
transform 1 0 2492 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_122
timestamp 1710899220
transform 1 0 2460 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_123
timestamp 1710899220
transform 1 0 2380 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_124
timestamp 1710899220
transform 1 0 2356 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_125
timestamp 1710899220
transform 1 0 2276 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_126
timestamp 1710899220
transform 1 0 2612 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_127
timestamp 1710899220
transform 1 0 2540 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_128
timestamp 1710899220
transform 1 0 2524 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_129
timestamp 1710899220
transform 1 0 2452 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_130
timestamp 1710899220
transform 1 0 2428 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_131
timestamp 1710899220
transform 1 0 2636 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_132
timestamp 1710899220
transform 1 0 2612 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_133
timestamp 1710899220
transform 1 0 2476 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_134
timestamp 1710899220
transform 1 0 2476 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_135
timestamp 1710899220
transform 1 0 2476 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_136
timestamp 1710899220
transform 1 0 2460 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_137
timestamp 1710899220
transform 1 0 2436 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_138
timestamp 1710899220
transform 1 0 2572 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_139
timestamp 1710899220
transform 1 0 2572 0 1 455
box -2 -2 2 2
use M2_M1  M2_M1_140
timestamp 1710899220
transform 1 0 2524 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_141
timestamp 1710899220
transform 1 0 2524 0 1 455
box -2 -2 2 2
use M2_M1  M2_M1_142
timestamp 1710899220
transform 1 0 2516 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_143
timestamp 1710899220
transform 1 0 2508 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_144
timestamp 1710899220
transform 1 0 1724 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_145
timestamp 1710899220
transform 1 0 1596 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_146
timestamp 1710899220
transform 1 0 1540 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_147
timestamp 1710899220
transform 1 0 1452 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_148
timestamp 1710899220
transform 1 0 1420 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_149
timestamp 1710899220
transform 1 0 1364 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_150
timestamp 1710899220
transform 1 0 1220 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_151
timestamp 1710899220
transform 1 0 1148 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_152
timestamp 1710899220
transform 1 0 1068 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_153
timestamp 1710899220
transform 1 0 852 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_154
timestamp 1710899220
transform 1 0 756 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_155
timestamp 1710899220
transform 1 0 684 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_156
timestamp 1710899220
transform 1 0 492 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_157
timestamp 1710899220
transform 1 0 484 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_158
timestamp 1710899220
transform 1 0 404 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_159
timestamp 1710899220
transform 1 0 276 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_160
timestamp 1710899220
transform 1 0 196 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_161
timestamp 1710899220
transform 1 0 124 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_162
timestamp 1710899220
transform 1 0 148 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_163
timestamp 1710899220
transform 1 0 76 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_164
timestamp 1710899220
transform 1 0 76 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_165
timestamp 1710899220
transform 1 0 164 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_166
timestamp 1710899220
transform 1 0 156 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_167
timestamp 1710899220
transform 1 0 124 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_168
timestamp 1710899220
transform 1 0 268 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_169
timestamp 1710899220
transform 1 0 268 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_170
timestamp 1710899220
transform 1 0 516 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_171
timestamp 1710899220
transform 1 0 420 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_172
timestamp 1710899220
transform 1 0 396 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_173
timestamp 1710899220
transform 1 0 444 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_174
timestamp 1710899220
transform 1 0 420 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_175
timestamp 1710899220
transform 1 0 492 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_176
timestamp 1710899220
transform 1 0 388 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_177
timestamp 1710899220
transform 1 0 644 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_178
timestamp 1710899220
transform 1 0 588 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_179
timestamp 1710899220
transform 1 0 764 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_180
timestamp 1710899220
transform 1 0 700 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_181
timestamp 1710899220
transform 1 0 700 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_182
timestamp 1710899220
transform 1 0 628 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_183
timestamp 1710899220
transform 1 0 716 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_184
timestamp 1710899220
transform 1 0 692 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_185
timestamp 1710899220
transform 1 0 828 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_186
timestamp 1710899220
transform 1 0 692 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_187
timestamp 1710899220
transform 1 0 844 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_188
timestamp 1710899220
transform 1 0 820 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_189
timestamp 1710899220
transform 1 0 1228 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_190
timestamp 1710899220
transform 1 0 1172 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_191
timestamp 1710899220
transform 1 0 1164 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_192
timestamp 1710899220
transform 1 0 932 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_193
timestamp 1710899220
transform 1 0 1012 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_194
timestamp 1710899220
transform 1 0 988 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_195
timestamp 1710899220
transform 1 0 1292 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_196
timestamp 1710899220
transform 1 0 1012 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_197
timestamp 1710899220
transform 1 0 1308 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_198
timestamp 1710899220
transform 1 0 1140 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_199
timestamp 1710899220
transform 1 0 1324 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_200
timestamp 1710899220
transform 1 0 1284 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_201
timestamp 1710899220
transform 1 0 1444 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_202
timestamp 1710899220
transform 1 0 1444 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_203
timestamp 1710899220
transform 1 0 1372 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_204
timestamp 1710899220
transform 1 0 1204 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_205
timestamp 1710899220
transform 1 0 1276 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_206
timestamp 1710899220
transform 1 0 1252 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_207
timestamp 1710899220
transform 1 0 1628 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_208
timestamp 1710899220
transform 1 0 1492 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_209
timestamp 1710899220
transform 1 0 1644 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_210
timestamp 1710899220
transform 1 0 1620 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_211
timestamp 1710899220
transform 1 0 1564 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_212
timestamp 1710899220
transform 1 0 1564 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_213
timestamp 1710899220
transform 1 0 1460 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_214
timestamp 1710899220
transform 1 0 1388 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_215
timestamp 1710899220
transform 1 0 1428 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_216
timestamp 1710899220
transform 1 0 1428 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_217
timestamp 1710899220
transform 1 0 1636 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_218
timestamp 1710899220
transform 1 0 1636 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_219
timestamp 1710899220
transform 1 0 1748 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_220
timestamp 1710899220
transform 1 0 1668 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_221
timestamp 1710899220
transform 1 0 1644 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_222
timestamp 1710899220
transform 1 0 1628 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_223
timestamp 1710899220
transform 1 0 1532 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_224
timestamp 1710899220
transform 1 0 1508 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_225
timestamp 1710899220
transform 1 0 1708 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_226
timestamp 1710899220
transform 1 0 1436 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_227
timestamp 1710899220
transform 1 0 1396 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_228
timestamp 1710899220
transform 1 0 1348 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_229
timestamp 1710899220
transform 1 0 1332 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_230
timestamp 1710899220
transform 1 0 1684 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_231
timestamp 1710899220
transform 1 0 1460 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_232
timestamp 1710899220
transform 1 0 1420 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_233
timestamp 1710899220
transform 1 0 1364 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_234
timestamp 1710899220
transform 1 0 1356 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_235
timestamp 1710899220
transform 1 0 1652 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_236
timestamp 1710899220
transform 1 0 1636 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_237
timestamp 1710899220
transform 1 0 1564 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_238
timestamp 1710899220
transform 1 0 1548 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_239
timestamp 1710899220
transform 1 0 1540 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_240
timestamp 1710899220
transform 1 0 1588 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_241
timestamp 1710899220
transform 1 0 1572 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_242
timestamp 1710899220
transform 1 0 1556 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_243
timestamp 1710899220
transform 1 0 1548 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_244
timestamp 1710899220
transform 1 0 1540 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_245
timestamp 1710899220
transform 1 0 1524 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_246
timestamp 1710899220
transform 1 0 1516 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_247
timestamp 1710899220
transform 1 0 1500 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_248
timestamp 1710899220
transform 1 0 1436 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_249
timestamp 1710899220
transform 1 0 1420 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_250
timestamp 1710899220
transform 1 0 1356 0 1 1695
box -2 -2 2 2
use M2_M1  M2_M1_251
timestamp 1710899220
transform 1 0 1324 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_252
timestamp 1710899220
transform 1 0 804 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_253
timestamp 1710899220
transform 1 0 740 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_254
timestamp 1710899220
transform 1 0 732 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_255
timestamp 1710899220
transform 1 0 716 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_256
timestamp 1710899220
transform 1 0 660 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_257
timestamp 1710899220
transform 1 0 628 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_258
timestamp 1710899220
transform 1 0 596 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_259
timestamp 1710899220
transform 1 0 572 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_260
timestamp 1710899220
transform 1 0 548 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_261
timestamp 1710899220
transform 1 0 540 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_262
timestamp 1710899220
transform 1 0 532 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_263
timestamp 1710899220
transform 1 0 1196 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_264
timestamp 1710899220
transform 1 0 1172 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_265
timestamp 1710899220
transform 1 0 1148 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_266
timestamp 1710899220
transform 1 0 1124 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_267
timestamp 1710899220
transform 1 0 1332 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_268
timestamp 1710899220
transform 1 0 1332 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_269
timestamp 1710899220
transform 1 0 1324 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_270
timestamp 1710899220
transform 1 0 1220 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_271
timestamp 1710899220
transform 1 0 1092 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_272
timestamp 1710899220
transform 1 0 732 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_273
timestamp 1710899220
transform 1 0 716 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_274
timestamp 1710899220
transform 1 0 1356 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_275
timestamp 1710899220
transform 1 0 1316 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_276
timestamp 1710899220
transform 1 0 1308 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_277
timestamp 1710899220
transform 1 0 1292 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_278
timestamp 1710899220
transform 1 0 1348 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_279
timestamp 1710899220
transform 1 0 1340 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_280
timestamp 1710899220
transform 1 0 1324 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_281
timestamp 1710899220
transform 1 0 1292 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_282
timestamp 1710899220
transform 1 0 1284 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_283
timestamp 1710899220
transform 1 0 1340 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_284
timestamp 1710899220
transform 1 0 1332 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_285
timestamp 1710899220
transform 1 0 1324 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_286
timestamp 1710899220
transform 1 0 1100 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_287
timestamp 1710899220
transform 1 0 964 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_288
timestamp 1710899220
transform 1 0 764 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_289
timestamp 1710899220
transform 1 0 764 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_290
timestamp 1710899220
transform 1 0 1380 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_291
timestamp 1710899220
transform 1 0 1364 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_292
timestamp 1710899220
transform 1 0 1356 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_293
timestamp 1710899220
transform 1 0 1068 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_294
timestamp 1710899220
transform 1 0 884 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_295
timestamp 1710899220
transform 1 0 788 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_296
timestamp 1710899220
transform 1 0 788 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_297
timestamp 1710899220
transform 1 0 1380 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_298
timestamp 1710899220
transform 1 0 1348 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_299
timestamp 1710899220
transform 1 0 1348 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_300
timestamp 1710899220
transform 1 0 1340 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_301
timestamp 1710899220
transform 1 0 1308 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_302
timestamp 1710899220
transform 1 0 732 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_303
timestamp 1710899220
transform 1 0 724 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_304
timestamp 1710899220
transform 1 0 1100 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_305
timestamp 1710899220
transform 1 0 1060 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_306
timestamp 1710899220
transform 1 0 804 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_307
timestamp 1710899220
transform 1 0 780 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_308
timestamp 1710899220
transform 1 0 764 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_309
timestamp 1710899220
transform 1 0 1028 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_310
timestamp 1710899220
transform 1 0 980 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_311
timestamp 1710899220
transform 1 0 900 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_312
timestamp 1710899220
transform 1 0 732 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_313
timestamp 1710899220
transform 1 0 716 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_314
timestamp 1710899220
transform 1 0 1260 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_315
timestamp 1710899220
transform 1 0 1244 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_316
timestamp 1710899220
transform 1 0 1236 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_317
timestamp 1710899220
transform 1 0 804 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_318
timestamp 1710899220
transform 1 0 788 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_319
timestamp 1710899220
transform 1 0 2124 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_320
timestamp 1710899220
transform 1 0 2092 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_321
timestamp 1710899220
transform 1 0 1380 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_322
timestamp 1710899220
transform 1 0 1268 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_323
timestamp 1710899220
transform 1 0 1212 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_324
timestamp 1710899220
transform 1 0 1052 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_325
timestamp 1710899220
transform 1 0 724 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_326
timestamp 1710899220
transform 1 0 708 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_327
timestamp 1710899220
transform 1 0 1500 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_328
timestamp 1710899220
transform 1 0 1180 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_329
timestamp 1710899220
transform 1 0 1140 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_330
timestamp 1710899220
transform 1 0 692 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_331
timestamp 1710899220
transform 1 0 676 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_332
timestamp 1710899220
transform 1 0 660 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_333
timestamp 1710899220
transform 1 0 1156 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_334
timestamp 1710899220
transform 1 0 1052 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_335
timestamp 1710899220
transform 1 0 980 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_336
timestamp 1710899220
transform 1 0 828 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_337
timestamp 1710899220
transform 1 0 508 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_338
timestamp 1710899220
transform 1 0 460 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_339
timestamp 1710899220
transform 1 0 1012 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_340
timestamp 1710899220
transform 1 0 988 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_341
timestamp 1710899220
transform 1 0 852 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_342
timestamp 1710899220
transform 1 0 652 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_343
timestamp 1710899220
transform 1 0 428 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_344
timestamp 1710899220
transform 1 0 252 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_345
timestamp 1710899220
transform 1 0 1924 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_346
timestamp 1710899220
transform 1 0 1916 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_347
timestamp 1710899220
transform 1 0 1684 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_348
timestamp 1710899220
transform 1 0 1636 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_349
timestamp 1710899220
transform 1 0 1604 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_350
timestamp 1710899220
transform 1 0 1540 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_351
timestamp 1710899220
transform 1 0 2020 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_352
timestamp 1710899220
transform 1 0 1972 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_353
timestamp 1710899220
transform 1 0 1900 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_354
timestamp 1710899220
transform 1 0 1748 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_355
timestamp 1710899220
transform 1 0 1548 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_356
timestamp 1710899220
transform 1 0 1068 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_357
timestamp 1710899220
transform 1 0 1916 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_358
timestamp 1710899220
transform 1 0 1828 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_359
timestamp 1710899220
transform 1 0 1796 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_360
timestamp 1710899220
transform 1 0 1932 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_361
timestamp 1710899220
transform 1 0 1884 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_362
timestamp 1710899220
transform 1 0 1812 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_363
timestamp 1710899220
transform 1 0 1804 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_364
timestamp 1710899220
transform 1 0 444 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_365
timestamp 1710899220
transform 1 0 420 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_366
timestamp 1710899220
transform 1 0 404 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_367
timestamp 1710899220
transform 1 0 1012 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_368
timestamp 1710899220
transform 1 0 980 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_369
timestamp 1710899220
transform 1 0 1004 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_370
timestamp 1710899220
transform 1 0 932 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_371
timestamp 1710899220
transform 1 0 924 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_372
timestamp 1710899220
transform 1 0 1036 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_373
timestamp 1710899220
transform 1 0 988 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_374
timestamp 1710899220
transform 1 0 988 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_375
timestamp 1710899220
transform 1 0 972 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_376
timestamp 1710899220
transform 1 0 1948 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_377
timestamp 1710899220
transform 1 0 1884 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_378
timestamp 1710899220
transform 1 0 1844 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_379
timestamp 1710899220
transform 1 0 1620 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_380
timestamp 1710899220
transform 1 0 1652 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_381
timestamp 1710899220
transform 1 0 1620 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_382
timestamp 1710899220
transform 1 0 1476 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_383
timestamp 1710899220
transform 1 0 836 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_384
timestamp 1710899220
transform 1 0 780 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_385
timestamp 1710899220
transform 1 0 1148 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_386
timestamp 1710899220
transform 1 0 924 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_387
timestamp 1710899220
transform 1 0 876 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_388
timestamp 1710899220
transform 1 0 484 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_389
timestamp 1710899220
transform 1 0 276 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_390
timestamp 1710899220
transform 1 0 220 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_391
timestamp 1710899220
transform 1 0 732 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_392
timestamp 1710899220
transform 1 0 564 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_393
timestamp 1710899220
transform 1 0 524 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_394
timestamp 1710899220
transform 1 0 804 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_395
timestamp 1710899220
transform 1 0 732 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_396
timestamp 1710899220
transform 1 0 516 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_397
timestamp 1710899220
transform 1 0 348 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_398
timestamp 1710899220
transform 1 0 348 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_399
timestamp 1710899220
transform 1 0 724 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_400
timestamp 1710899220
transform 1 0 684 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_401
timestamp 1710899220
transform 1 0 1012 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_402
timestamp 1710899220
transform 1 0 1012 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_403
timestamp 1710899220
transform 1 0 980 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_404
timestamp 1710899220
transform 1 0 980 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_405
timestamp 1710899220
transform 1 0 940 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_406
timestamp 1710899220
transform 1 0 796 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_407
timestamp 1710899220
transform 1 0 748 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_408
timestamp 1710899220
transform 1 0 548 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_409
timestamp 1710899220
transform 1 0 540 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_410
timestamp 1710899220
transform 1 0 804 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_411
timestamp 1710899220
transform 1 0 772 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_412
timestamp 1710899220
transform 1 0 756 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_413
timestamp 1710899220
transform 1 0 740 0 1 1355
box -2 -2 2 2
use M2_M1  M2_M1_414
timestamp 1710899220
transform 1 0 740 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_415
timestamp 1710899220
transform 1 0 724 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_416
timestamp 1710899220
transform 1 0 508 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_417
timestamp 1710899220
transform 1 0 252 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_418
timestamp 1710899220
transform 1 0 204 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_419
timestamp 1710899220
transform 1 0 180 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_420
timestamp 1710899220
transform 1 0 836 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_421
timestamp 1710899220
transform 1 0 812 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_422
timestamp 1710899220
transform 1 0 788 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_423
timestamp 1710899220
transform 1 0 812 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_424
timestamp 1710899220
transform 1 0 764 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_425
timestamp 1710899220
transform 1 0 1636 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_426
timestamp 1710899220
transform 1 0 1180 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_427
timestamp 1710899220
transform 1 0 1132 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_428
timestamp 1710899220
transform 1 0 908 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_429
timestamp 1710899220
transform 1 0 1596 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_430
timestamp 1710899220
transform 1 0 1564 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_431
timestamp 1710899220
transform 1 0 1780 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_432
timestamp 1710899220
transform 1 0 1716 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_433
timestamp 1710899220
transform 1 0 1684 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_434
timestamp 1710899220
transform 1 0 2020 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_435
timestamp 1710899220
transform 1 0 1988 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_436
timestamp 1710899220
transform 1 0 1332 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_437
timestamp 1710899220
transform 1 0 1300 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_438
timestamp 1710899220
transform 1 0 1292 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_439
timestamp 1710899220
transform 1 0 1268 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_440
timestamp 1710899220
transform 1 0 1228 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_441
timestamp 1710899220
transform 1 0 1180 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_442
timestamp 1710899220
transform 1 0 1140 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_443
timestamp 1710899220
transform 1 0 1124 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_444
timestamp 1710899220
transform 1 0 1004 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_445
timestamp 1710899220
transform 1 0 964 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_446
timestamp 1710899220
transform 1 0 948 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_447
timestamp 1710899220
transform 1 0 932 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_448
timestamp 1710899220
transform 1 0 780 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_449
timestamp 1710899220
transform 1 0 732 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_450
timestamp 1710899220
transform 1 0 724 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_451
timestamp 1710899220
transform 1 0 724 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_452
timestamp 1710899220
transform 1 0 716 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_453
timestamp 1710899220
transform 1 0 996 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_454
timestamp 1710899220
transform 1 0 972 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_455
timestamp 1710899220
transform 1 0 900 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_456
timestamp 1710899220
transform 1 0 804 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_457
timestamp 1710899220
transform 1 0 692 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_458
timestamp 1710899220
transform 1 0 692 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_459
timestamp 1710899220
transform 1 0 692 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_460
timestamp 1710899220
transform 1 0 684 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_461
timestamp 1710899220
transform 1 0 1340 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_462
timestamp 1710899220
transform 1 0 1324 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_463
timestamp 1710899220
transform 1 0 1292 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_464
timestamp 1710899220
transform 1 0 1164 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_465
timestamp 1710899220
transform 1 0 1132 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_466
timestamp 1710899220
transform 1 0 1116 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_467
timestamp 1710899220
transform 1 0 1100 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_468
timestamp 1710899220
transform 1 0 1076 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_469
timestamp 1710899220
transform 1 0 1004 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_470
timestamp 1710899220
transform 1 0 1004 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_471
timestamp 1710899220
transform 1 0 932 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_472
timestamp 1710899220
transform 1 0 684 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_473
timestamp 1710899220
transform 1 0 644 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_474
timestamp 1710899220
transform 1 0 612 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_475
timestamp 1710899220
transform 1 0 604 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_476
timestamp 1710899220
transform 1 0 524 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_477
timestamp 1710899220
transform 1 0 524 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_478
timestamp 1710899220
transform 1 0 332 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_479
timestamp 1710899220
transform 1 0 332 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_480
timestamp 1710899220
transform 1 0 268 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_481
timestamp 1710899220
transform 1 0 236 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_482
timestamp 1710899220
transform 1 0 1140 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_483
timestamp 1710899220
transform 1 0 1100 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_484
timestamp 1710899220
transform 1 0 1092 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_485
timestamp 1710899220
transform 1 0 1084 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_486
timestamp 1710899220
transform 1 0 1044 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_487
timestamp 1710899220
transform 1 0 892 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_488
timestamp 1710899220
transform 1 0 788 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_489
timestamp 1710899220
transform 1 0 668 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_490
timestamp 1710899220
transform 1 0 668 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_491
timestamp 1710899220
transform 1 0 660 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_492
timestamp 1710899220
transform 1 0 636 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_493
timestamp 1710899220
transform 1 0 628 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_494
timestamp 1710899220
transform 1 0 340 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_495
timestamp 1710899220
transform 1 0 308 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_496
timestamp 1710899220
transform 1 0 308 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_497
timestamp 1710899220
transform 1 0 284 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_498
timestamp 1710899220
transform 1 0 244 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_499
timestamp 1710899220
transform 1 0 188 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_500
timestamp 1710899220
transform 1 0 172 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_501
timestamp 1710899220
transform 1 0 484 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_502
timestamp 1710899220
transform 1 0 468 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_503
timestamp 1710899220
transform 1 0 444 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_504
timestamp 1710899220
transform 1 0 308 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_505
timestamp 1710899220
transform 1 0 276 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_506
timestamp 1710899220
transform 1 0 260 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_507
timestamp 1710899220
transform 1 0 260 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_508
timestamp 1710899220
transform 1 0 252 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_509
timestamp 1710899220
transform 1 0 196 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_510
timestamp 1710899220
transform 1 0 148 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_511
timestamp 1710899220
transform 1 0 1244 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_512
timestamp 1710899220
transform 1 0 1244 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_513
timestamp 1710899220
transform 1 0 1196 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_514
timestamp 1710899220
transform 1 0 1180 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_515
timestamp 1710899220
transform 1 0 1020 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_516
timestamp 1710899220
transform 1 0 940 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_517
timestamp 1710899220
transform 1 0 900 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_518
timestamp 1710899220
transform 1 0 1100 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_519
timestamp 1710899220
transform 1 0 1068 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_520
timestamp 1710899220
transform 1 0 1684 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_521
timestamp 1710899220
transform 1 0 1684 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_522
timestamp 1710899220
transform 1 0 1396 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_523
timestamp 1710899220
transform 1 0 1364 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_524
timestamp 1710899220
transform 1 0 1076 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_525
timestamp 1710899220
transform 1 0 1052 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_526
timestamp 1710899220
transform 1 0 1052 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_527
timestamp 1710899220
transform 1 0 1036 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_528
timestamp 1710899220
transform 1 0 1724 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_529
timestamp 1710899220
transform 1 0 1676 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_530
timestamp 1710899220
transform 1 0 1644 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_531
timestamp 1710899220
transform 1 0 1596 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_532
timestamp 1710899220
transform 1 0 1348 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_533
timestamp 1710899220
transform 1 0 1228 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_534
timestamp 1710899220
transform 1 0 1196 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_535
timestamp 1710899220
transform 1 0 820 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_536
timestamp 1710899220
transform 1 0 788 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_537
timestamp 1710899220
transform 1 0 756 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_538
timestamp 1710899220
transform 1 0 732 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_539
timestamp 1710899220
transform 1 0 732 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_540
timestamp 1710899220
transform 1 0 596 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_541
timestamp 1710899220
transform 1 0 580 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_542
timestamp 1710899220
transform 1 0 1308 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_543
timestamp 1710899220
transform 1 0 1276 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_544
timestamp 1710899220
transform 1 0 1276 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_545
timestamp 1710899220
transform 1 0 1244 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_546
timestamp 1710899220
transform 1 0 1084 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_547
timestamp 1710899220
transform 1 0 732 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_548
timestamp 1710899220
transform 1 0 692 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_549
timestamp 1710899220
transform 1 0 716 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_550
timestamp 1710899220
transform 1 0 708 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_551
timestamp 1710899220
transform 1 0 668 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_552
timestamp 1710899220
transform 1 0 580 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_553
timestamp 1710899220
transform 1 0 556 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_554
timestamp 1710899220
transform 1 0 364 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_555
timestamp 1710899220
transform 1 0 548 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_556
timestamp 1710899220
transform 1 0 500 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_557
timestamp 1710899220
transform 1 0 396 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_558
timestamp 1710899220
transform 1 0 332 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_559
timestamp 1710899220
transform 1 0 1716 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_560
timestamp 1710899220
transform 1 0 1700 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_561
timestamp 1710899220
transform 1 0 556 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_562
timestamp 1710899220
transform 1 0 540 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_563
timestamp 1710899220
transform 1 0 492 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_564
timestamp 1710899220
transform 1 0 340 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_565
timestamp 1710899220
transform 1 0 300 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_566
timestamp 1710899220
transform 1 0 1148 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_567
timestamp 1710899220
transform 1 0 1148 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_568
timestamp 1710899220
transform 1 0 1084 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_569
timestamp 1710899220
transform 1 0 1020 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_570
timestamp 1710899220
transform 1 0 1044 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_571
timestamp 1710899220
transform 1 0 1020 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_572
timestamp 1710899220
transform 1 0 964 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_573
timestamp 1710899220
transform 1 0 844 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_574
timestamp 1710899220
transform 1 0 844 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_575
timestamp 1710899220
transform 1 0 828 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_576
timestamp 1710899220
transform 1 0 804 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_577
timestamp 1710899220
transform 1 0 756 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_578
timestamp 1710899220
transform 1 0 836 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_579
timestamp 1710899220
transform 1 0 756 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_580
timestamp 1710899220
transform 1 0 580 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_581
timestamp 1710899220
transform 1 0 556 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_582
timestamp 1710899220
transform 1 0 532 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_583
timestamp 1710899220
transform 1 0 836 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_584
timestamp 1710899220
transform 1 0 676 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_585
timestamp 1710899220
transform 1 0 652 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_586
timestamp 1710899220
transform 1 0 372 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_587
timestamp 1710899220
transform 1 0 324 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_588
timestamp 1710899220
transform 1 0 1388 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_589
timestamp 1710899220
transform 1 0 796 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_590
timestamp 1710899220
transform 1 0 396 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_591
timestamp 1710899220
transform 1 0 372 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_592
timestamp 1710899220
transform 1 0 1036 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_593
timestamp 1710899220
transform 1 0 1036 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_594
timestamp 1710899220
transform 1 0 996 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_595
timestamp 1710899220
transform 1 0 916 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_596
timestamp 1710899220
transform 1 0 892 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_597
timestamp 1710899220
transform 1 0 1276 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_598
timestamp 1710899220
transform 1 0 1164 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_599
timestamp 1710899220
transform 1 0 1132 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_600
timestamp 1710899220
transform 1 0 1116 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_601
timestamp 1710899220
transform 1 0 1300 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_602
timestamp 1710899220
transform 1 0 1268 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_603
timestamp 1710899220
transform 1 0 1204 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_604
timestamp 1710899220
transform 1 0 1172 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_605
timestamp 1710899220
transform 1 0 1684 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_606
timestamp 1710899220
transform 1 0 1636 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_607
timestamp 1710899220
transform 1 0 1564 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_608
timestamp 1710899220
transform 1 0 1412 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_609
timestamp 1710899220
transform 1 0 1284 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_610
timestamp 1710899220
transform 1 0 1620 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_611
timestamp 1710899220
transform 1 0 1604 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_612
timestamp 1710899220
transform 1 0 1484 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_613
timestamp 1710899220
transform 1 0 1380 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_614
timestamp 1710899220
transform 1 0 1684 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_615
timestamp 1710899220
transform 1 0 1660 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_616
timestamp 1710899220
transform 1 0 1452 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_617
timestamp 1710899220
transform 1 0 1388 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_618
timestamp 1710899220
transform 1 0 1364 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_619
timestamp 1710899220
transform 1 0 1708 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_620
timestamp 1710899220
transform 1 0 1692 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_621
timestamp 1710899220
transform 1 0 2012 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_622
timestamp 1710899220
transform 1 0 1964 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_623
timestamp 1710899220
transform 1 0 1844 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_624
timestamp 1710899220
transform 1 0 1804 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_625
timestamp 1710899220
transform 1 0 1796 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_626
timestamp 1710899220
transform 1 0 1764 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_627
timestamp 1710899220
transform 1 0 2004 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_628
timestamp 1710899220
transform 1 0 1972 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_629
timestamp 1710899220
transform 1 0 1948 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_630
timestamp 1710899220
transform 1 0 1812 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_631
timestamp 1710899220
transform 1 0 1796 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_632
timestamp 1710899220
transform 1 0 1836 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_633
timestamp 1710899220
transform 1 0 1716 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_634
timestamp 1710899220
transform 1 0 1676 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_635
timestamp 1710899220
transform 1 0 2012 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_636
timestamp 1710899220
transform 1 0 1980 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_637
timestamp 1710899220
transform 1 0 1820 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_638
timestamp 1710899220
transform 1 0 1788 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_639
timestamp 1710899220
transform 1 0 1756 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_640
timestamp 1710899220
transform 1 0 1652 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_641
timestamp 1710899220
transform 1 0 1644 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_642
timestamp 1710899220
transform 1 0 1556 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_643
timestamp 1710899220
transform 1 0 1396 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_644
timestamp 1710899220
transform 1 0 1835 0 1 924
box -2 -2 2 2
use M2_M1  M2_M1_645
timestamp 1710899220
transform 1 0 1804 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_646
timestamp 1710899220
transform 1 0 1516 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_647
timestamp 1710899220
transform 1 0 1460 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_648
timestamp 1710899220
transform 1 0 1396 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_649
timestamp 1710899220
transform 1 0 1684 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_650
timestamp 1710899220
transform 1 0 1676 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_651
timestamp 1710899220
transform 1 0 1644 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_652
timestamp 1710899220
transform 1 0 1876 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_653
timestamp 1710899220
transform 1 0 1772 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_654
timestamp 1710899220
transform 1 0 1724 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_655
timestamp 1710899220
transform 1 0 1628 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_656
timestamp 1710899220
transform 1 0 1524 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_657
timestamp 1710899220
transform 1 0 1980 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_658
timestamp 1710899220
transform 1 0 1948 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_659
timestamp 1710899220
transform 1 0 1828 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_660
timestamp 1710899220
transform 1 0 1764 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_661
timestamp 1710899220
transform 1 0 1756 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_662
timestamp 1710899220
transform 1 0 1988 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_663
timestamp 1710899220
transform 1 0 1956 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_664
timestamp 1710899220
transform 1 0 1932 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_665
timestamp 1710899220
transform 1 0 1820 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_666
timestamp 1710899220
transform 1 0 1796 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_667
timestamp 1710899220
transform 1 0 1780 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_668
timestamp 1710899220
transform 1 0 1740 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_669
timestamp 1710899220
transform 1 0 1524 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_670
timestamp 1710899220
transform 1 0 1428 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_671
timestamp 1710899220
transform 1 0 2028 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_672
timestamp 1710899220
transform 1 0 1860 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_673
timestamp 1710899220
transform 1 0 1788 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_674
timestamp 1710899220
transform 1 0 1564 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_675
timestamp 1710899220
transform 1 0 1508 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_676
timestamp 1710899220
transform 1 0 1508 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_677
timestamp 1710899220
transform 1 0 1428 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_678
timestamp 1710899220
transform 1 0 1596 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_679
timestamp 1710899220
transform 1 0 1548 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_680
timestamp 1710899220
transform 1 0 1532 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_681
timestamp 1710899220
transform 1 0 1556 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_682
timestamp 1710899220
transform 1 0 1500 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_683
timestamp 1710899220
transform 1 0 1492 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_684
timestamp 1710899220
transform 1 0 1748 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_685
timestamp 1710899220
transform 1 0 1748 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_686
timestamp 1710899220
transform 1 0 740 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_687
timestamp 1710899220
transform 1 0 700 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_688
timestamp 1710899220
transform 1 0 692 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_689
timestamp 1710899220
transform 1 0 380 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_690
timestamp 1710899220
transform 1 0 348 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_691
timestamp 1710899220
transform 1 0 348 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_692
timestamp 1710899220
transform 1 0 308 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_693
timestamp 1710899220
transform 1 0 332 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_694
timestamp 1710899220
transform 1 0 324 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_695
timestamp 1710899220
transform 1 0 284 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_696
timestamp 1710899220
transform 1 0 1132 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_697
timestamp 1710899220
transform 1 0 1132 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_698
timestamp 1710899220
transform 1 0 1011 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_699
timestamp 1710899220
transform 1 0 1004 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_700
timestamp 1710899220
transform 1 0 844 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_701
timestamp 1710899220
transform 1 0 780 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_702
timestamp 1710899220
transform 1 0 756 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_703
timestamp 1710899220
transform 1 0 548 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_704
timestamp 1710899220
transform 1 0 516 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_705
timestamp 1710899220
transform 1 0 348 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_706
timestamp 1710899220
transform 1 0 308 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_707
timestamp 1710899220
transform 1 0 420 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_708
timestamp 1710899220
transform 1 0 388 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_709
timestamp 1710899220
transform 1 0 356 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_710
timestamp 1710899220
transform 1 0 1012 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_711
timestamp 1710899220
transform 1 0 980 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_712
timestamp 1710899220
transform 1 0 1188 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_713
timestamp 1710899220
transform 1 0 1156 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_714
timestamp 1710899220
transform 1 0 1700 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_715
timestamp 1710899220
transform 1 0 1660 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_716
timestamp 1710899220
transform 1 0 1636 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_717
timestamp 1710899220
transform 1 0 1620 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_718
timestamp 1710899220
transform 1 0 1588 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_719
timestamp 1710899220
transform 1 0 1700 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_720
timestamp 1710899220
transform 1 0 1652 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_721
timestamp 1710899220
transform 1 0 1636 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_722
timestamp 1710899220
transform 1 0 1628 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_723
timestamp 1710899220
transform 1 0 2028 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_724
timestamp 1710899220
transform 1 0 1988 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_725
timestamp 1710899220
transform 1 0 1964 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_726
timestamp 1710899220
transform 1 0 1940 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_727
timestamp 1710899220
transform 1 0 1892 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_728
timestamp 1710899220
transform 1 0 2028 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_729
timestamp 1710899220
transform 1 0 1988 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_730
timestamp 1710899220
transform 1 0 1956 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_731
timestamp 1710899220
transform 1 0 1908 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_732
timestamp 1710899220
transform 1 0 2004 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_733
timestamp 1710899220
transform 1 0 1996 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_734
timestamp 1710899220
transform 1 0 1980 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_735
timestamp 1710899220
transform 1 0 1964 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_736
timestamp 1710899220
transform 1 0 1684 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_737
timestamp 1710899220
transform 1 0 1628 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_738
timestamp 1710899220
transform 1 0 1572 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_739
timestamp 1710899220
transform 1 0 1804 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_740
timestamp 1710899220
transform 1 0 1788 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_741
timestamp 1710899220
transform 1 0 1772 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_742
timestamp 1710899220
transform 1 0 1756 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_743
timestamp 1710899220
transform 1 0 1892 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_744
timestamp 1710899220
transform 1 0 1852 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_745
timestamp 1710899220
transform 1 0 1772 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_746
timestamp 1710899220
transform 1 0 1724 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_747
timestamp 1710899220
transform 1 0 1996 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_748
timestamp 1710899220
transform 1 0 1948 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_749
timestamp 1710899220
transform 1 0 1932 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_750
timestamp 1710899220
transform 1 0 2004 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_751
timestamp 1710899220
transform 1 0 1956 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_752
timestamp 1710899220
transform 1 0 1924 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_753
timestamp 1710899220
transform 1 0 1892 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_754
timestamp 1710899220
transform 1 0 2052 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_755
timestamp 1710899220
transform 1 0 2012 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_756
timestamp 1710899220
transform 1 0 1908 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_757
timestamp 1710899220
transform 1 0 1852 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_758
timestamp 1710899220
transform 1 0 2316 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_759
timestamp 1710899220
transform 1 0 2268 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_760
timestamp 1710899220
transform 1 0 2284 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_761
timestamp 1710899220
transform 1 0 2268 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_762
timestamp 1710899220
transform 1 0 2564 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_763
timestamp 1710899220
transform 1 0 2548 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_764
timestamp 1710899220
transform 1 0 2516 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_765
timestamp 1710899220
transform 1 0 2516 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_766
timestamp 1710899220
transform 1 0 2532 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_767
timestamp 1710899220
transform 1 0 2476 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_768
timestamp 1710899220
transform 1 0 2476 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_769
timestamp 1710899220
transform 1 0 2396 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_770
timestamp 1710899220
transform 1 0 2364 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_771
timestamp 1710899220
transform 1 0 2348 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_772
timestamp 1710899220
transform 1 0 2348 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_773
timestamp 1710899220
transform 1 0 2532 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_774
timestamp 1710899220
transform 1 0 2508 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_775
timestamp 1710899220
transform 1 0 2412 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_776
timestamp 1710899220
transform 1 0 2484 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_777
timestamp 1710899220
transform 1 0 2396 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_778
timestamp 1710899220
transform 1 0 2316 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_779
timestamp 1710899220
transform 1 0 2572 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_780
timestamp 1710899220
transform 1 0 2532 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_781
timestamp 1710899220
transform 1 0 2500 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_782
timestamp 1710899220
transform 1 0 2468 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_783
timestamp 1710899220
transform 1 0 2572 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_784
timestamp 1710899220
transform 1 0 2508 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_785
timestamp 1710899220
transform 1 0 2444 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_786
timestamp 1710899220
transform 1 0 2428 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_787
timestamp 1710899220
transform 1 0 2548 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_788
timestamp 1710899220
transform 1 0 2436 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_789
timestamp 1710899220
transform 1 0 2372 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_790
timestamp 1710899220
transform 1 0 2332 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_791
timestamp 1710899220
transform 1 0 2276 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_792
timestamp 1710899220
transform 1 0 2548 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_793
timestamp 1710899220
transform 1 0 2404 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_794
timestamp 1710899220
transform 1 0 2628 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_795
timestamp 1710899220
transform 1 0 2596 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_796
timestamp 1710899220
transform 1 0 2588 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_797
timestamp 1710899220
transform 1 0 2588 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_798
timestamp 1710899220
transform 1 0 2580 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_799
timestamp 1710899220
transform 1 0 2572 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_800
timestamp 1710899220
transform 1 0 2628 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_801
timestamp 1710899220
transform 1 0 2404 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_802
timestamp 1710899220
transform 1 0 2468 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_803
timestamp 1710899220
transform 1 0 2412 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_804
timestamp 1710899220
transform 1 0 2340 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_805
timestamp 1710899220
transform 1 0 2292 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_806
timestamp 1710899220
transform 1 0 2452 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_807
timestamp 1710899220
transform 1 0 2452 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_808
timestamp 1710899220
transform 1 0 2156 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_809
timestamp 1710899220
transform 1 0 2156 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_810
timestamp 1710899220
transform 1 0 2292 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_811
timestamp 1710899220
transform 1 0 2260 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_812
timestamp 1710899220
transform 1 0 2236 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_813
timestamp 1710899220
transform 1 0 2060 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_814
timestamp 1710899220
transform 1 0 2268 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_815
timestamp 1710899220
transform 1 0 2236 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_816
timestamp 1710899220
transform 1 0 2188 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_817
timestamp 1710899220
transform 1 0 2132 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_818
timestamp 1710899220
transform 1 0 2228 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_819
timestamp 1710899220
transform 1 0 2196 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_820
timestamp 1710899220
transform 1 0 2180 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_821
timestamp 1710899220
transform 1 0 2484 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_822
timestamp 1710899220
transform 1 0 2460 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_823
timestamp 1710899220
transform 1 0 1252 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_824
timestamp 1710899220
transform 1 0 1156 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_825
timestamp 1710899220
transform 1 0 1028 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_826
timestamp 1710899220
transform 1 0 948 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_827
timestamp 1710899220
transform 1 0 908 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_828
timestamp 1710899220
transform 1 0 1228 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_829
timestamp 1710899220
transform 1 0 1220 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_830
timestamp 1710899220
transform 1 0 1188 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_831
timestamp 1710899220
transform 1 0 1156 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_832
timestamp 1710899220
transform 1 0 1004 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_833
timestamp 1710899220
transform 1 0 900 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_834
timestamp 1710899220
transform 1 0 876 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_835
timestamp 1710899220
transform 1 0 1092 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_836
timestamp 1710899220
transform 1 0 940 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_837
timestamp 1710899220
transform 1 0 852 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_838
timestamp 1710899220
transform 1 0 700 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_839
timestamp 1710899220
transform 1 0 668 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_840
timestamp 1710899220
transform 1 0 516 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_841
timestamp 1710899220
transform 1 0 724 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_842
timestamp 1710899220
transform 1 0 716 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_843
timestamp 1710899220
transform 1 0 524 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_844
timestamp 1710899220
transform 1 0 444 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_845
timestamp 1710899220
transform 1 0 292 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_846
timestamp 1710899220
transform 1 0 284 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_847
timestamp 1710899220
transform 1 0 740 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_848
timestamp 1710899220
transform 1 0 700 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_849
timestamp 1710899220
transform 1 0 484 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_850
timestamp 1710899220
transform 1 0 268 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_851
timestamp 1710899220
transform 1 0 268 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_852
timestamp 1710899220
transform 1 0 228 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_853
timestamp 1710899220
transform 1 0 148 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_854
timestamp 1710899220
transform 1 0 236 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_855
timestamp 1710899220
transform 1 0 228 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_856
timestamp 1710899220
transform 1 0 356 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_857
timestamp 1710899220
transform 1 0 268 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_858
timestamp 1710899220
transform 1 0 268 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_859
timestamp 1710899220
transform 1 0 268 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_860
timestamp 1710899220
transform 1 0 484 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_861
timestamp 1710899220
transform 1 0 396 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_862
timestamp 1710899220
transform 1 0 292 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_863
timestamp 1710899220
transform 1 0 540 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_864
timestamp 1710899220
transform 1 0 524 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_865
timestamp 1710899220
transform 1 0 604 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_866
timestamp 1710899220
transform 1 0 588 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_867
timestamp 1710899220
transform 1 0 476 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_868
timestamp 1710899220
transform 1 0 540 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_869
timestamp 1710899220
transform 1 0 516 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_870
timestamp 1710899220
transform 1 0 660 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_871
timestamp 1710899220
transform 1 0 572 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_872
timestamp 1710899220
transform 1 0 532 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_873
timestamp 1710899220
transform 1 0 908 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_874
timestamp 1710899220
transform 1 0 908 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_875
timestamp 1710899220
transform 1 0 860 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_876
timestamp 1710899220
transform 1 0 780 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_877
timestamp 1710899220
transform 1 0 788 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_878
timestamp 1710899220
transform 1 0 700 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_879
timestamp 1710899220
transform 1 0 684 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_880
timestamp 1710899220
transform 1 0 796 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_881
timestamp 1710899220
transform 1 0 780 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_882
timestamp 1710899220
transform 1 0 860 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_883
timestamp 1710899220
transform 1 0 844 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_884
timestamp 1710899220
transform 1 0 980 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_885
timestamp 1710899220
transform 1 0 892 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_886
timestamp 1710899220
transform 1 0 852 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_887
timestamp 1710899220
transform 1 0 1252 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_888
timestamp 1710899220
transform 1 0 1236 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_889
timestamp 1710899220
transform 1 0 1164 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_890
timestamp 1710899220
transform 1 0 1076 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_891
timestamp 1710899220
transform 1 0 1060 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_892
timestamp 1710899220
transform 1 0 1108 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_893
timestamp 1710899220
transform 1 0 1020 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_894
timestamp 1710899220
transform 1 0 860 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_895
timestamp 1710899220
transform 1 0 1340 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_896
timestamp 1710899220
transform 1 0 1308 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_897
timestamp 1710899220
transform 1 0 1460 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_898
timestamp 1710899220
transform 1 0 1372 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_899
timestamp 1710899220
transform 1 0 1316 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_900
timestamp 1710899220
transform 1 0 1588 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_901
timestamp 1710899220
transform 1 0 1500 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_902
timestamp 1710899220
transform 1 0 1332 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_903
timestamp 1710899220
transform 1 0 1500 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_904
timestamp 1710899220
transform 1 0 1484 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_905
timestamp 1710899220
transform 1 0 1348 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_906
timestamp 1710899220
transform 1 0 1332 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_907
timestamp 1710899220
transform 1 0 1284 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_908
timestamp 1710899220
transform 1 0 1284 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_909
timestamp 1710899220
transform 1 0 1660 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_910
timestamp 1710899220
transform 1 0 1644 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_911
timestamp 1710899220
transform 1 0 1780 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_912
timestamp 1710899220
transform 1 0 1692 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_913
timestamp 1710899220
transform 1 0 1652 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_914
timestamp 1710899220
transform 1 0 1580 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_915
timestamp 1710899220
transform 1 0 1420 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_916
timestamp 1710899220
transform 1 0 1372 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_917
timestamp 1710899220
transform 1 0 1692 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_918
timestamp 1710899220
transform 1 0 1596 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_919
timestamp 1710899220
transform 1 0 1604 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_920
timestamp 1710899220
transform 1 0 1588 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_921
timestamp 1710899220
transform 1 0 1812 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_922
timestamp 1710899220
transform 1 0 1708 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_923
timestamp 1710899220
transform 1 0 1740 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_924
timestamp 1710899220
transform 1 0 1740 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_925
timestamp 1710899220
transform 1 0 1668 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_926
timestamp 1710899220
transform 1 0 1644 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_927
timestamp 1710899220
transform 1 0 1612 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_928
timestamp 1710899220
transform 1 0 1572 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_929
timestamp 1710899220
transform 1 0 1540 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_930
timestamp 1710899220
transform 1 0 1532 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_931
timestamp 1710899220
transform 1 0 1468 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_932
timestamp 1710899220
transform 1 0 1692 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_933
timestamp 1710899220
transform 1 0 1660 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_934
timestamp 1710899220
transform 1 0 1644 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_935
timestamp 1710899220
transform 1 0 1492 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_936
timestamp 1710899220
transform 1 0 1460 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_937
timestamp 1710899220
transform 1 0 1476 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_938
timestamp 1710899220
transform 1 0 1420 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_939
timestamp 1710899220
transform 1 0 1580 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_940
timestamp 1710899220
transform 1 0 1564 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_941
timestamp 1710899220
transform 1 0 1260 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_942
timestamp 1710899220
transform 1 0 1244 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_943
timestamp 1710899220
transform 1 0 1228 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_944
timestamp 1710899220
transform 1 0 1204 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_945
timestamp 1710899220
transform 1 0 1348 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_946
timestamp 1710899220
transform 1 0 1268 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_947
timestamp 1710899220
transform 1 0 1644 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_948
timestamp 1710899220
transform 1 0 1620 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_949
timestamp 1710899220
transform 1 0 1516 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_950
timestamp 1710899220
transform 1 0 1500 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_951
timestamp 1710899220
transform 1 0 1316 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_952
timestamp 1710899220
transform 1 0 1284 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_953
timestamp 1710899220
transform 1 0 2236 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_954
timestamp 1710899220
transform 1 0 2212 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_955
timestamp 1710899220
transform 1 0 2180 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_956
timestamp 1710899220
transform 1 0 2660 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_957
timestamp 1710899220
transform 1 0 2620 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_958
timestamp 1710899220
transform 1 0 2612 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_959
timestamp 1710899220
transform 1 0 2572 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_960
timestamp 1710899220
transform 1 0 2500 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_961
timestamp 1710899220
transform 1 0 2460 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_962
timestamp 1710899220
transform 1 0 2316 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_963
timestamp 1710899220
transform 1 0 2292 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_964
timestamp 1710899220
transform 1 0 2332 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_965
timestamp 1710899220
transform 1 0 2332 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_966
timestamp 1710899220
transform 1 0 2508 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_967
timestamp 1710899220
transform 1 0 2468 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_968
timestamp 1710899220
transform 1 0 2628 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_969
timestamp 1710899220
transform 1 0 2588 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_970
timestamp 1710899220
transform 1 0 2612 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_971
timestamp 1710899220
transform 1 0 2612 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_972
timestamp 1710899220
transform 1 0 2324 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_973
timestamp 1710899220
transform 1 0 2284 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_974
timestamp 1710899220
transform 1 0 2324 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_975
timestamp 1710899220
transform 1 0 2284 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_976
timestamp 1710899220
transform 1 0 2660 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_977
timestamp 1710899220
transform 1 0 2636 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_978
timestamp 1710899220
transform 1 0 2596 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_979
timestamp 1710899220
transform 1 0 2556 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_980
timestamp 1710899220
transform 1 0 2612 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_981
timestamp 1710899220
transform 1 0 2572 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_982
timestamp 1710899220
transform 1 0 2660 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_983
timestamp 1710899220
transform 1 0 2620 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_984
timestamp 1710899220
transform 1 0 2444 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_985
timestamp 1710899220
transform 1 0 2404 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_986
timestamp 1710899220
transform 1 0 2612 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_987
timestamp 1710899220
transform 1 0 2572 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_988
timestamp 1710899220
transform 1 0 2604 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_989
timestamp 1710899220
transform 1 0 2604 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_990
timestamp 1710899220
transform 1 0 2460 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_991
timestamp 1710899220
transform 1 0 2420 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_992
timestamp 1710899220
transform 1 0 2332 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_993
timestamp 1710899220
transform 1 0 2332 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_994
timestamp 1710899220
transform 1 0 2356 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_995
timestamp 1710899220
transform 1 0 2316 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_996
timestamp 1710899220
transform 1 0 2092 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_997
timestamp 1710899220
transform 1 0 2068 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_998
timestamp 1710899220
transform 1 0 2236 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_999
timestamp 1710899220
transform 1 0 2196 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1000
timestamp 1710899220
transform 1 0 1932 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1001
timestamp 1710899220
transform 1 0 1892 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1002
timestamp 1710899220
transform 1 0 1916 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1003
timestamp 1710899220
transform 1 0 1876 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1004
timestamp 1710899220
transform 1 0 1924 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1005
timestamp 1710899220
transform 1 0 1876 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1006
timestamp 1710899220
transform 1 0 1860 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1007
timestamp 1710899220
transform 1 0 1820 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1008
timestamp 1710899220
transform 1 0 1916 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1009
timestamp 1710899220
transform 1 0 1876 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1010
timestamp 1710899220
transform 1 0 2084 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1011
timestamp 1710899220
transform 1 0 2044 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1012
timestamp 1710899220
transform 1 0 2284 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1013
timestamp 1710899220
transform 1 0 2236 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1014
timestamp 1710899220
transform 1 0 2132 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1015
timestamp 1710899220
transform 1 0 2084 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1016
timestamp 1710899220
transform 1 0 2372 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1017
timestamp 1710899220
transform 1 0 2332 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1018
timestamp 1710899220
transform 1 0 2260 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1019
timestamp 1710899220
transform 1 0 2212 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1020
timestamp 1710899220
transform 1 0 1820 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1021
timestamp 1710899220
transform 1 0 1788 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1022
timestamp 1710899220
transform 1 0 1460 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1023
timestamp 1710899220
transform 1 0 1316 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1024
timestamp 1710899220
transform 1 0 1308 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1025
timestamp 1710899220
transform 1 0 1156 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1026
timestamp 1710899220
transform 1 0 1156 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1027
timestamp 1710899220
transform 1 0 2092 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1028
timestamp 1710899220
transform 1 0 2052 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1029
timestamp 1710899220
transform 1 0 2268 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1030
timestamp 1710899220
transform 1 0 2260 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1031
timestamp 1710899220
transform 1 0 2172 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1032
timestamp 1710899220
transform 1 0 2116 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1033
timestamp 1710899220
transform 1 0 2052 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1034
timestamp 1710899220
transform 1 0 2020 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1035
timestamp 1710899220
transform 1 0 1180 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1036
timestamp 1710899220
transform 1 0 916 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_1037
timestamp 1710899220
transform 1 0 868 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1038
timestamp 1710899220
transform 1 0 1092 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1039
timestamp 1710899220
transform 1 0 892 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1040
timestamp 1710899220
transform 1 0 844 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1041
timestamp 1710899220
transform 1 0 1716 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1042
timestamp 1710899220
transform 1 0 1716 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1043
timestamp 1710899220
transform 1 0 1700 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1044
timestamp 1710899220
transform 1 0 1044 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1045
timestamp 1710899220
transform 1 0 948 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1046
timestamp 1710899220
transform 1 0 844 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1047
timestamp 1710899220
transform 1 0 820 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1048
timestamp 1710899220
transform 1 0 812 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1049
timestamp 1710899220
transform 1 0 812 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1050
timestamp 1710899220
transform 1 0 1420 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1051
timestamp 1710899220
transform 1 0 1420 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1052
timestamp 1710899220
transform 1 0 1372 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1053
timestamp 1710899220
transform 1 0 1748 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1054
timestamp 1710899220
transform 1 0 1748 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1055
timestamp 1710899220
transform 1 0 1732 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1056
timestamp 1710899220
transform 1 0 692 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1057
timestamp 1710899220
transform 1 0 668 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1058
timestamp 1710899220
transform 1 0 660 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1059
timestamp 1710899220
transform 1 0 660 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_1060
timestamp 1710899220
transform 1 0 1076 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1061
timestamp 1710899220
transform 1 0 924 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1062
timestamp 1710899220
transform 1 0 924 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1063
timestamp 1710899220
transform 1 0 1180 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1064
timestamp 1710899220
transform 1 0 1148 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1065
timestamp 1710899220
transform 1 0 1148 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1066
timestamp 1710899220
transform 1 0 1156 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1067
timestamp 1710899220
transform 1 0 1108 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1068
timestamp 1710899220
transform 1 0 1100 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1069
timestamp 1710899220
transform 1 0 1900 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1070
timestamp 1710899220
transform 1 0 1852 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1071
timestamp 1710899220
transform 1 0 1804 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1072
timestamp 1710899220
transform 1 0 1716 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1073
timestamp 1710899220
transform 1 0 1716 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1074
timestamp 1710899220
transform 1 0 1692 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1075
timestamp 1710899220
transform 1 0 652 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1076
timestamp 1710899220
transform 1 0 628 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1077
timestamp 1710899220
transform 1 0 620 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1078
timestamp 1710899220
transform 1 0 620 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1079
timestamp 1710899220
transform 1 0 1084 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_1080
timestamp 1710899220
transform 1 0 1036 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1081
timestamp 1710899220
transform 1 0 1284 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1082
timestamp 1710899220
transform 1 0 1260 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1083
timestamp 1710899220
transform 1 0 1252 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1084
timestamp 1710899220
transform 1 0 1252 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1085
timestamp 1710899220
transform 1 0 1196 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1086
timestamp 1710899220
transform 1 0 1124 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1087
timestamp 1710899220
transform 1 0 1124 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1088
timestamp 1710899220
transform 1 0 1540 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1089
timestamp 1710899220
transform 1 0 1516 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1090
timestamp 1710899220
transform 1 0 1508 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1091
timestamp 1710899220
transform 1 0 1508 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1092
timestamp 1710899220
transform 1 0 1580 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1093
timestamp 1710899220
transform 1 0 1564 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1094
timestamp 1710899220
transform 1 0 1028 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1095
timestamp 1710899220
transform 1 0 980 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1096
timestamp 1710899220
transform 1 0 1060 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1097
timestamp 1710899220
transform 1 0 988 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1098
timestamp 1710899220
transform 1 0 988 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1099
timestamp 1710899220
transform 1 0 1372 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1100
timestamp 1710899220
transform 1 0 1324 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1101
timestamp 1710899220
transform 1 0 1324 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1102
timestamp 1710899220
transform 1 0 1380 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1103
timestamp 1710899220
transform 1 0 1348 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1104
timestamp 1710899220
transform 1 0 1332 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1105
timestamp 1710899220
transform 1 0 1644 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1106
timestamp 1710899220
transform 1 0 1644 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1107
timestamp 1710899220
transform 1 0 1612 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1108
timestamp 1710899220
transform 1 0 1596 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1109
timestamp 1710899220
transform 1 0 1836 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1110
timestamp 1710899220
transform 1 0 1788 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1111
timestamp 1710899220
transform 1 0 1708 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1112
timestamp 1710899220
transform 1 0 1668 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1113
timestamp 1710899220
transform 1 0 2588 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1114
timestamp 1710899220
transform 1 0 2572 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1115
timestamp 1710899220
transform 1 0 2540 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1116
timestamp 1710899220
transform 1 0 2476 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1117
timestamp 1710899220
transform 1 0 2444 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1118
timestamp 1710899220
transform 1 0 2420 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1119
timestamp 1710899220
transform 1 0 2396 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1120
timestamp 1710899220
transform 1 0 2340 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1121
timestamp 1710899220
transform 1 0 2300 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1122
timestamp 1710899220
transform 1 0 2292 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1123
timestamp 1710899220
transform 1 0 2284 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1124
timestamp 1710899220
transform 1 0 1980 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1125
timestamp 1710899220
transform 1 0 1892 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1126
timestamp 1710899220
transform 1 0 1844 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1127
timestamp 1710899220
transform 1 0 2588 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1128
timestamp 1710899220
transform 1 0 2588 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1129
timestamp 1710899220
transform 1 0 2588 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1130
timestamp 1710899220
transform 1 0 2588 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1131
timestamp 1710899220
transform 1 0 2572 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1132
timestamp 1710899220
transform 1 0 2572 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1133
timestamp 1710899220
transform 1 0 2564 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1134
timestamp 1710899220
transform 1 0 2436 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1135
timestamp 1710899220
transform 1 0 2420 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1136
timestamp 1710899220
transform 1 0 2332 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1137
timestamp 1710899220
transform 1 0 2308 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1138
timestamp 1710899220
transform 1 0 2284 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1139
timestamp 1710899220
transform 1 0 2236 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1140
timestamp 1710899220
transform 1 0 2236 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1141
timestamp 1710899220
transform 1 0 2348 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1142
timestamp 1710899220
transform 1 0 2252 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1143
timestamp 1710899220
transform 1 0 2212 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1144
timestamp 1710899220
transform 1 0 2164 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1145
timestamp 1710899220
transform 1 0 2124 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1146
timestamp 1710899220
transform 1 0 2068 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1147
timestamp 1710899220
transform 1 0 2036 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1148
timestamp 1710899220
transform 1 0 1996 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1149
timestamp 1710899220
transform 1 0 1964 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1150
timestamp 1710899220
transform 1 0 1844 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1151
timestamp 1710899220
transform 1 0 1828 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1152
timestamp 1710899220
transform 1 0 1828 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1153
timestamp 1710899220
transform 1 0 1828 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1154
timestamp 1710899220
transform 1 0 1772 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1155
timestamp 1710899220
transform 1 0 2068 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1156
timestamp 1710899220
transform 1 0 2068 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1157
timestamp 1710899220
transform 1 0 2068 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1158
timestamp 1710899220
transform 1 0 2052 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1159
timestamp 1710899220
transform 1 0 2044 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1160
timestamp 1710899220
transform 1 0 2044 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1161
timestamp 1710899220
transform 1 0 2020 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1162
timestamp 1710899220
transform 1 0 1956 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1163
timestamp 1710899220
transform 1 0 1916 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1164
timestamp 1710899220
transform 1 0 1724 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1165
timestamp 1710899220
transform 1 0 1676 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1166
timestamp 1710899220
transform 1 0 1676 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1167
timestamp 1710899220
transform 1 0 1572 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1168
timestamp 1710899220
transform 1 0 1564 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1169
timestamp 1710899220
transform 1 0 1236 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1170
timestamp 1710899220
transform 1 0 1172 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1171
timestamp 1710899220
transform 1 0 1156 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1172
timestamp 1710899220
transform 1 0 1060 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1173
timestamp 1710899220
transform 1 0 964 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1174
timestamp 1710899220
transform 1 0 924 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1175
timestamp 1710899220
transform 1 0 828 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1176
timestamp 1710899220
transform 1 0 596 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1177
timestamp 1710899220
transform 1 0 452 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1178
timestamp 1710899220
transform 1 0 244 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1179
timestamp 1710899220
transform 1 0 244 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1180
timestamp 1710899220
transform 1 0 188 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1181
timestamp 1710899220
transform 1 0 180 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1182
timestamp 1710899220
transform 1 0 180 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1183
timestamp 1710899220
transform 1 0 1972 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1184
timestamp 1710899220
transform 1 0 1860 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1185
timestamp 1710899220
transform 1 0 1852 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1186
timestamp 1710899220
transform 1 0 1844 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1187
timestamp 1710899220
transform 1 0 1772 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1188
timestamp 1710899220
transform 1 0 1564 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1189
timestamp 1710899220
transform 1 0 1524 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1190
timestamp 1710899220
transform 1 0 1468 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1191
timestamp 1710899220
transform 1 0 1468 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1192
timestamp 1710899220
transform 1 0 1436 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1193
timestamp 1710899220
transform 1 0 1436 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1194
timestamp 1710899220
transform 1 0 1364 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1195
timestamp 1710899220
transform 1 0 1324 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1196
timestamp 1710899220
transform 1 0 1268 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1197
timestamp 1710899220
transform 1 0 1260 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1198
timestamp 1710899220
transform 1 0 1164 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1199
timestamp 1710899220
transform 1 0 1116 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1200
timestamp 1710899220
transform 1 0 1076 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1201
timestamp 1710899220
transform 1 0 868 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1202
timestamp 1710899220
transform 1 0 860 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1203
timestamp 1710899220
transform 1 0 764 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1204
timestamp 1710899220
transform 1 0 748 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1205
timestamp 1710899220
transform 1 0 668 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1206
timestamp 1710899220
transform 1 0 580 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1207
timestamp 1710899220
transform 1 0 564 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1208
timestamp 1710899220
transform 1 0 556 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1209
timestamp 1710899220
transform 1 0 452 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1210
timestamp 1710899220
transform 1 0 412 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1211
timestamp 1710899220
transform 1 0 2180 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1212
timestamp 1710899220
transform 1 0 2140 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1213
timestamp 1710899220
transform 1 0 2044 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1214
timestamp 1710899220
transform 1 0 1948 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1215
timestamp 1710899220
transform 1 0 1900 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1216
timestamp 1710899220
transform 1 0 1884 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1217
timestamp 1710899220
transform 1 0 1796 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1218
timestamp 1710899220
transform 1 0 1588 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1219
timestamp 1710899220
transform 1 0 1396 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1220
timestamp 1710899220
transform 1 0 1364 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1221
timestamp 1710899220
transform 1 0 1228 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1222
timestamp 1710899220
transform 1 0 1228 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1223
timestamp 1710899220
transform 1 0 1212 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1224
timestamp 1710899220
transform 1 0 1108 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1225
timestamp 1710899220
transform 1 0 1764 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1226
timestamp 1710899220
transform 1 0 1444 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1227
timestamp 1710899220
transform 1 0 1204 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1228
timestamp 1710899220
transform 1 0 1020 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1229
timestamp 1710899220
transform 1 0 948 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1230
timestamp 1710899220
transform 1 0 924 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1231
timestamp 1710899220
transform 1 0 884 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1232
timestamp 1710899220
transform 1 0 844 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1233
timestamp 1710899220
transform 1 0 820 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1234
timestamp 1710899220
transform 1 0 780 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1235
timestamp 1710899220
transform 1 0 756 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1236
timestamp 1710899220
transform 1 0 700 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1237
timestamp 1710899220
transform 1 0 540 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1238
timestamp 1710899220
transform 1 0 476 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1239
timestamp 1710899220
transform 1 0 1852 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1240
timestamp 1710899220
transform 1 0 1820 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1241
timestamp 1710899220
transform 1 0 1804 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1242
timestamp 1710899220
transform 1 0 1772 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1243
timestamp 1710899220
transform 1 0 1764 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1244
timestamp 1710899220
transform 1 0 1684 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1245
timestamp 1710899220
transform 1 0 1644 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1246
timestamp 1710899220
transform 1 0 1604 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1247
timestamp 1710899220
transform 1 0 1444 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1248
timestamp 1710899220
transform 1 0 1412 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1249
timestamp 1710899220
transform 1 0 1236 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1250
timestamp 1710899220
transform 1 0 1148 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1251
timestamp 1710899220
transform 1 0 1036 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1252
timestamp 1710899220
transform 1 0 996 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1253
timestamp 1710899220
transform 1 0 1940 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1254
timestamp 1710899220
transform 1 0 1932 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1255
timestamp 1710899220
transform 1 0 2268 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1256
timestamp 1710899220
transform 1 0 2060 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1257
timestamp 1710899220
transform 1 0 2028 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1258
timestamp 1710899220
transform 1 0 2004 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1259
timestamp 1710899220
transform 1 0 1820 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1260
timestamp 1710899220
transform 1 0 1300 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1261
timestamp 1710899220
transform 1 0 1244 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1262
timestamp 1710899220
transform 1 0 1220 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1263
timestamp 1710899220
transform 1 0 1844 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1264
timestamp 1710899220
transform 1 0 1804 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1265
timestamp 1710899220
transform 1 0 1772 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1266
timestamp 1710899220
transform 1 0 1748 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1267
timestamp 1710899220
transform 1 0 1476 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1268
timestamp 1710899220
transform 1 0 1468 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1269
timestamp 1710899220
transform 1 0 1452 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1270
timestamp 1710899220
transform 1 0 1452 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1271
timestamp 1710899220
transform 1 0 1428 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1272
timestamp 1710899220
transform 1 0 1428 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1273
timestamp 1710899220
transform 1 0 1420 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_1274
timestamp 1710899220
transform 1 0 1404 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1275
timestamp 1710899220
transform 1 0 1396 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_1276
timestamp 1710899220
transform 1 0 1388 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1277
timestamp 1710899220
transform 1 0 1372 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1278
timestamp 1710899220
transform 1 0 1364 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_1279
timestamp 1710899220
transform 1 0 1324 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1280
timestamp 1710899220
transform 1 0 1284 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1281
timestamp 1710899220
transform 1 0 1268 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1282
timestamp 1710899220
transform 1 0 1220 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1283
timestamp 1710899220
transform 1 0 1124 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1284
timestamp 1710899220
transform 1 0 1004 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1285
timestamp 1710899220
transform 1 0 876 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1286
timestamp 1710899220
transform 1 0 828 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1287
timestamp 1710899220
transform 1 0 756 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1288
timestamp 1710899220
transform 1 0 724 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1289
timestamp 1710899220
transform 1 0 716 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_1290
timestamp 1710899220
transform 1 0 700 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1291
timestamp 1710899220
transform 1 0 684 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1292
timestamp 1710899220
transform 1 0 676 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1293
timestamp 1710899220
transform 1 0 660 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1294
timestamp 1710899220
transform 1 0 1812 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1295
timestamp 1710899220
transform 1 0 1804 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1296
timestamp 1710899220
transform 1 0 1764 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1297
timestamp 1710899220
transform 1 0 1764 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1298
timestamp 1710899220
transform 1 0 1764 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1299
timestamp 1710899220
transform 1 0 1548 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1300
timestamp 1710899220
transform 1 0 1532 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1301
timestamp 1710899220
transform 1 0 1492 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1302
timestamp 1710899220
transform 1 0 1420 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1303
timestamp 1710899220
transform 1 0 1404 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1304
timestamp 1710899220
transform 1 0 1396 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1305
timestamp 1710899220
transform 1 0 1332 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1306
timestamp 1710899220
transform 1 0 1316 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1307
timestamp 1710899220
transform 1 0 1292 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1308
timestamp 1710899220
transform 1 0 1172 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1309
timestamp 1710899220
transform 1 0 1100 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1310
timestamp 1710899220
transform 1 0 972 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1311
timestamp 1710899220
transform 1 0 868 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1312
timestamp 1710899220
transform 1 0 812 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1313
timestamp 1710899220
transform 1 0 812 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1314
timestamp 1710899220
transform 1 0 668 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1315
timestamp 1710899220
transform 1 0 636 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1316
timestamp 1710899220
transform 1 0 620 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1317
timestamp 1710899220
transform 1 0 612 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1318
timestamp 1710899220
transform 1 0 540 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1319
timestamp 1710899220
transform 1 0 524 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1320
timestamp 1710899220
transform 1 0 1148 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1321
timestamp 1710899220
transform 1 0 1124 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1322
timestamp 1710899220
transform 1 0 1092 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1323
timestamp 1710899220
transform 1 0 996 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1324
timestamp 1710899220
transform 1 0 956 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1325
timestamp 1710899220
transform 1 0 780 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1326
timestamp 1710899220
transform 1 0 740 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1327
timestamp 1710899220
transform 1 0 508 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1328
timestamp 1710899220
transform 1 0 348 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1329
timestamp 1710899220
transform 1 0 340 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1330
timestamp 1710899220
transform 1 0 276 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1331
timestamp 1710899220
transform 1 0 276 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1332
timestamp 1710899220
transform 1 0 276 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1333
timestamp 1710899220
transform 1 0 2004 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1334
timestamp 1710899220
transform 1 0 1988 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1335
timestamp 1710899220
transform 1 0 1980 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1336
timestamp 1710899220
transform 1 0 1964 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1337
timestamp 1710899220
transform 1 0 1956 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1338
timestamp 1710899220
transform 1 0 1948 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1339
timestamp 1710899220
transform 1 0 1860 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1340
timestamp 1710899220
transform 1 0 1852 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1341
timestamp 1710899220
transform 1 0 1812 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1342
timestamp 1710899220
transform 1 0 1660 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1343
timestamp 1710899220
transform 1 0 1652 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1344
timestamp 1710899220
transform 1 0 1628 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1345
timestamp 1710899220
transform 1 0 1580 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1346
timestamp 1710899220
transform 1 0 2620 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1347
timestamp 1710899220
transform 1 0 2556 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1348
timestamp 1710899220
transform 1 0 2532 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1349
timestamp 1710899220
transform 1 0 2532 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1350
timestamp 1710899220
transform 1 0 2532 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1351
timestamp 1710899220
transform 1 0 2532 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1352
timestamp 1710899220
transform 1 0 2532 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1353
timestamp 1710899220
transform 1 0 2516 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1354
timestamp 1710899220
transform 1 0 2516 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1355
timestamp 1710899220
transform 1 0 2516 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1356
timestamp 1710899220
transform 1 0 2516 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1357
timestamp 1710899220
transform 1 0 2444 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1358
timestamp 1710899220
transform 1 0 2348 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1359
timestamp 1710899220
transform 1 0 2348 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1360
timestamp 1710899220
transform 1 0 2340 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1361
timestamp 1710899220
transform 1 0 2324 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1362
timestamp 1710899220
transform 1 0 2316 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1363
timestamp 1710899220
transform 1 0 2292 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1364
timestamp 1710899220
transform 1 0 2284 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1365
timestamp 1710899220
transform 1 0 2572 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1366
timestamp 1710899220
transform 1 0 2452 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1367
timestamp 1710899220
transform 1 0 2300 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1368
timestamp 1710899220
transform 1 0 2268 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1369
timestamp 1710899220
transform 1 0 2268 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1370
timestamp 1710899220
transform 1 0 2252 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1371
timestamp 1710899220
transform 1 0 2236 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1372
timestamp 1710899220
transform 1 0 2140 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1373
timestamp 1710899220
transform 1 0 2140 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1374
timestamp 1710899220
transform 1 0 2140 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1375
timestamp 1710899220
transform 1 0 2116 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1376
timestamp 1710899220
transform 1 0 1948 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1377
timestamp 1710899220
transform 1 0 1940 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1378
timestamp 1710899220
transform 1 0 1940 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_1379
timestamp 1710899220
transform 1 0 1940 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1380
timestamp 1710899220
transform 1 0 1932 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1381
timestamp 1710899220
transform 1 0 1900 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1382
timestamp 1710899220
transform 1 0 1900 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1383
timestamp 1710899220
transform 1 0 1916 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1384
timestamp 1710899220
transform 1 0 1892 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1385
timestamp 1710899220
transform 1 0 1908 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1386
timestamp 1710899220
transform 1 0 1844 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1387
timestamp 1710899220
transform 1 0 1820 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_1388
timestamp 1710899220
transform 1 0 2172 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1389
timestamp 1710899220
transform 1 0 2076 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_1390
timestamp 1710899220
transform 1 0 2036 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1391
timestamp 1710899220
transform 1 0 2020 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1392
timestamp 1710899220
transform 1 0 2004 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_1393
timestamp 1710899220
transform 1 0 1988 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1394
timestamp 1710899220
transform 1 0 1964 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1395
timestamp 1710899220
transform 1 0 1940 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1396
timestamp 1710899220
transform 1 0 1932 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1397
timestamp 1710899220
transform 1 0 1844 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1398
timestamp 1710899220
transform 1 0 1612 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1399
timestamp 1710899220
transform 1 0 1180 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1400
timestamp 1710899220
transform 1 0 1156 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1401
timestamp 1710899220
transform 1 0 1028 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1402
timestamp 1710899220
transform 1 0 1004 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1403
timestamp 1710899220
transform 1 0 812 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1404
timestamp 1710899220
transform 1 0 716 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1405
timestamp 1710899220
transform 1 0 340 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1406
timestamp 1710899220
transform 1 0 332 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1407
timestamp 1710899220
transform 1 0 308 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1408
timestamp 1710899220
transform 1 0 1148 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1409
timestamp 1710899220
transform 1 0 1004 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_1410
timestamp 1710899220
transform 1 0 972 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1411
timestamp 1710899220
transform 1 0 924 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1412
timestamp 1710899220
transform 1 0 852 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1413
timestamp 1710899220
transform 1 0 828 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_1414
timestamp 1710899220
transform 1 0 828 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1415
timestamp 1710899220
transform 1 0 796 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1416
timestamp 1710899220
transform 1 0 684 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_1417
timestamp 1710899220
transform 1 0 644 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1418
timestamp 1710899220
transform 1 0 596 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1419
timestamp 1710899220
transform 1 0 596 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1420
timestamp 1710899220
transform 1 0 596 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_1421
timestamp 1710899220
transform 1 0 596 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1422
timestamp 1710899220
transform 1 0 572 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1423
timestamp 1710899220
transform 1 0 492 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1424
timestamp 1710899220
transform 1 0 444 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1425
timestamp 1710899220
transform 1 0 444 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1426
timestamp 1710899220
transform 1 0 1748 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1427
timestamp 1710899220
transform 1 0 1716 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1428
timestamp 1710899220
transform 1 0 1708 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1429
timestamp 1710899220
transform 1 0 1684 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1430
timestamp 1710899220
transform 1 0 1668 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1431
timestamp 1710899220
transform 1 0 1612 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1432
timestamp 1710899220
transform 1 0 1588 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1433
timestamp 1710899220
transform 1 0 1556 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1434
timestamp 1710899220
transform 1 0 1404 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1435
timestamp 1710899220
transform 1 0 1348 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1436
timestamp 1710899220
transform 1 0 1316 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1437
timestamp 1710899220
transform 1 0 1300 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1438
timestamp 1710899220
transform 1 0 1284 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1439
timestamp 1710899220
transform 1 0 1260 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1440
timestamp 1710899220
transform 1 0 1460 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1441
timestamp 1710899220
transform 1 0 1356 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1442
timestamp 1710899220
transform 1 0 1284 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1443
timestamp 1710899220
transform 1 0 1260 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1444
timestamp 1710899220
transform 1 0 1252 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1445
timestamp 1710899220
transform 1 0 1228 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1446
timestamp 1710899220
transform 1 0 1220 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1447
timestamp 1710899220
transform 1 0 1188 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1448
timestamp 1710899220
transform 1 0 1180 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1449
timestamp 1710899220
transform 1 0 1156 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1450
timestamp 1710899220
transform 1 0 1148 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1451
timestamp 1710899220
transform 1 0 1124 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1452
timestamp 1710899220
transform 1 0 1092 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1453
timestamp 1710899220
transform 1 0 1932 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1454
timestamp 1710899220
transform 1 0 1908 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1455
timestamp 1710899220
transform 1 0 2012 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1456
timestamp 1710899220
transform 1 0 1996 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1457
timestamp 1710899220
transform 1 0 1948 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1458
timestamp 1710899220
transform 1 0 1876 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1459
timestamp 1710899220
transform 1 0 2228 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1460
timestamp 1710899220
transform 1 0 2204 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1461
timestamp 1710899220
transform 1 0 2044 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1462
timestamp 1710899220
transform 1 0 1932 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1463
timestamp 1710899220
transform 1 0 1924 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1464
timestamp 1710899220
transform 1 0 1644 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1465
timestamp 1710899220
transform 1 0 1868 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1466
timestamp 1710899220
transform 1 0 1860 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1467
timestamp 1710899220
transform 1 0 1844 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1468
timestamp 1710899220
transform 1 0 1732 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1469
timestamp 1710899220
transform 1 0 1732 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1470
timestamp 1710899220
transform 1 0 1604 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1471
timestamp 1710899220
transform 1 0 1588 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1472
timestamp 1710899220
transform 1 0 1524 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1473
timestamp 1710899220
transform 1 0 1380 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1474
timestamp 1710899220
transform 1 0 1332 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1475
timestamp 1710899220
transform 1 0 1316 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1476
timestamp 1710899220
transform 1 0 1044 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1477
timestamp 1710899220
transform 1 0 1004 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1478
timestamp 1710899220
transform 1 0 988 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1479
timestamp 1710899220
transform 1 0 964 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1480
timestamp 1710899220
transform 1 0 940 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1481
timestamp 1710899220
transform 1 0 876 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1482
timestamp 1710899220
transform 1 0 852 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1483
timestamp 1710899220
transform 1 0 828 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1484
timestamp 1710899220
transform 1 0 676 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1485
timestamp 1710899220
transform 1 0 636 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1486
timestamp 1710899220
transform 1 0 2588 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1487
timestamp 1710899220
transform 1 0 2548 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1488
timestamp 1710899220
transform 1 0 2548 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1489
timestamp 1710899220
transform 1 0 2388 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1490
timestamp 1710899220
transform 1 0 2348 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1491
timestamp 1710899220
transform 1 0 2308 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1492
timestamp 1710899220
transform 1 0 2292 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1493
timestamp 1710899220
transform 1 0 2276 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1494
timestamp 1710899220
transform 1 0 2172 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1495
timestamp 1710899220
transform 1 0 2164 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1496
timestamp 1710899220
transform 1 0 2132 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1497
timestamp 1710899220
transform 1 0 2116 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1498
timestamp 1710899220
transform 1 0 2028 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1499
timestamp 1710899220
transform 1 0 1972 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1500
timestamp 1710899220
transform 1 0 1956 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1501
timestamp 1710899220
transform 1 0 1956 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1502
timestamp 1710899220
transform 1 0 1932 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1503
timestamp 1710899220
transform 1 0 2652 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1504
timestamp 1710899220
transform 1 0 2604 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1505
timestamp 1710899220
transform 1 0 2564 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1506
timestamp 1710899220
transform 1 0 2564 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1507
timestamp 1710899220
transform 1 0 2548 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1508
timestamp 1710899220
transform 1 0 2532 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1509
timestamp 1710899220
transform 1 0 2532 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1510
timestamp 1710899220
transform 1 0 2532 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1511
timestamp 1710899220
transform 1 0 2484 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1512
timestamp 1710899220
transform 1 0 2364 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1513
timestamp 1710899220
transform 1 0 2364 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1514
timestamp 1710899220
transform 1 0 2340 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1515
timestamp 1710899220
transform 1 0 2316 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1516
timestamp 1710899220
transform 1 0 2300 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1517
timestamp 1710899220
transform 1 0 2188 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1518
timestamp 1710899220
transform 1 0 2052 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1519
timestamp 1710899220
transform 1 0 1964 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1520
timestamp 1710899220
transform 1 0 1452 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1521
timestamp 1710899220
transform 1 0 1324 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_1522
timestamp 1710899220
transform 1 0 1260 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_1523
timestamp 1710899220
transform 1 0 1124 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1524
timestamp 1710899220
transform 1 0 1124 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1525
timestamp 1710899220
transform 1 0 1092 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_1526
timestamp 1710899220
transform 1 0 1068 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1527
timestamp 1710899220
transform 1 0 1044 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1528
timestamp 1710899220
transform 1 0 1012 0 1 785
box -2 -2 2 2
use M2_M1  M2_M1_1529
timestamp 1710899220
transform 1 0 2476 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_1530
timestamp 1710899220
transform 1 0 2404 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_1531
timestamp 1710899220
transform 1 0 2348 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_1532
timestamp 1710899220
transform 1 0 2348 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_1533
timestamp 1710899220
transform 1 0 2324 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1534
timestamp 1710899220
transform 1 0 2268 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1535
timestamp 1710899220
transform 1 0 2172 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1536
timestamp 1710899220
transform 1 0 2148 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1537
timestamp 1710899220
transform 1 0 1956 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_1538
timestamp 1710899220
transform 1 0 1916 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_1539
timestamp 1710899220
transform 1 0 148 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_1540
timestamp 1710899220
transform 1 0 140 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1541
timestamp 1710899220
transform 1 0 132 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1542
timestamp 1710899220
transform 1 0 2268 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1543
timestamp 1710899220
transform 1 0 2236 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1544
timestamp 1710899220
transform 1 0 2180 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1545
timestamp 1710899220
transform 1 0 2588 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1546
timestamp 1710899220
transform 1 0 2588 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1547
timestamp 1710899220
transform 1 0 2588 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1548
timestamp 1710899220
transform 1 0 2540 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1549
timestamp 1710899220
transform 1 0 2492 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1550
timestamp 1710899220
transform 1 0 2340 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1551
timestamp 1710899220
transform 1 0 2284 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1552
timestamp 1710899220
transform 1 0 2252 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1553
timestamp 1710899220
transform 1 0 2204 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1554
timestamp 1710899220
transform 1 0 2164 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1555
timestamp 1710899220
transform 1 0 2156 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1556
timestamp 1710899220
transform 1 0 2140 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1557
timestamp 1710899220
transform 1 0 2100 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1558
timestamp 1710899220
transform 1 0 2084 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1559
timestamp 1710899220
transform 1 0 220 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1560
timestamp 1710899220
transform 1 0 100 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1561
timestamp 1710899220
transform 1 0 100 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1562
timestamp 1710899220
transform 1 0 228 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_1563
timestamp 1710899220
transform 1 0 180 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1564
timestamp 1710899220
transform 1 0 220 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1565
timestamp 1710899220
transform 1 0 204 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1566
timestamp 1710899220
transform 1 0 180 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1567
timestamp 1710899220
transform 1 0 852 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1568
timestamp 1710899220
transform 1 0 804 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1569
timestamp 1710899220
transform 1 0 300 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1570
timestamp 1710899220
transform 1 0 204 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1571
timestamp 1710899220
transform 1 0 172 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1572
timestamp 1710899220
transform 1 0 412 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1573
timestamp 1710899220
transform 1 0 308 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1574
timestamp 1710899220
transform 1 0 276 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1575
timestamp 1710899220
transform 1 0 516 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1576
timestamp 1710899220
transform 1 0 420 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1577
timestamp 1710899220
transform 1 0 388 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1578
timestamp 1710899220
transform 1 0 1316 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1579
timestamp 1710899220
transform 1 0 1252 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1580
timestamp 1710899220
transform 1 0 244 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1581
timestamp 1710899220
transform 1 0 164 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1582
timestamp 1710899220
transform 1 0 140 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1583
timestamp 1710899220
transform 1 0 132 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1584
timestamp 1710899220
transform 1 0 132 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1585
timestamp 1710899220
transform 1 0 76 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1586
timestamp 1710899220
transform 1 0 1260 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_1587
timestamp 1710899220
transform 1 0 1212 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1588
timestamp 1710899220
transform 1 0 196 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1589
timestamp 1710899220
transform 1 0 132 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1590
timestamp 1710899220
transform 1 0 76 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1591
timestamp 1710899220
transform 1 0 148 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1592
timestamp 1710899220
transform 1 0 132 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1593
timestamp 1710899220
transform 1 0 164 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1594
timestamp 1710899220
transform 1 0 132 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1595
timestamp 1710899220
transform 1 0 340 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1596
timestamp 1710899220
transform 1 0 252 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1597
timestamp 1710899220
transform 1 0 220 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1598
timestamp 1710899220
transform 1 0 156 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_1599
timestamp 1710899220
transform 1 0 156 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1600
timestamp 1710899220
transform 1 0 348 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1601
timestamp 1710899220
transform 1 0 124 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1602
timestamp 1710899220
transform 1 0 492 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1603
timestamp 1710899220
transform 1 0 252 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1604
timestamp 1710899220
transform 1 0 644 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1605
timestamp 1710899220
transform 1 0 396 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1606
timestamp 1710899220
transform 1 0 964 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1607
timestamp 1710899220
transform 1 0 548 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1608
timestamp 1710899220
transform 1 0 1084 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1609
timestamp 1710899220
transform 1 0 868 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1610
timestamp 1710899220
transform 1 0 1204 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1611
timestamp 1710899220
transform 1 0 988 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1612
timestamp 1710899220
transform 1 0 1156 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1613
timestamp 1710899220
transform 1 0 1100 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1614
timestamp 1710899220
transform 1 0 244 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1615
timestamp 1710899220
transform 1 0 116 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1616
timestamp 1710899220
transform 1 0 236 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_1617
timestamp 1710899220
transform 1 0 228 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1618
timestamp 1710899220
transform 1 0 420 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1619
timestamp 1710899220
transform 1 0 244 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1620
timestamp 1710899220
transform 1 0 412 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_1621
timestamp 1710899220
transform 1 0 388 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1622
timestamp 1710899220
transform 1 0 420 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1623
timestamp 1710899220
transform 1 0 148 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1624
timestamp 1710899220
transform 1 0 412 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_1625
timestamp 1710899220
transform 1 0 316 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1626
timestamp 1710899220
transform 1 0 636 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1627
timestamp 1710899220
transform 1 0 380 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1628
timestamp 1710899220
transform 1 0 628 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_1629
timestamp 1710899220
transform 1 0 540 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1630
timestamp 1710899220
transform 1 0 652 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1631
timestamp 1710899220
transform 1 0 324 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1632
timestamp 1710899220
transform 1 0 636 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_1633
timestamp 1710899220
transform 1 0 540 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1634
timestamp 1710899220
transform 1 0 452 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1635
timestamp 1710899220
transform 1 0 308 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1636
timestamp 1710899220
transform 1 0 500 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1637
timestamp 1710899220
transform 1 0 500 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1638
timestamp 1710899220
transform 1 0 844 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1639
timestamp 1710899220
transform 1 0 532 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1640
timestamp 1710899220
transform 1 0 852 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1641
timestamp 1710899220
transform 1 0 836 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_1642
timestamp 1710899220
transform 1 0 892 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1643
timestamp 1710899220
transform 1 0 532 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1644
timestamp 1710899220
transform 1 0 884 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_1645
timestamp 1710899220
transform 1 0 748 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1646
timestamp 1710899220
transform 1 0 772 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1647
timestamp 1710899220
transform 1 0 548 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1648
timestamp 1710899220
transform 1 0 812 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1649
timestamp 1710899220
transform 1 0 740 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1650
timestamp 1710899220
transform 1 0 1044 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1651
timestamp 1710899220
transform 1 0 852 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1652
timestamp 1710899220
transform 1 0 1036 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_1653
timestamp 1710899220
transform 1 0 980 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1654
timestamp 1710899220
transform 1 0 724 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1655
timestamp 1710899220
transform 1 0 684 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1656
timestamp 1710899220
transform 1 0 972 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1657
timestamp 1710899220
transform 1 0 724 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1658
timestamp 1710899220
transform 1 0 1084 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1659
timestamp 1710899220
transform 1 0 948 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1660
timestamp 1710899220
transform 1 0 1124 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1661
timestamp 1710899220
transform 1 0 1108 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1662
timestamp 1710899220
transform 1 0 100 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1663
timestamp 1710899220
transform 1 0 100 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1664
timestamp 1710899220
transform 1 0 252 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1665
timestamp 1710899220
transform 1 0 140 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1666
timestamp 1710899220
transform 1 0 452 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1667
timestamp 1710899220
transform 1 0 316 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1668
timestamp 1710899220
transform 1 0 676 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1669
timestamp 1710899220
transform 1 0 436 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1670
timestamp 1710899220
transform 1 0 748 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1671
timestamp 1710899220
transform 1 0 732 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1672
timestamp 1710899220
transform 1 0 276 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1673
timestamp 1710899220
transform 1 0 132 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1674
timestamp 1710899220
transform 1 0 428 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1675
timestamp 1710899220
transform 1 0 324 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1676
timestamp 1710899220
transform 1 0 500 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1677
timestamp 1710899220
transform 1 0 428 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1678
timestamp 1710899220
transform 1 0 740 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_1679
timestamp 1710899220
transform 1 0 716 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1680
timestamp 1710899220
transform 1 0 700 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1681
timestamp 1710899220
transform 1 0 660 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1682
timestamp 1710899220
transform 1 0 476 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1683
timestamp 1710899220
transform 1 0 308 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1684
timestamp 1710899220
transform 1 0 660 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1685
timestamp 1710899220
transform 1 0 540 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1686
timestamp 1710899220
transform 1 0 820 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1687
timestamp 1710899220
transform 1 0 788 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1688
timestamp 1710899220
transform 1 0 652 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1689
timestamp 1710899220
transform 1 0 652 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_1690
timestamp 1710899220
transform 1 0 1092 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1691
timestamp 1710899220
transform 1 0 1092 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_1692
timestamp 1710899220
transform 1 0 884 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1693
timestamp 1710899220
transform 1 0 532 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1694
timestamp 1710899220
transform 1 0 852 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1695
timestamp 1710899220
transform 1 0 796 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1696
timestamp 1710899220
transform 1 0 980 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1697
timestamp 1710899220
transform 1 0 940 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1698
timestamp 1710899220
transform 1 0 1132 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1699
timestamp 1710899220
transform 1 0 1068 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1700
timestamp 1710899220
transform 1 0 1196 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1701
timestamp 1710899220
transform 1 0 1124 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1702
timestamp 1710899220
transform 1 0 908 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1703
timestamp 1710899220
transform 1 0 780 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1704
timestamp 1710899220
transform 1 0 948 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1705
timestamp 1710899220
transform 1 0 932 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1706
timestamp 1710899220
transform 1 0 1156 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1707
timestamp 1710899220
transform 1 0 1132 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1708
timestamp 1710899220
transform 1 0 1556 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1709
timestamp 1710899220
transform 1 0 1516 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1710
timestamp 1710899220
transform 1 0 1708 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1711
timestamp 1710899220
transform 1 0 1636 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1712
timestamp 1710899220
transform 1 0 1788 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1713
timestamp 1710899220
transform 1 0 1724 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1714
timestamp 1710899220
transform 1 0 1820 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_1715
timestamp 1710899220
transform 1 0 1700 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1716
timestamp 1710899220
transform 1 0 1604 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1717
timestamp 1710899220
transform 1 0 1404 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1718
timestamp 1710899220
transform 1 0 1628 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1719
timestamp 1710899220
transform 1 0 1548 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1720
timestamp 1710899220
transform 1 0 1716 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1721
timestamp 1710899220
transform 1 0 1676 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1722
timestamp 1710899220
transform 1 0 1804 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1723
timestamp 1710899220
transform 1 0 1764 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1724
timestamp 1710899220
transform 1 0 1372 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1725
timestamp 1710899220
transform 1 0 1332 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1726
timestamp 1710899220
transform 1 0 1524 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1727
timestamp 1710899220
transform 1 0 1428 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1728
timestamp 1710899220
transform 1 0 1612 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1729
timestamp 1710899220
transform 1 0 1572 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1730
timestamp 1710899220
transform 1 0 1484 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1731
timestamp 1710899220
transform 1 0 1444 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1732
timestamp 1710899220
transform 1 0 1188 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1733
timestamp 1710899220
transform 1 0 1148 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1734
timestamp 1710899220
transform 1 0 1276 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1735
timestamp 1710899220
transform 1 0 1228 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1736
timestamp 1710899220
transform 1 0 1132 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1737
timestamp 1710899220
transform 1 0 1092 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1738
timestamp 1710899220
transform 1 0 1004 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1739
timestamp 1710899220
transform 1 0 964 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1740
timestamp 1710899220
transform 1 0 972 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1741
timestamp 1710899220
transform 1 0 940 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1742
timestamp 1710899220
transform 1 0 820 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1743
timestamp 1710899220
transform 1 0 764 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1744
timestamp 1710899220
transform 1 0 812 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1745
timestamp 1710899220
transform 1 0 772 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1746
timestamp 1710899220
transform 1 0 684 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1747
timestamp 1710899220
transform 1 0 644 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1748
timestamp 1710899220
transform 1 0 644 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1749
timestamp 1710899220
transform 1 0 636 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1750
timestamp 1710899220
transform 1 0 564 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1751
timestamp 1710899220
transform 1 0 500 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1752
timestamp 1710899220
transform 1 0 508 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1753
timestamp 1710899220
transform 1 0 468 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1754
timestamp 1710899220
transform 1 0 380 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1755
timestamp 1710899220
transform 1 0 340 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1756
timestamp 1710899220
transform 1 0 372 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1757
timestamp 1710899220
transform 1 0 364 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1758
timestamp 1710899220
transform 1 0 268 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1759
timestamp 1710899220
transform 1 0 220 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1760
timestamp 1710899220
transform 1 0 220 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1761
timestamp 1710899220
transform 1 0 132 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1762
timestamp 1710899220
transform 1 0 204 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1763
timestamp 1710899220
transform 1 0 124 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1764
timestamp 1710899220
transform 1 0 404 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1765
timestamp 1710899220
transform 1 0 404 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1766
timestamp 1710899220
transform 1 0 428 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1767
timestamp 1710899220
transform 1 0 276 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1768
timestamp 1710899220
transform 1 0 292 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1769
timestamp 1710899220
transform 1 0 244 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1770
timestamp 1710899220
transform 1 0 708 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1771
timestamp 1710899220
transform 1 0 708 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1772
timestamp 1710899220
transform 1 0 732 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1773
timestamp 1710899220
transform 1 0 580 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1774
timestamp 1710899220
transform 1 0 596 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1775
timestamp 1710899220
transform 1 0 548 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1776
timestamp 1710899220
transform 1 0 1140 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1777
timestamp 1710899220
transform 1 0 1028 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1778
timestamp 1710899220
transform 1 0 1044 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1779
timestamp 1710899220
transform 1 0 900 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_1780
timestamp 1710899220
transform 1 0 916 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1781
timestamp 1710899220
transform 1 0 868 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1782
timestamp 1710899220
transform 1 0 1500 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1783
timestamp 1710899220
transform 1 0 1476 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1784
timestamp 1710899220
transform 1 0 1532 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1785
timestamp 1710899220
transform 1 0 1380 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1786
timestamp 1710899220
transform 1 0 1396 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1787
timestamp 1710899220
transform 1 0 1348 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1788
timestamp 1710899220
transform 1 0 1572 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1789
timestamp 1710899220
transform 1 0 1572 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1790
timestamp 1710899220
transform 1 0 1692 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1791
timestamp 1710899220
transform 1 0 1628 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1792
timestamp 1710899220
transform 1 0 1716 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1793
timestamp 1710899220
transform 1 0 1668 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1794
timestamp 1710899220
transform 1 0 1740 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1795
timestamp 1710899220
transform 1 0 1732 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1796
timestamp 1710899220
transform 1 0 1756 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1797
timestamp 1710899220
transform 1 0 1756 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1798
timestamp 1710899220
transform 1 0 1788 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_1799
timestamp 1710899220
transform 1 0 1716 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1800
timestamp 1710899220
transform 1 0 2236 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1801
timestamp 1710899220
transform 1 0 2220 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1802
timestamp 1710899220
transform 1 0 2084 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1803
timestamp 1710899220
transform 1 0 2068 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_1804
timestamp 1710899220
transform 1 0 1588 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1805
timestamp 1710899220
transform 1 0 1516 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1806
timestamp 1710899220
transform 1 0 1428 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1807
timestamp 1710899220
transform 1 0 1396 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1808
timestamp 1710899220
transform 1 0 1380 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1809
timestamp 1710899220
transform 1 0 1516 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1810
timestamp 1710899220
transform 1 0 1476 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1811
timestamp 1710899220
transform 1 0 1460 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1812
timestamp 1710899220
transform 1 0 1420 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1813
timestamp 1710899220
transform 1 0 1340 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_1814
timestamp 1710899220
transform 1 0 1436 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1815
timestamp 1710899220
transform 1 0 1404 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1816
timestamp 1710899220
transform 1 0 1356 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1817
timestamp 1710899220
transform 1 0 1332 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1818
timestamp 1710899220
transform 1 0 1252 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_1819
timestamp 1710899220
transform 1 0 1260 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1820
timestamp 1710899220
transform 1 0 1220 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1821
timestamp 1710899220
transform 1 0 1140 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1822
timestamp 1710899220
transform 1 0 1100 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_1823
timestamp 1710899220
transform 1 0 1092 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1824
timestamp 1710899220
transform 1 0 996 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1825
timestamp 1710899220
transform 1 0 980 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1826
timestamp 1710899220
transform 1 0 956 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1827
timestamp 1710899220
transform 1 0 892 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_1828
timestamp 1710899220
transform 1 0 884 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1829
timestamp 1710899220
transform 1 0 700 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1830
timestamp 1710899220
transform 1 0 660 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1831
timestamp 1710899220
transform 1 0 636 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1832
timestamp 1710899220
transform 1 0 532 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1833
timestamp 1710899220
transform 1 0 508 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1834
timestamp 1710899220
transform 1 0 452 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1835
timestamp 1710899220
transform 1 0 428 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1836
timestamp 1710899220
transform 1 0 388 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1837
timestamp 1710899220
transform 1 0 364 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1838
timestamp 1710899220
transform 1 0 292 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_1839
timestamp 1710899220
transform 1 0 340 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1840
timestamp 1710899220
transform 1 0 332 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1841
timestamp 1710899220
transform 1 0 316 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1842
timestamp 1710899220
transform 1 0 244 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1843
timestamp 1710899220
transform 1 0 228 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1844
timestamp 1710899220
transform 1 0 220 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1845
timestamp 1710899220
transform 1 0 196 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1846
timestamp 1710899220
transform 1 0 132 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1847
timestamp 1710899220
transform 1 0 124 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1848
timestamp 1710899220
transform 1 0 180 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1849
timestamp 1710899220
transform 1 0 132 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1850
timestamp 1710899220
transform 1 0 76 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1851
timestamp 1710899220
transform 1 0 2124 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1852
timestamp 1710899220
transform 1 0 2004 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1853
timestamp 1710899220
transform 1 0 2092 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1854
timestamp 1710899220
transform 1 0 2036 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1855
timestamp 1710899220
transform 1 0 2012 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1856
timestamp 1710899220
transform 1 0 1948 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1857
timestamp 1710899220
transform 1 0 2068 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1858
timestamp 1710899220
transform 1 0 2028 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1859
timestamp 1710899220
transform 1 0 2220 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1860
timestamp 1710899220
transform 1 0 2188 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1861
timestamp 1710899220
transform 1 0 2244 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1862
timestamp 1710899220
transform 1 0 2228 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1863
timestamp 1710899220
transform 1 0 2060 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1864
timestamp 1710899220
transform 1 0 1988 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1865
timestamp 1710899220
transform 1 0 220 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1866
timestamp 1710899220
transform 1 0 148 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1867
timestamp 1710899220
transform 1 0 124 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1868
timestamp 1710899220
transform 1 0 252 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1869
timestamp 1710899220
transform 1 0 212 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_1870
timestamp 1710899220
transform 1 0 180 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1871
timestamp 1710899220
transform 1 0 364 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1872
timestamp 1710899220
transform 1 0 340 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_1873
timestamp 1710899220
transform 1 0 284 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1874
timestamp 1710899220
transform 1 0 484 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1875
timestamp 1710899220
transform 1 0 484 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_1876
timestamp 1710899220
transform 1 0 460 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1877
timestamp 1710899220
transform 1 0 396 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1878
timestamp 1710899220
transform 1 0 636 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_1879
timestamp 1710899220
transform 1 0 540 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1880
timestamp 1710899220
transform 1 0 500 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1881
timestamp 1710899220
transform 1 0 956 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_1882
timestamp 1710899220
transform 1 0 788 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1883
timestamp 1710899220
transform 1 0 1076 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_1884
timestamp 1710899220
transform 1 0 996 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1885
timestamp 1710899220
transform 1 0 1196 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_1886
timestamp 1710899220
transform 1 0 1148 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1887
timestamp 1710899220
transform 1 0 1212 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1888
timestamp 1710899220
transform 1 0 1204 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1889
timestamp 1710899220
transform 1 0 1372 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1890
timestamp 1710899220
transform 1 0 1300 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1891
timestamp 1710899220
transform 1 0 1284 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1892
timestamp 1710899220
transform 1 0 2308 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_1893
timestamp 1710899220
transform 1 0 2204 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1894
timestamp 1710899220
transform 1 0 2156 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1895
timestamp 1710899220
transform 1 0 2076 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1896
timestamp 1710899220
transform 1 0 1892 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1897
timestamp 1710899220
transform 1 0 1764 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1898
timestamp 1710899220
transform 1 0 1596 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1899
timestamp 1710899220
transform 1 0 1548 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1900
timestamp 1710899220
transform 1 0 1532 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1901
timestamp 1710899220
transform 1 0 1500 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_1902
timestamp 1710899220
transform 1 0 1420 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1903
timestamp 1710899220
transform 1 0 1348 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1904
timestamp 1710899220
transform 1 0 1340 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1905
timestamp 1710899220
transform 1 0 1268 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1906
timestamp 1710899220
transform 1 0 1164 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1907
timestamp 1710899220
transform 1 0 1140 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1908
timestamp 1710899220
transform 1 0 1116 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1909
timestamp 1710899220
transform 1 0 980 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1910
timestamp 1710899220
transform 1 0 940 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1911
timestamp 1710899220
transform 1 0 1356 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1912
timestamp 1710899220
transform 1 0 1036 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1913
timestamp 1710899220
transform 1 0 1388 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1914
timestamp 1710899220
transform 1 0 1340 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1915
timestamp 1710899220
transform 1 0 2044 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1916
timestamp 1710899220
transform 1 0 1676 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1917
timestamp 1710899220
transform 1 0 1580 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1918
timestamp 1710899220
transform 1 0 1444 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1919
timestamp 1710899220
transform 1 0 1564 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1920
timestamp 1710899220
transform 1 0 1548 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1921
timestamp 1710899220
transform 1 0 1380 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1922
timestamp 1710899220
transform 1 0 1372 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1923
timestamp 1710899220
transform 1 0 1236 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1924
timestamp 1710899220
transform 1 0 692 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_1925
timestamp 1710899220
transform 1 0 668 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1926
timestamp 1710899220
transform 1 0 1092 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1927
timestamp 1710899220
transform 1 0 708 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1928
timestamp 1710899220
transform 1 0 1284 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1929
timestamp 1710899220
transform 1 0 1164 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1930
timestamp 1710899220
transform 1 0 1100 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1931
timestamp 1710899220
transform 1 0 1068 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1932
timestamp 1710899220
transform 1 0 1692 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1933
timestamp 1710899220
transform 1 0 1660 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1934
timestamp 1710899220
transform 1 0 1636 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1935
timestamp 1710899220
transform 1 0 1228 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1936
timestamp 1710899220
transform 1 0 1196 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1937
timestamp 1710899220
transform 1 0 1108 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1938
timestamp 1710899220
transform 1 0 1060 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1939
timestamp 1710899220
transform 1 0 956 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1940
timestamp 1710899220
transform 1 0 932 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1941
timestamp 1710899220
transform 1 0 1148 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1942
timestamp 1710899220
transform 1 0 1076 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1943
timestamp 1710899220
transform 1 0 1308 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1944
timestamp 1710899220
transform 1 0 1156 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1945
timestamp 1710899220
transform 1 0 1132 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1946
timestamp 1710899220
transform 1 0 1132 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1947
timestamp 1710899220
transform 1 0 652 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1948
timestamp 1710899220
transform 1 0 628 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1949
timestamp 1710899220
transform 1 0 1124 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1950
timestamp 1710899220
transform 1 0 660 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1951
timestamp 1710899220
transform 1 0 1580 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1952
timestamp 1710899220
transform 1 0 1564 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1953
timestamp 1710899220
transform 1 0 1532 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1954
timestamp 1710899220
transform 1 0 1260 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1955
timestamp 1710899220
transform 1 0 1212 0 1 1755
box -2 -2 2 2
use M2_M1  M2_M1_1956
timestamp 1710899220
transform 1 0 1140 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1957
timestamp 1710899220
transform 1 0 1108 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1958
timestamp 1710899220
transform 1 0 1156 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1959
timestamp 1710899220
transform 1 0 1124 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1960
timestamp 1710899220
transform 1 0 1188 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1961
timestamp 1710899220
transform 1 0 1036 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1962
timestamp 1710899220
transform 1 0 1724 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1963
timestamp 1710899220
transform 1 0 1684 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1964
timestamp 1710899220
transform 1 0 1644 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1965
timestamp 1710899220
transform 1 0 1324 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1966
timestamp 1710899220
transform 1 0 1292 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1967
timestamp 1710899220
transform 1 0 1172 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1968
timestamp 1710899220
transform 1 0 1164 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1969
timestamp 1710899220
transform 1 0 1404 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1970
timestamp 1710899220
transform 1 0 1300 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1971
timestamp 1710899220
transform 1 0 1268 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1972
timestamp 1710899220
transform 1 0 1020 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1973
timestamp 1710899220
transform 1 0 996 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1974
timestamp 1710899220
transform 1 0 1180 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1975
timestamp 1710899220
transform 1 0 1060 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1976
timestamp 1710899220
transform 1 0 1228 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1977
timestamp 1710899220
transform 1 0 1172 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1978
timestamp 1710899220
transform 1 0 1588 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1979
timestamp 1710899220
transform 1 0 1580 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1980
timestamp 1710899220
transform 1 0 1252 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1981
timestamp 1710899220
transform 1 0 1188 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1982
timestamp 1710899220
transform 1 0 844 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1983
timestamp 1710899220
transform 1 0 820 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1984
timestamp 1710899220
transform 1 0 1260 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1985
timestamp 1710899220
transform 1 0 852 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1986
timestamp 1710899220
transform 1 0 1180 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1987
timestamp 1710899220
transform 1 0 1156 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1988
timestamp 1710899220
transform 1 0 1252 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1989
timestamp 1710899220
transform 1 0 1180 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1990
timestamp 1710899220
transform 1 0 1292 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1991
timestamp 1710899220
transform 1 0 1284 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1992
timestamp 1710899220
transform 1 0 1252 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1993
timestamp 1710899220
transform 1 0 1236 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1994
timestamp 1710899220
transform 1 0 1132 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1995
timestamp 1710899220
transform 1 0 1108 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1996
timestamp 1710899220
transform 1 0 1220 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1997
timestamp 1710899220
transform 1 0 1164 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1998
timestamp 1710899220
transform 1 0 1324 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1999
timestamp 1710899220
transform 1 0 1324 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2000
timestamp 1710899220
transform 1 0 1212 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2001
timestamp 1710899220
transform 1 0 1204 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2002
timestamp 1710899220
transform 1 0 1284 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2003
timestamp 1710899220
transform 1 0 1260 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2004
timestamp 1710899220
transform 1 0 1292 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2005
timestamp 1710899220
transform 1 0 1284 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2006
timestamp 1710899220
transform 1 0 1156 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2007
timestamp 1710899220
transform 1 0 1132 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2008
timestamp 1710899220
transform 1 0 1244 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2009
timestamp 1710899220
transform 1 0 1196 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2010
timestamp 1710899220
transform 1 0 1316 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2011
timestamp 1710899220
transform 1 0 1316 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2012
timestamp 1710899220
transform 1 0 1412 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2013
timestamp 1710899220
transform 1 0 1340 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2014
timestamp 1710899220
transform 1 0 1316 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2015
timestamp 1710899220
transform 1 0 1300 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2016
timestamp 1710899220
transform 1 0 1284 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2017
timestamp 1710899220
transform 1 0 1092 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2018
timestamp 1710899220
transform 1 0 1788 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2019
timestamp 1710899220
transform 1 0 1684 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2020
timestamp 1710899220
transform 1 0 1652 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2021
timestamp 1710899220
transform 1 0 1652 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2022
timestamp 1710899220
transform 1 0 1532 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2023
timestamp 1710899220
transform 1 0 1508 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2024
timestamp 1710899220
transform 1 0 1748 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2025
timestamp 1710899220
transform 1 0 1724 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2026
timestamp 1710899220
transform 1 0 1716 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2027
timestamp 1710899220
transform 1 0 1684 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2028
timestamp 1710899220
transform 1 0 1716 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2029
timestamp 1710899220
transform 1 0 1692 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2030
timestamp 1710899220
transform 1 0 1556 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2031
timestamp 1710899220
transform 1 0 1532 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2032
timestamp 1710899220
transform 1 0 1636 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_2033
timestamp 1710899220
transform 1 0 1636 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2034
timestamp 1710899220
transform 1 0 1612 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2035
timestamp 1710899220
transform 1 0 1572 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2036
timestamp 1710899220
transform 1 0 1572 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2037
timestamp 1710899220
transform 1 0 1540 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2038
timestamp 1710899220
transform 1 0 1516 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2039
timestamp 1710899220
transform 1 0 1556 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2040
timestamp 1710899220
transform 1 0 1548 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2041
timestamp 1710899220
transform 1 0 1612 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2042
timestamp 1710899220
transform 1 0 1572 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2043
timestamp 1710899220
transform 1 0 1588 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2044
timestamp 1710899220
transform 1 0 1548 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2045
timestamp 1710899220
transform 1 0 1668 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2046
timestamp 1710899220
transform 1 0 1628 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2047
timestamp 1710899220
transform 1 0 1524 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2048
timestamp 1710899220
transform 1 0 1500 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2049
timestamp 1710899220
transform 1 0 1484 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2050
timestamp 1710899220
transform 1 0 1484 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2051
timestamp 1710899220
transform 1 0 1860 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2052
timestamp 1710899220
transform 1 0 1820 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2053
timestamp 1710899220
transform 1 0 1748 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2054
timestamp 1710899220
transform 1 0 1724 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2055
timestamp 1710899220
transform 1 0 1676 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2056
timestamp 1710899220
transform 1 0 1620 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2057
timestamp 1710899220
transform 1 0 1780 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2058
timestamp 1710899220
transform 1 0 1756 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2059
timestamp 1710899220
transform 1 0 1716 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2060
timestamp 1710899220
transform 1 0 1580 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2061
timestamp 1710899220
transform 1 0 2148 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2062
timestamp 1710899220
transform 1 0 2108 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2063
timestamp 1710899220
transform 1 0 2028 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2064
timestamp 1710899220
transform 1 0 1540 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_2065
timestamp 1710899220
transform 1 0 1524 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2066
timestamp 1710899220
transform 1 0 1380 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2067
timestamp 1710899220
transform 1 0 1340 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2068
timestamp 1710899220
transform 1 0 1924 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2069
timestamp 1710899220
transform 1 0 1604 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2070
timestamp 1710899220
transform 1 0 1540 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2071
timestamp 1710899220
transform 1 0 1420 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2072
timestamp 1710899220
transform 1 0 1340 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2073
timestamp 1710899220
transform 1 0 1332 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2074
timestamp 1710899220
transform 1 0 1372 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2075
timestamp 1710899220
transform 1 0 1348 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2076
timestamp 1710899220
transform 1 0 1572 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2077
timestamp 1710899220
transform 1 0 1548 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2078
timestamp 1710899220
transform 1 0 1452 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2079
timestamp 1710899220
transform 1 0 1428 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2080
timestamp 1710899220
transform 1 0 2148 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2081
timestamp 1710899220
transform 1 0 2132 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2082
timestamp 1710899220
transform 1 0 2236 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2083
timestamp 1710899220
transform 1 0 2180 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_2084
timestamp 1710899220
transform 1 0 2172 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2085
timestamp 1710899220
transform 1 0 2164 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2086
timestamp 1710899220
transform 1 0 2140 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_2087
timestamp 1710899220
transform 1 0 2132 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2088
timestamp 1710899220
transform 1 0 2148 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2089
timestamp 1710899220
transform 1 0 2036 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2090
timestamp 1710899220
transform 1 0 2244 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2091
timestamp 1710899220
transform 1 0 2156 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_2092
timestamp 1710899220
transform 1 0 2300 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2093
timestamp 1710899220
transform 1 0 2268 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2094
timestamp 1710899220
transform 1 0 2212 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2095
timestamp 1710899220
transform 1 0 2212 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2096
timestamp 1710899220
transform 1 0 2244 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2097
timestamp 1710899220
transform 1 0 2220 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_2098
timestamp 1710899220
transform 1 0 2364 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2099
timestamp 1710899220
transform 1 0 2324 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2100
timestamp 1710899220
transform 1 0 980 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2101
timestamp 1710899220
transform 1 0 892 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2102
timestamp 1710899220
transform 1 0 692 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2103
timestamp 1710899220
transform 1 0 588 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2104
timestamp 1710899220
transform 1 0 964 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2105
timestamp 1710899220
transform 1 0 868 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2106
timestamp 1710899220
transform 1 0 652 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2107
timestamp 1710899220
transform 1 0 524 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2108
timestamp 1710899220
transform 1 0 1060 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2109
timestamp 1710899220
transform 1 0 996 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2110
timestamp 1710899220
transform 1 0 1004 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2111
timestamp 1710899220
transform 1 0 932 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2112
timestamp 1710899220
transform 1 0 1028 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2113
timestamp 1710899220
transform 1 0 972 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2114
timestamp 1710899220
transform 1 0 892 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2115
timestamp 1710899220
transform 1 0 828 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2116
timestamp 1710899220
transform 1 0 844 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2117
timestamp 1710899220
transform 1 0 748 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2118
timestamp 1710899220
transform 1 0 1180 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2119
timestamp 1710899220
transform 1 0 1084 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2120
timestamp 1710899220
transform 1 0 1132 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2121
timestamp 1710899220
transform 1 0 1044 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2122
timestamp 1710899220
transform 1 0 1284 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2123
timestamp 1710899220
transform 1 0 1196 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2124
timestamp 1710899220
transform 1 0 1156 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2125
timestamp 1710899220
transform 1 0 1068 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2126
timestamp 1710899220
transform 1 0 1348 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2127
timestamp 1710899220
transform 1 0 1276 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2128
timestamp 1710899220
transform 1 0 1420 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2129
timestamp 1710899220
transform 1 0 1356 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2130
timestamp 1710899220
transform 1 0 868 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2131
timestamp 1710899220
transform 1 0 804 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2132
timestamp 1710899220
transform 1 0 1468 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2133
timestamp 1710899220
transform 1 0 1396 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2134
timestamp 1710899220
transform 1 0 1876 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2135
timestamp 1710899220
transform 1 0 1876 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2136
timestamp 1710899220
transform 1 0 1788 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2137
timestamp 1710899220
transform 1 0 1748 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2138
timestamp 1710899220
transform 1 0 1540 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2139
timestamp 1710899220
transform 1 0 1468 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2140
timestamp 1710899220
transform 1 0 1668 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2141
timestamp 1710899220
transform 1 0 1628 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2142
timestamp 1710899220
transform 1 0 1620 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2143
timestamp 1710899220
transform 1 0 1620 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2144
timestamp 1710899220
transform 1 0 1908 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2145
timestamp 1710899220
transform 1 0 1868 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2146
timestamp 1710899220
transform 1 0 1796 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2147
timestamp 1710899220
transform 1 0 1756 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2148
timestamp 1710899220
transform 1 0 1828 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2149
timestamp 1710899220
transform 1 0 1788 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2150
timestamp 1710899220
transform 1 0 1372 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2151
timestamp 1710899220
transform 1 0 1252 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2152
timestamp 1710899220
transform 1 0 1372 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2153
timestamp 1710899220
transform 1 0 1284 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2154
timestamp 1710899220
transform 1 0 1628 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2155
timestamp 1710899220
transform 1 0 1588 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2156
timestamp 1710899220
transform 1 0 1452 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2157
timestamp 1710899220
transform 1 0 1452 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2158
timestamp 1710899220
transform 1 0 2180 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2159
timestamp 1710899220
transform 1 0 2148 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2160
timestamp 1710899220
transform 1 0 1372 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2161
timestamp 1710899220
transform 1 0 1356 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2162
timestamp 1710899220
transform 1 0 1396 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2163
timestamp 1710899220
transform 1 0 1364 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2164
timestamp 1710899220
transform 1 0 1364 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2165
timestamp 1710899220
transform 1 0 1340 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2166
timestamp 1710899220
transform 1 0 1348 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2167
timestamp 1710899220
transform 1 0 1284 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2168
timestamp 1710899220
transform 1 0 1412 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2169
timestamp 1710899220
transform 1 0 1372 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2170
timestamp 1710899220
transform 1 0 1428 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2171
timestamp 1710899220
transform 1 0 1340 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2172
timestamp 1710899220
transform 1 0 1452 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2173
timestamp 1710899220
transform 1 0 1316 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2174
timestamp 1710899220
transform 1 0 1380 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2175
timestamp 1710899220
transform 1 0 1356 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2176
timestamp 1710899220
transform 1 0 1428 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2177
timestamp 1710899220
transform 1 0 1372 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2178
timestamp 1710899220
transform 1 0 1404 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2179
timestamp 1710899220
transform 1 0 1340 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2180
timestamp 1710899220
transform 1 0 1212 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2181
timestamp 1710899220
transform 1 0 1196 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2182
timestamp 1710899220
transform 1 0 756 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2183
timestamp 1710899220
transform 1 0 740 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2184
timestamp 1710899220
transform 1 0 684 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2185
timestamp 1710899220
transform 1 0 668 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2186
timestamp 1710899220
transform 1 0 708 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2187
timestamp 1710899220
transform 1 0 644 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2188
timestamp 1710899220
transform 1 0 876 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2189
timestamp 1710899220
transform 1 0 860 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2190
timestamp 1710899220
transform 1 0 724 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2191
timestamp 1710899220
transform 1 0 684 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2192
timestamp 1710899220
transform 1 0 780 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2193
timestamp 1710899220
transform 1 0 660 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2194
timestamp 1710899220
transform 1 0 756 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2195
timestamp 1710899220
transform 1 0 708 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2196
timestamp 1710899220
transform 1 0 700 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2197
timestamp 1710899220
transform 1 0 700 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2198
timestamp 1710899220
transform 1 0 532 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2199
timestamp 1710899220
transform 1 0 524 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2200
timestamp 1710899220
transform 1 0 260 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2201
timestamp 1710899220
transform 1 0 172 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2202
timestamp 1710899220
transform 1 0 276 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_2203
timestamp 1710899220
transform 1 0 212 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2204
timestamp 1710899220
transform 1 0 164 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2205
timestamp 1710899220
transform 1 0 124 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2206
timestamp 1710899220
transform 1 0 404 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2207
timestamp 1710899220
transform 1 0 404 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_2208
timestamp 1710899220
transform 1 0 340 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2209
timestamp 1710899220
transform 1 0 324 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2210
timestamp 1710899220
transform 1 0 308 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2211
timestamp 1710899220
transform 1 0 308 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2212
timestamp 1710899220
transform 1 0 308 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2213
timestamp 1710899220
transform 1 0 300 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2214
timestamp 1710899220
transform 1 0 260 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2215
timestamp 1710899220
transform 1 0 268 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_2216
timestamp 1710899220
transform 1 0 212 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2217
timestamp 1710899220
transform 1 0 188 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2218
timestamp 1710899220
transform 1 0 284 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_2219
timestamp 1710899220
transform 1 0 260 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2220
timestamp 1710899220
transform 1 0 204 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2221
timestamp 1710899220
transform 1 0 756 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2222
timestamp 1710899220
transform 1 0 716 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2223
timestamp 1710899220
transform 1 0 644 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2224
timestamp 1710899220
transform 1 0 620 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2225
timestamp 1710899220
transform 1 0 620 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2226
timestamp 1710899220
transform 1 0 820 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_2227
timestamp 1710899220
transform 1 0 812 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2228
timestamp 1710899220
transform 1 0 812 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2229
timestamp 1710899220
transform 1 0 716 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2230
timestamp 1710899220
transform 1 0 1164 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2231
timestamp 1710899220
transform 1 0 1140 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2232
timestamp 1710899220
transform 1 0 1460 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2233
timestamp 1710899220
transform 1 0 1428 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2234
timestamp 1710899220
transform 1 0 1396 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2235
timestamp 1710899220
transform 1 0 1300 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2236
timestamp 1710899220
transform 1 0 1116 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2237
timestamp 1710899220
transform 1 0 1580 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2238
timestamp 1710899220
transform 1 0 1444 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2239
timestamp 1710899220
transform 1 0 1428 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2240
timestamp 1710899220
transform 1 0 1412 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2241
timestamp 1710899220
transform 1 0 1156 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2242
timestamp 1710899220
transform 1 0 1652 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2243
timestamp 1710899220
transform 1 0 1444 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2244
timestamp 1710899220
transform 1 0 1412 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2245
timestamp 1710899220
transform 1 0 1076 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2246
timestamp 1710899220
transform 1 0 1588 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2247
timestamp 1710899220
transform 1 0 1572 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2248
timestamp 1710899220
transform 1 0 1548 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2249
timestamp 1710899220
transform 1 0 1548 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2250
timestamp 1710899220
transform 1 0 1604 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2251
timestamp 1710899220
transform 1 0 1484 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2252
timestamp 1710899220
transform 1 0 2340 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2253
timestamp 1710899220
transform 1 0 2276 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2254
timestamp 1710899220
transform 1 0 2244 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2255
timestamp 1710899220
transform 1 0 2140 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2256
timestamp 1710899220
transform 1 0 2236 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2257
timestamp 1710899220
transform 1 0 2164 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2258
timestamp 1710899220
transform 1 0 2148 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2259
timestamp 1710899220
transform 1 0 2108 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2260
timestamp 1710899220
transform 1 0 2036 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2261
timestamp 1710899220
transform 1 0 1932 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2262
timestamp 1710899220
transform 1 0 2004 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2263
timestamp 1710899220
transform 1 0 1892 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2264
timestamp 1710899220
transform 1 0 2036 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2265
timestamp 1710899220
transform 1 0 1932 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2266
timestamp 1710899220
transform 1 0 2036 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2267
timestamp 1710899220
transform 1 0 1932 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2268
timestamp 1710899220
transform 1 0 2052 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_2269
timestamp 1710899220
transform 1 0 1948 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2270
timestamp 1710899220
transform 1 0 2132 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2271
timestamp 1710899220
transform 1 0 2004 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2272
timestamp 1710899220
transform 1 0 2468 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2273
timestamp 1710899220
transform 1 0 2364 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2274
timestamp 1710899220
transform 1 0 2428 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2275
timestamp 1710899220
transform 1 0 2324 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2276
timestamp 1710899220
transform 1 0 2444 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2277
timestamp 1710899220
transform 1 0 2340 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2278
timestamp 1710899220
transform 1 0 2444 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2279
timestamp 1710899220
transform 1 0 2340 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2280
timestamp 1710899220
transform 1 0 2412 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2281
timestamp 1710899220
transform 1 0 2292 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2282
timestamp 1710899220
transform 1 0 2436 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2283
timestamp 1710899220
transform 1 0 2316 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2284
timestamp 1710899220
transform 1 0 2564 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2285
timestamp 1710899220
transform 1 0 2508 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2286
timestamp 1710899220
transform 1 0 2644 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2287
timestamp 1710899220
transform 1 0 2580 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2288
timestamp 1710899220
transform 1 0 1460 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2289
timestamp 1710899220
transform 1 0 1276 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2290
timestamp 1710899220
transform 1 0 1452 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2291
timestamp 1710899220
transform 1 0 1364 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2292
timestamp 1710899220
transform 1 0 1780 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2293
timestamp 1710899220
transform 1 0 1276 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2294
timestamp 1710899220
transform 1 0 1556 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2295
timestamp 1710899220
transform 1 0 1492 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2296
timestamp 1710899220
transform 1 0 1628 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2297
timestamp 1710899220
transform 1 0 1556 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2298
timestamp 1710899220
transform 1 0 1540 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2299
timestamp 1710899220
transform 1 0 1532 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2300
timestamp 1710899220
transform 1 0 1372 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2301
timestamp 1710899220
transform 1 0 1612 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2302
timestamp 1710899220
transform 1 0 1556 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2303
timestamp 1710899220
transform 1 0 1476 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2304
timestamp 1710899220
transform 1 0 1452 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2305
timestamp 1710899220
transform 1 0 1276 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2306
timestamp 1710899220
transform 1 0 1452 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2307
timestamp 1710899220
transform 1 0 1364 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2308
timestamp 1710899220
transform 1 0 2156 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2309
timestamp 1710899220
transform 1 0 2012 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2310
timestamp 1710899220
transform 1 0 1996 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2311
timestamp 1710899220
transform 1 0 1988 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2312
timestamp 1710899220
transform 1 0 1916 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2313
timestamp 1710899220
transform 1 0 1884 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2314
timestamp 1710899220
transform 1 0 1692 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2315
timestamp 1710899220
transform 1 0 1692 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2316
timestamp 1710899220
transform 1 0 1660 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2317
timestamp 1710899220
transform 1 0 1124 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2318
timestamp 1710899220
transform 1 0 540 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2319
timestamp 1710899220
transform 1 0 380 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2320
timestamp 1710899220
transform 1 0 372 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2321
timestamp 1710899220
transform 1 0 2252 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2322
timestamp 1710899220
transform 1 0 2188 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2323
timestamp 1710899220
transform 1 0 2188 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2324
timestamp 1710899220
transform 1 0 2172 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2325
timestamp 1710899220
transform 1 0 2284 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2326
timestamp 1710899220
transform 1 0 2164 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2327
timestamp 1710899220
transform 1 0 2164 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2328
timestamp 1710899220
transform 1 0 2204 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2329
timestamp 1710899220
transform 1 0 2132 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2330
timestamp 1710899220
transform 1 0 2108 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2331
timestamp 1710899220
transform 1 0 2260 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2332
timestamp 1710899220
transform 1 0 2260 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_2333
timestamp 1710899220
transform 1 0 2268 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_2334
timestamp 1710899220
transform 1 0 2220 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2335
timestamp 1710899220
transform 1 0 1812 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2336
timestamp 1710899220
transform 1 0 1812 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2337
timestamp 1710899220
transform 1 0 1788 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2338
timestamp 1710899220
transform 1 0 1844 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2339
timestamp 1710899220
transform 1 0 1836 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_2340
timestamp 1710899220
transform 1 0 2012 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2341
timestamp 1710899220
transform 1 0 2012 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2342
timestamp 1710899220
transform 1 0 1868 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2343
timestamp 1710899220
transform 1 0 1852 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2344
timestamp 1710899220
transform 1 0 1844 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2345
timestamp 1710899220
transform 1 0 1828 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2346
timestamp 1710899220
transform 1 0 1756 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2347
timestamp 1710899220
transform 1 0 1724 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2348
timestamp 1710899220
transform 1 0 1980 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2349
timestamp 1710899220
transform 1 0 1972 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2350
timestamp 1710899220
transform 1 0 1940 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2351
timestamp 1710899220
transform 1 0 1772 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2352
timestamp 1710899220
transform 1 0 1772 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2353
timestamp 1710899220
transform 1 0 1684 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2354
timestamp 1710899220
transform 1 0 1732 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2355
timestamp 1710899220
transform 1 0 1692 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2356
timestamp 1710899220
transform 1 0 1524 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2357
timestamp 1710899220
transform 1 0 1716 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2358
timestamp 1710899220
transform 1 0 1580 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2359
timestamp 1710899220
transform 1 0 1980 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2360
timestamp 1710899220
transform 1 0 1804 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2361
timestamp 1710899220
transform 1 0 1716 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2362
timestamp 1710899220
transform 1 0 1732 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2363
timestamp 1710899220
transform 1 0 1540 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2364
timestamp 1710899220
transform 1 0 1548 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2365
timestamp 1710899220
transform 1 0 1540 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2366
timestamp 1710899220
transform 1 0 1516 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2367
timestamp 1710899220
transform 1 0 1420 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2368
timestamp 1710899220
transform 1 0 1284 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2369
timestamp 1710899220
transform 1 0 1524 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_2370
timestamp 1710899220
transform 1 0 1484 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2371
timestamp 1710899220
transform 1 0 1468 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_2372
timestamp 1710899220
transform 1 0 1404 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2373
timestamp 1710899220
transform 1 0 1372 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_2374
timestamp 1710899220
transform 1 0 1500 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_2375
timestamp 1710899220
transform 1 0 1492 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2376
timestamp 1710899220
transform 1 0 1444 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2377
timestamp 1710899220
transform 1 0 1764 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2378
timestamp 1710899220
transform 1 0 1716 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_2379
timestamp 1710899220
transform 1 0 1532 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2380
timestamp 1710899220
transform 1 0 1484 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2381
timestamp 1710899220
transform 1 0 1508 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_2382
timestamp 1710899220
transform 1 0 1396 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2383
timestamp 1710899220
transform 1 0 1412 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2384
timestamp 1710899220
transform 1 0 1388 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2385
timestamp 1710899220
transform 1 0 1060 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2386
timestamp 1710899220
transform 1 0 1372 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_2387
timestamp 1710899220
transform 1 0 1364 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2388
timestamp 1710899220
transform 1 0 1420 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_2389
timestamp 1710899220
transform 1 0 1404 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2390
timestamp 1710899220
transform 1 0 1068 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2391
timestamp 1710899220
transform 1 0 1052 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_2392
timestamp 1710899220
transform 1 0 1788 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2393
timestamp 1710899220
transform 1 0 1740 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2394
timestamp 1710899220
transform 1 0 1260 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2395
timestamp 1710899220
transform 1 0 1244 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2396
timestamp 1710899220
transform 1 0 1268 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2397
timestamp 1710899220
transform 1 0 1236 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2398
timestamp 1710899220
transform 1 0 1812 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2399
timestamp 1710899220
transform 1 0 1228 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_2400
timestamp 1710899220
transform 1 0 1252 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2401
timestamp 1710899220
transform 1 0 580 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2402
timestamp 1710899220
transform 1 0 1244 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_2403
timestamp 1710899220
transform 1 0 884 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2404
timestamp 1710899220
transform 1 0 1292 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2405
timestamp 1710899220
transform 1 0 1260 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2406
timestamp 1710899220
transform 1 0 2660 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2407
timestamp 1710899220
transform 1 0 2596 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2408
timestamp 1710899220
transform 1 0 2540 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2409
timestamp 1710899220
transform 1 0 2524 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2410
timestamp 1710899220
transform 1 0 2476 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2411
timestamp 1710899220
transform 1 0 2452 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2412
timestamp 1710899220
transform 1 0 2332 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2413
timestamp 1710899220
transform 1 0 2300 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2414
timestamp 1710899220
transform 1 0 2324 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2415
timestamp 1710899220
transform 1 0 2308 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2416
timestamp 1710899220
transform 1 0 2524 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2417
timestamp 1710899220
transform 1 0 2508 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2418
timestamp 1710899220
transform 1 0 2644 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2419
timestamp 1710899220
transform 1 0 2628 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2420
timestamp 1710899220
transform 1 0 2556 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2421
timestamp 1710899220
transform 1 0 2556 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2422
timestamp 1710899220
transform 1 0 2356 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2423
timestamp 1710899220
transform 1 0 2324 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2424
timestamp 1710899220
transform 1 0 2356 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2425
timestamp 1710899220
transform 1 0 2324 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2426
timestamp 1710899220
transform 1 0 2660 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2427
timestamp 1710899220
transform 1 0 2556 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2428
timestamp 1710899220
transform 1 0 2548 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2429
timestamp 1710899220
transform 1 0 2524 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2430
timestamp 1710899220
transform 1 0 2556 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2431
timestamp 1710899220
transform 1 0 2540 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2432
timestamp 1710899220
transform 1 0 2660 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2433
timestamp 1710899220
transform 1 0 2540 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2434
timestamp 1710899220
transform 1 0 2348 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2435
timestamp 1710899220
transform 1 0 2340 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2436
timestamp 1710899220
transform 1 0 2556 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2437
timestamp 1710899220
transform 1 0 2540 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2438
timestamp 1710899220
transform 1 0 2596 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2439
timestamp 1710899220
transform 1 0 2580 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2440
timestamp 1710899220
transform 1 0 2396 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2441
timestamp 1710899220
transform 1 0 2380 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2442
timestamp 1710899220
transform 1 0 2316 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2443
timestamp 1710899220
transform 1 0 2300 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2444
timestamp 1710899220
transform 1 0 2284 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2445
timestamp 1710899220
transform 1 0 2268 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2446
timestamp 1710899220
transform 1 0 2036 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2447
timestamp 1710899220
transform 1 0 2020 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2448
timestamp 1710899220
transform 1 0 2180 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2449
timestamp 1710899220
transform 1 0 2164 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2450
timestamp 1710899220
transform 1 0 1964 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2451
timestamp 1710899220
transform 1 0 1932 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2452
timestamp 1710899220
transform 1 0 1948 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2453
timestamp 1710899220
transform 1 0 1916 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2454
timestamp 1710899220
transform 1 0 1948 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2455
timestamp 1710899220
transform 1 0 1916 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2456
timestamp 1710899220
transform 1 0 1908 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2457
timestamp 1710899220
transform 1 0 1876 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2458
timestamp 1710899220
transform 1 0 1948 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2459
timestamp 1710899220
transform 1 0 1916 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2460
timestamp 1710899220
transform 1 0 2124 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2461
timestamp 1710899220
transform 1 0 2092 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2462
timestamp 1710899220
transform 1 0 2196 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2463
timestamp 1710899220
transform 1 0 2180 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2464
timestamp 1710899220
transform 1 0 2156 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2465
timestamp 1710899220
transform 1 0 2124 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2466
timestamp 1710899220
transform 1 0 2308 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2467
timestamp 1710899220
transform 1 0 2292 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2468
timestamp 1710899220
transform 1 0 2284 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2469
timestamp 1710899220
transform 1 0 2252 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2470
timestamp 1710899220
transform 1 0 2060 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2471
timestamp 1710899220
transform 1 0 2036 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2472
timestamp 1710899220
transform 1 0 1964 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2473
timestamp 1710899220
transform 1 0 1956 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2474
timestamp 1710899220
transform 1 0 1948 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2475
timestamp 1710899220
transform 1 0 1756 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2476
timestamp 1710899220
transform 1 0 1724 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2477
timestamp 1710899220
transform 1 0 2036 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_2478
timestamp 1710899220
transform 1 0 2012 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2479
timestamp 1710899220
transform 1 0 1708 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_2480
timestamp 1710899220
transform 1 0 1636 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2481
timestamp 1710899220
transform 1 0 1724 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2482
timestamp 1710899220
transform 1 0 1700 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2483
timestamp 1710899220
transform 1 0 1692 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_2484
timestamp 1710899220
transform 1 0 1668 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_2485
timestamp 1710899220
transform 1 0 1676 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2486
timestamp 1710899220
transform 1 0 1636 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_2487
timestamp 1710899220
transform 1 0 1500 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2488
timestamp 1710899220
transform 1 0 1692 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2489
timestamp 1710899220
transform 1 0 1676 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2490
timestamp 1710899220
transform 1 0 596 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2491
timestamp 1710899220
transform 1 0 1812 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2492
timestamp 1710899220
transform 1 0 1652 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2493
timestamp 1710899220
transform 1 0 1612 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2494
timestamp 1710899220
transform 1 0 1628 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_2495
timestamp 1710899220
transform 1 0 1628 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_2496
timestamp 1710899220
transform 1 0 1796 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_2497
timestamp 1710899220
transform 1 0 1612 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_2498
timestamp 1710899220
transform 1 0 1068 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2499
timestamp 1710899220
transform 1 0 1628 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2500
timestamp 1710899220
transform 1 0 1572 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_2501
timestamp 1710899220
transform 1 0 772 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2502
timestamp 1710899220
transform 1 0 1596 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2503
timestamp 1710899220
transform 1 0 1044 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2504
timestamp 1710899220
transform 1 0 1660 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2505
timestamp 1710899220
transform 1 0 1076 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2506
timestamp 1710899220
transform 1 0 1668 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2507
timestamp 1710899220
transform 1 0 844 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2508
timestamp 1710899220
transform 1 0 1692 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2509
timestamp 1710899220
transform 1 0 1676 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_2510
timestamp 1710899220
transform 1 0 1740 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2511
timestamp 1710899220
transform 1 0 1692 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_2512
timestamp 1710899220
transform 1 0 1788 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2513
timestamp 1710899220
transform 1 0 1708 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2514
timestamp 1710899220
transform 1 0 1796 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2515
timestamp 1710899220
transform 1 0 1772 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2516
timestamp 1710899220
transform 1 0 1908 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2517
timestamp 1710899220
transform 1 0 1772 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2518
timestamp 1710899220
transform 1 0 1764 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_2519
timestamp 1710899220
transform 1 0 1756 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2520
timestamp 1710899220
transform 1 0 1740 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_2521
timestamp 1710899220
transform 1 0 1668 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2522
timestamp 1710899220
transform 1 0 1756 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2523
timestamp 1710899220
transform 1 0 1732 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2524
timestamp 1710899220
transform 1 0 580 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2525
timestamp 1710899220
transform 1 0 564 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2526
timestamp 1710899220
transform 1 0 604 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2527
timestamp 1710899220
transform 1 0 452 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2528
timestamp 1710899220
transform 1 0 1868 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2529
timestamp 1710899220
transform 1 0 1828 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2530
timestamp 1710899220
transform 1 0 1868 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2531
timestamp 1710899220
transform 1 0 1868 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2532
timestamp 1710899220
transform 1 0 1524 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2533
timestamp 1710899220
transform 1 0 1500 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2534
timestamp 1710899220
transform 1 0 1644 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_2535
timestamp 1710899220
transform 1 0 1580 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2536
timestamp 1710899220
transform 1 0 1036 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2537
timestamp 1710899220
transform 1 0 884 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2538
timestamp 1710899220
transform 1 0 772 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2539
timestamp 1710899220
transform 1 0 724 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2540
timestamp 1710899220
transform 1 0 1812 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_2541
timestamp 1710899220
transform 1 0 1804 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2542
timestamp 1710899220
transform 1 0 1668 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2543
timestamp 1710899220
transform 1 0 1580 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2544
timestamp 1710899220
transform 1 0 1956 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2545
timestamp 1710899220
transform 1 0 1908 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_2546
timestamp 1710899220
transform 1 0 1996 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2547
timestamp 1710899220
transform 1 0 1932 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2548
timestamp 1710899220
transform 1 0 1996 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2549
timestamp 1710899220
transform 1 0 1980 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2550
timestamp 1710899220
transform 1 0 1964 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2551
timestamp 1710899220
transform 1 0 1940 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2552
timestamp 1710899220
transform 1 0 2028 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2553
timestamp 1710899220
transform 1 0 1964 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2554
timestamp 1710899220
transform 1 0 1900 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2555
timestamp 1710899220
transform 1 0 1828 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2556
timestamp 1710899220
transform 1 0 1076 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2557
timestamp 1710899220
transform 1 0 1044 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2558
timestamp 1710899220
transform 1 0 1868 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2559
timestamp 1710899220
transform 1 0 1724 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2560
timestamp 1710899220
transform 1 0 1724 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2561
timestamp 1710899220
transform 1 0 1724 0 1 755
box -2 -2 2 2
use M2_M1  M2_M1_2562
timestamp 1710899220
transform 1 0 1732 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_2563
timestamp 1710899220
transform 1 0 1724 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2564
timestamp 1710899220
transform 1 0 1716 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_2565
timestamp 1710899220
transform 1 0 1708 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2566
timestamp 1710899220
transform 1 0 1740 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2567
timestamp 1710899220
transform 1 0 1644 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2568
timestamp 1710899220
transform 1 0 1644 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2569
timestamp 1710899220
transform 1 0 1572 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2570
timestamp 1710899220
transform 1 0 1692 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2571
timestamp 1710899220
transform 1 0 1652 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2572
timestamp 1710899220
transform 1 0 1684 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_2573
timestamp 1710899220
transform 1 0 1588 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2574
timestamp 1710899220
transform 1 0 1604 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2575
timestamp 1710899220
transform 1 0 1604 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2576
timestamp 1710899220
transform 1 0 1764 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2577
timestamp 1710899220
transform 1 0 1716 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_2578
timestamp 1710899220
transform 1 0 1732 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2579
timestamp 1710899220
transform 1 0 1716 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2580
timestamp 1710899220
transform 1 0 1876 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2581
timestamp 1710899220
transform 1 0 1708 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2582
timestamp 1710899220
transform 1 0 1932 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2583
timestamp 1710899220
transform 1 0 1884 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_2584
timestamp 1710899220
transform 1 0 1900 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2585
timestamp 1710899220
transform 1 0 1900 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2586
timestamp 1710899220
transform 1 0 1932 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2587
timestamp 1710899220
transform 1 0 1916 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2588
timestamp 1710899220
transform 1 0 1948 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2589
timestamp 1710899220
transform 1 0 1940 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2590
timestamp 1710899220
transform 1 0 836 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_2591
timestamp 1710899220
transform 1 0 524 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2592
timestamp 1710899220
transform 1 0 884 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2593
timestamp 1710899220
transform 1 0 852 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2594
timestamp 1710899220
transform 1 0 908 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2595
timestamp 1710899220
transform 1 0 860 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2596
timestamp 1710899220
transform 1 0 948 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2597
timestamp 1710899220
transform 1 0 868 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2598
timestamp 1710899220
transform 1 0 876 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_2599
timestamp 1710899220
transform 1 0 540 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2600
timestamp 1710899220
transform 1 0 540 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_2601
timestamp 1710899220
transform 1 0 396 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2602
timestamp 1710899220
transform 1 0 388 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2603
timestamp 1710899220
transform 1 0 372 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2604
timestamp 1710899220
transform 1 0 388 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2605
timestamp 1710899220
transform 1 0 356 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2606
timestamp 1710899220
transform 1 0 948 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2607
timestamp 1710899220
transform 1 0 932 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2608
timestamp 1710899220
transform 1 0 1004 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2609
timestamp 1710899220
transform 1 0 508 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2610
timestamp 1710899220
transform 1 0 508 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2611
timestamp 1710899220
transform 1 0 476 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2612
timestamp 1710899220
transform 1 0 500 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_2613
timestamp 1710899220
transform 1 0 452 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2614
timestamp 1710899220
transform 1 0 444 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2615
timestamp 1710899220
transform 1 0 444 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2616
timestamp 1710899220
transform 1 0 572 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2617
timestamp 1710899220
transform 1 0 444 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2618
timestamp 1710899220
transform 1 0 420 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2619
timestamp 1710899220
transform 1 0 412 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2620
timestamp 1710899220
transform 1 0 1028 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2621
timestamp 1710899220
transform 1 0 988 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2622
timestamp 1710899220
transform 1 0 1052 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2623
timestamp 1710899220
transform 1 0 1020 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2624
timestamp 1710899220
transform 1 0 1060 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_2625
timestamp 1710899220
transform 1 0 636 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2626
timestamp 1710899220
transform 1 0 1076 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2627
timestamp 1710899220
transform 1 0 1052 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2628
timestamp 1710899220
transform 1 0 1036 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2629
timestamp 1710899220
transform 1 0 948 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2630
timestamp 1710899220
transform 1 0 1036 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2631
timestamp 1710899220
transform 1 0 988 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2632
timestamp 1710899220
transform 1 0 1620 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2633
timestamp 1710899220
transform 1 0 1028 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_2634
timestamp 1710899220
transform 1 0 1708 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2635
timestamp 1710899220
transform 1 0 1620 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_2636
timestamp 1710899220
transform 1 0 1788 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2637
timestamp 1710899220
transform 1 0 1692 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2638
timestamp 1710899220
transform 1 0 1740 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2639
timestamp 1710899220
transform 1 0 1708 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2640
timestamp 1710899220
transform 1 0 1100 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2641
timestamp 1710899220
transform 1 0 972 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2642
timestamp 1710899220
transform 1 0 612 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2643
timestamp 1710899220
transform 1 0 412 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2644
timestamp 1710899220
transform 1 0 620 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2645
timestamp 1710899220
transform 1 0 540 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2646
timestamp 1710899220
transform 1 0 804 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2647
timestamp 1710899220
transform 1 0 628 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_2648
timestamp 1710899220
transform 1 0 932 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2649
timestamp 1710899220
transform 1 0 772 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2650
timestamp 1710899220
transform 1 0 804 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_2651
timestamp 1710899220
transform 1 0 780 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2652
timestamp 1710899220
transform 1 0 772 0 1 695
box -2 -2 2 2
use M2_M1  M2_M1_2653
timestamp 1710899220
transform 1 0 772 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2654
timestamp 1710899220
transform 1 0 652 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2655
timestamp 1710899220
transform 1 0 524 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2656
timestamp 1710899220
transform 1 0 1860 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2657
timestamp 1710899220
transform 1 0 1836 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2658
timestamp 1710899220
transform 1 0 724 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2659
timestamp 1710899220
transform 1 0 684 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2660
timestamp 1710899220
transform 1 0 1732 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2661
timestamp 1710899220
transform 1 0 1524 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2662
timestamp 1710899220
transform 1 0 1436 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2663
timestamp 1710899220
transform 1 0 1276 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2664
timestamp 1710899220
transform 1 0 1452 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2665
timestamp 1710899220
transform 1 0 1332 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2666
timestamp 1710899220
transform 1 0 1324 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2667
timestamp 1710899220
transform 1 0 1300 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2668
timestamp 1710899220
transform 1 0 1260 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2669
timestamp 1710899220
transform 1 0 1252 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2670
timestamp 1710899220
transform 1 0 1820 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2671
timestamp 1710899220
transform 1 0 1404 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2672
timestamp 1710899220
transform 1 0 1780 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2673
timestamp 1710899220
transform 1 0 1428 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2674
timestamp 1710899220
transform 1 0 1548 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2675
timestamp 1710899220
transform 1 0 1396 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2676
timestamp 1710899220
transform 1 0 1420 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2677
timestamp 1710899220
transform 1 0 1364 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2678
timestamp 1710899220
transform 1 0 1420 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2679
timestamp 1710899220
transform 1 0 1372 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2680
timestamp 1710899220
transform 1 0 1780 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2681
timestamp 1710899220
transform 1 0 1420 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2682
timestamp 1710899220
transform 1 0 1836 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2683
timestamp 1710899220
transform 1 0 1436 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2684
timestamp 1710899220
transform 1 0 1788 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2685
timestamp 1710899220
transform 1 0 1484 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2686
timestamp 1710899220
transform 1 0 1388 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2687
timestamp 1710899220
transform 1 0 1388 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2688
timestamp 1710899220
transform 1 0 1508 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2689
timestamp 1710899220
transform 1 0 1460 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2690
timestamp 1710899220
transform 1 0 1452 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2691
timestamp 1710899220
transform 1 0 1420 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2692
timestamp 1710899220
transform 1 0 1332 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2693
timestamp 1710899220
transform 1 0 1292 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2694
timestamp 1710899220
transform 1 0 916 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2695
timestamp 1710899220
transform 1 0 820 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2696
timestamp 1710899220
transform 1 0 828 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2697
timestamp 1710899220
transform 1 0 764 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2698
timestamp 1710899220
transform 1 0 676 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2699
timestamp 1710899220
transform 1 0 676 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2700
timestamp 1710899220
transform 1 0 644 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2701
timestamp 1710899220
transform 1 0 644 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2702
timestamp 1710899220
transform 1 0 996 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2703
timestamp 1710899220
transform 1 0 988 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2704
timestamp 1710899220
transform 1 0 1116 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2705
timestamp 1710899220
transform 1 0 1116 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2706
timestamp 1710899220
transform 1 0 684 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2707
timestamp 1710899220
transform 1 0 564 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2708
timestamp 1710899220
transform 1 0 628 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2709
timestamp 1710899220
transform 1 0 540 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2710
timestamp 1710899220
transform 1 0 708 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2711
timestamp 1710899220
transform 1 0 660 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2712
timestamp 1710899220
transform 1 0 2116 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2713
timestamp 1710899220
transform 1 0 1748 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2714
timestamp 1710899220
transform 1 0 1284 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2715
timestamp 1710899220
transform 1 0 2164 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2716
timestamp 1710899220
transform 1 0 1972 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2717
timestamp 1710899220
transform 1 0 1500 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2718
timestamp 1710899220
transform 1 0 1372 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2719
timestamp 1710899220
transform 1 0 1348 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2720
timestamp 1710899220
transform 1 0 1196 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2721
timestamp 1710899220
transform 1 0 1196 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2722
timestamp 1710899220
transform 1 0 1516 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2723
timestamp 1710899220
transform 1 0 1436 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2724
timestamp 1710899220
transform 1 0 1412 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2725
timestamp 1710899220
transform 1 0 1412 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2726
timestamp 1710899220
transform 1 0 1356 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2727
timestamp 1710899220
transform 1 0 1260 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2728
timestamp 1710899220
transform 1 0 1300 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2729
timestamp 1710899220
transform 1 0 1300 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2730
timestamp 1710899220
transform 1 0 1268 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2731
timestamp 1710899220
transform 1 0 1268 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2732
timestamp 1710899220
transform 1 0 196 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2733
timestamp 1710899220
transform 1 0 1460 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2734
timestamp 1710899220
transform 1 0 1380 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2735
timestamp 1710899220
transform 1 0 1292 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2736
timestamp 1710899220
transform 1 0 1252 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2737
timestamp 1710899220
transform 1 0 1004 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2738
timestamp 1710899220
transform 1 0 1292 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2739
timestamp 1710899220
transform 1 0 1292 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2740
timestamp 1710899220
transform 1 0 1284 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2741
timestamp 1710899220
transform 1 0 1236 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2742
timestamp 1710899220
transform 1 0 172 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2743
timestamp 1710899220
transform 1 0 1732 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2744
timestamp 1710899220
transform 1 0 1708 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2745
timestamp 1710899220
transform 1 0 1284 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2746
timestamp 1710899220
transform 1 0 1268 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2747
timestamp 1710899220
transform 1 0 1228 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2748
timestamp 1710899220
transform 1 0 1108 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2749
timestamp 1710899220
transform 1 0 252 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2750
timestamp 1710899220
transform 1 0 1284 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2751
timestamp 1710899220
transform 1 0 1188 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2752
timestamp 1710899220
transform 1 0 1172 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2753
timestamp 1710899220
transform 1 0 1668 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2754
timestamp 1710899220
transform 1 0 1596 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2755
timestamp 1710899220
transform 1 0 1220 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2756
timestamp 1710899220
transform 1 0 1716 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2757
timestamp 1710899220
transform 1 0 1660 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2758
timestamp 1710899220
transform 1 0 1628 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2759
timestamp 1710899220
transform 1 0 1516 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2760
timestamp 1710899220
transform 1 0 1516 0 1 1245
box -2 -2 2 2
use M2_M1  M2_M1_2761
timestamp 1710899220
transform 1 0 1508 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2762
timestamp 1710899220
transform 1 0 1436 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2763
timestamp 1710899220
transform 1 0 1596 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2764
timestamp 1710899220
transform 1 0 1420 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2765
timestamp 1710899220
transform 1 0 1348 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2766
timestamp 1710899220
transform 1 0 1252 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2767
timestamp 1710899220
transform 1 0 1236 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2768
timestamp 1710899220
transform 1 0 1532 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2769
timestamp 1710899220
transform 1 0 1484 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2770
timestamp 1710899220
transform 1 0 1412 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2771
timestamp 1710899220
transform 1 0 1388 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2772
timestamp 1710899220
transform 1 0 1356 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2773
timestamp 1710899220
transform 1 0 1092 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2774
timestamp 1710899220
transform 1 0 924 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2775
timestamp 1710899220
transform 1 0 908 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2776
timestamp 1710899220
transform 1 0 844 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2777
timestamp 1710899220
transform 1 0 828 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2778
timestamp 1710899220
transform 1 0 812 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2779
timestamp 1710899220
transform 1 0 812 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2780
timestamp 1710899220
transform 1 0 788 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2781
timestamp 1710899220
transform 1 0 860 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2782
timestamp 1710899220
transform 1 0 836 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2783
timestamp 1710899220
transform 1 0 956 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2784
timestamp 1710899220
transform 1 0 844 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2785
timestamp 1710899220
transform 1 0 908 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2786
timestamp 1710899220
transform 1 0 884 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2787
timestamp 1710899220
transform 1 0 796 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2788
timestamp 1710899220
transform 1 0 772 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2789
timestamp 1710899220
transform 1 0 1100 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2790
timestamp 1710899220
transform 1 0 1036 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2791
timestamp 1710899220
transform 1 0 948 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2792
timestamp 1710899220
transform 1 0 948 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2793
timestamp 1710899220
transform 1 0 1116 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2794
timestamp 1710899220
transform 1 0 1060 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2795
timestamp 1710899220
transform 1 0 988 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2796
timestamp 1710899220
transform 1 0 964 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2797
timestamp 1710899220
transform 1 0 1148 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2798
timestamp 1710899220
transform 1 0 1108 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2799
timestamp 1710899220
transform 1 0 884 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2800
timestamp 1710899220
transform 1 0 1172 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2801
timestamp 1710899220
transform 1 0 988 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2802
timestamp 1710899220
transform 1 0 1004 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2803
timestamp 1710899220
transform 1 0 980 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2804
timestamp 1710899220
transform 1 0 940 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2805
timestamp 1710899220
transform 1 0 996 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2806
timestamp 1710899220
transform 1 0 996 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2807
timestamp 1710899220
transform 1 0 1124 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2808
timestamp 1710899220
transform 1 0 1012 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2809
timestamp 1710899220
transform 1 0 892 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2810
timestamp 1710899220
transform 1 0 852 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2811
timestamp 1710899220
transform 1 0 876 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2812
timestamp 1710899220
transform 1 0 836 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2813
timestamp 1710899220
transform 1 0 796 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2814
timestamp 1710899220
transform 1 0 852 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_2815
timestamp 1710899220
transform 1 0 788 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2816
timestamp 1710899220
transform 1 0 1004 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2817
timestamp 1710899220
transform 1 0 988 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2818
timestamp 1710899220
transform 1 0 1004 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2819
timestamp 1710899220
transform 1 0 980 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2820
timestamp 1710899220
transform 1 0 1052 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2821
timestamp 1710899220
transform 1 0 988 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2822
timestamp 1710899220
transform 1 0 1084 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2823
timestamp 1710899220
transform 1 0 1068 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2824
timestamp 1710899220
transform 1 0 1028 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2825
timestamp 1710899220
transform 1 0 740 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2826
timestamp 1710899220
transform 1 0 740 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2827
timestamp 1710899220
transform 1 0 732 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2828
timestamp 1710899220
transform 1 0 732 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2829
timestamp 1710899220
transform 1 0 948 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2830
timestamp 1710899220
transform 1 0 780 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_2831
timestamp 1710899220
transform 1 0 780 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2832
timestamp 1710899220
transform 1 0 1036 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2833
timestamp 1710899220
transform 1 0 892 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2834
timestamp 1710899220
transform 1 0 860 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2835
timestamp 1710899220
transform 1 0 804 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2836
timestamp 1710899220
transform 1 0 900 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2837
timestamp 1710899220
transform 1 0 883 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2838
timestamp 1710899220
transform 1 0 860 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2839
timestamp 1710899220
transform 1 0 836 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2840
timestamp 1710899220
transform 1 0 924 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2841
timestamp 1710899220
transform 1 0 876 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2842
timestamp 1710899220
transform 1 0 932 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2843
timestamp 1710899220
transform 1 0 916 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2844
timestamp 1710899220
transform 1 0 812 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2845
timestamp 1710899220
transform 1 0 772 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2846
timestamp 1710899220
transform 1 0 764 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2847
timestamp 1710899220
transform 1 0 756 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2848
timestamp 1710899220
transform 1 0 828 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2849
timestamp 1710899220
transform 1 0 812 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2850
timestamp 1710899220
transform 1 0 756 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2851
timestamp 1710899220
transform 1 0 1132 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2852
timestamp 1710899220
transform 1 0 1108 0 1 1217
box -2 -2 2 2
use M2_M1  M2_M1_2853
timestamp 1710899220
transform 1 0 1036 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2854
timestamp 1710899220
transform 1 0 964 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2855
timestamp 1710899220
transform 1 0 980 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2856
timestamp 1710899220
transform 1 0 964 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_2857
timestamp 1710899220
transform 1 0 924 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2858
timestamp 1710899220
transform 1 0 908 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2859
timestamp 1710899220
transform 1 0 1036 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2860
timestamp 1710899220
transform 1 0 964 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2861
timestamp 1710899220
transform 1 0 1068 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2862
timestamp 1710899220
transform 1 0 1004 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2863
timestamp 1710899220
transform 1 0 972 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2864
timestamp 1710899220
transform 1 0 916 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2865
timestamp 1710899220
transform 1 0 1044 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2866
timestamp 1710899220
transform 1 0 1020 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2867
timestamp 1710899220
transform 1 0 932 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2868
timestamp 1710899220
transform 1 0 844 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_2869
timestamp 1710899220
transform 1 0 844 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2870
timestamp 1710899220
transform 1 0 916 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2871
timestamp 1710899220
transform 1 0 892 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2872
timestamp 1710899220
transform 1 0 876 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2873
timestamp 1710899220
transform 1 0 852 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2874
timestamp 1710899220
transform 1 0 932 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2875
timestamp 1710899220
transform 1 0 876 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2876
timestamp 1710899220
transform 1 0 844 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2877
timestamp 1710899220
transform 1 0 836 0 1 1355
box -2 -2 2 2
use M2_M1  M2_M1_2878
timestamp 1710899220
transform 1 0 788 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2879
timestamp 1710899220
transform 1 0 1052 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2880
timestamp 1710899220
transform 1 0 1004 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2881
timestamp 1710899220
transform 1 0 1020 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2882
timestamp 1710899220
transform 1 0 860 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2883
timestamp 1710899220
transform 1 0 964 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2884
timestamp 1710899220
transform 1 0 948 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2885
timestamp 1710899220
transform 1 0 988 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2886
timestamp 1710899220
transform 1 0 900 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2887
timestamp 1710899220
transform 1 0 868 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2888
timestamp 1710899220
transform 1 0 860 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2889
timestamp 1710899220
transform 1 0 868 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2890
timestamp 1710899220
transform 1 0 804 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2891
timestamp 1710899220
transform 1 0 756 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2892
timestamp 1710899220
transform 1 0 708 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2893
timestamp 1710899220
transform 1 0 764 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2894
timestamp 1710899220
transform 1 0 716 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2895
timestamp 1710899220
transform 1 0 764 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2896
timestamp 1710899220
transform 1 0 700 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2897
timestamp 1710899220
transform 1 0 756 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2898
timestamp 1710899220
transform 1 0 708 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2899
timestamp 1710899220
transform 1 0 884 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2900
timestamp 1710899220
transform 1 0 796 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2901
timestamp 1710899220
transform 1 0 908 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2902
timestamp 1710899220
transform 1 0 876 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2903
timestamp 1710899220
transform 1 0 804 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2904
timestamp 1710899220
transform 1 0 772 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2905
timestamp 1710899220
transform 1 0 788 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2906
timestamp 1710899220
transform 1 0 708 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2907
timestamp 1710899220
transform 1 0 676 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2908
timestamp 1710899220
transform 1 0 532 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2909
timestamp 1710899220
transform 1 0 676 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2910
timestamp 1710899220
transform 1 0 652 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2911
timestamp 1710899220
transform 1 0 684 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2912
timestamp 1710899220
transform 1 0 676 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2913
timestamp 1710899220
transform 1 0 668 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2914
timestamp 1710899220
transform 1 0 644 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2915
timestamp 1710899220
transform 1 0 644 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2916
timestamp 1710899220
transform 1 0 612 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2917
timestamp 1710899220
transform 1 0 588 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2918
timestamp 1710899220
transform 1 0 580 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2919
timestamp 1710899220
transform 1 0 564 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2920
timestamp 1710899220
transform 1 0 564 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2921
timestamp 1710899220
transform 1 0 708 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2922
timestamp 1710899220
transform 1 0 700 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2923
timestamp 1710899220
transform 1 0 684 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2924
timestamp 1710899220
transform 1 0 660 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2925
timestamp 1710899220
transform 1 0 604 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2926
timestamp 1710899220
transform 1 0 596 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2927
timestamp 1710899220
transform 1 0 580 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2928
timestamp 1710899220
transform 1 0 628 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2929
timestamp 1710899220
transform 1 0 628 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2930
timestamp 1710899220
transform 1 0 556 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2931
timestamp 1710899220
transform 1 0 516 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2932
timestamp 1710899220
transform 1 0 516 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2933
timestamp 1710899220
transform 1 0 516 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2934
timestamp 1710899220
transform 1 0 516 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2935
timestamp 1710899220
transform 1 0 660 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2936
timestamp 1710899220
transform 1 0 660 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2937
timestamp 1710899220
transform 1 0 596 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2938
timestamp 1710899220
transform 1 0 540 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2939
timestamp 1710899220
transform 1 0 540 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2940
timestamp 1710899220
transform 1 0 532 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2941
timestamp 1710899220
transform 1 0 524 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2942
timestamp 1710899220
transform 1 0 732 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2943
timestamp 1710899220
transform 1 0 652 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2944
timestamp 1710899220
transform 1 0 724 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2945
timestamp 1710899220
transform 1 0 700 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2946
timestamp 1710899220
transform 1 0 724 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2947
timestamp 1710899220
transform 1 0 636 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2948
timestamp 1710899220
transform 1 0 700 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2949
timestamp 1710899220
transform 1 0 588 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2950
timestamp 1710899220
transform 1 0 700 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2951
timestamp 1710899220
transform 1 0 676 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2952
timestamp 1710899220
transform 1 0 612 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2953
timestamp 1710899220
transform 1 0 532 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2954
timestamp 1710899220
transform 1 0 612 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2955
timestamp 1710899220
transform 1 0 588 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2956
timestamp 1710899220
transform 1 0 788 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2957
timestamp 1710899220
transform 1 0 780 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2958
timestamp 1710899220
transform 1 0 764 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2959
timestamp 1710899220
transform 1 0 628 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2960
timestamp 1710899220
transform 1 0 780 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2961
timestamp 1710899220
transform 1 0 764 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2962
timestamp 1710899220
transform 1 0 716 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2963
timestamp 1710899220
transform 1 0 652 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2964
timestamp 1710899220
transform 1 0 716 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2965
timestamp 1710899220
transform 1 0 692 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2966
timestamp 1710899220
transform 1 0 596 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2967
timestamp 1710899220
transform 1 0 524 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2968
timestamp 1710899220
transform 1 0 596 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2969
timestamp 1710899220
transform 1 0 572 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2970
timestamp 1710899220
transform 1 0 244 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2971
timestamp 1710899220
transform 1 0 212 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2972
timestamp 1710899220
transform 1 0 236 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2973
timestamp 1710899220
transform 1 0 212 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2974
timestamp 1710899220
transform 1 0 324 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2975
timestamp 1710899220
transform 1 0 180 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2976
timestamp 1710899220
transform 1 0 284 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2977
timestamp 1710899220
transform 1 0 188 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2978
timestamp 1710899220
transform 1 0 612 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2979
timestamp 1710899220
transform 1 0 260 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2980
timestamp 1710899220
transform 1 0 396 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2981
timestamp 1710899220
transform 1 0 268 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2982
timestamp 1710899220
transform 1 0 468 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2983
timestamp 1710899220
transform 1 0 372 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2984
timestamp 1710899220
transform 1 0 412 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2985
timestamp 1710899220
transform 1 0 380 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2986
timestamp 1710899220
transform 1 0 588 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2987
timestamp 1710899220
transform 1 0 548 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2988
timestamp 1710899220
transform 1 0 548 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2989
timestamp 1710899220
transform 1 0 452 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2990
timestamp 1710899220
transform 1 0 380 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2991
timestamp 1710899220
transform 1 0 356 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2992
timestamp 1710899220
transform 1 0 348 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2993
timestamp 1710899220
transform 1 0 628 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2994
timestamp 1710899220
transform 1 0 580 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2995
timestamp 1710899220
transform 1 0 572 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2996
timestamp 1710899220
transform 1 0 484 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2997
timestamp 1710899220
transform 1 0 420 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2998
timestamp 1710899220
transform 1 0 380 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2999
timestamp 1710899220
transform 1 0 364 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3000
timestamp 1710899220
transform 1 0 628 0 1 1217
box -2 -2 2 2
use M2_M1  M2_M1_3001
timestamp 1710899220
transform 1 0 604 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3002
timestamp 1710899220
transform 1 0 540 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3003
timestamp 1710899220
transform 1 0 452 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3004
timestamp 1710899220
transform 1 0 436 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3005
timestamp 1710899220
transform 1 0 420 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3006
timestamp 1710899220
transform 1 0 420 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3007
timestamp 1710899220
transform 1 0 644 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3008
timestamp 1710899220
transform 1 0 644 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3009
timestamp 1710899220
transform 1 0 556 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3010
timestamp 1710899220
transform 1 0 500 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3011
timestamp 1710899220
transform 1 0 476 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3012
timestamp 1710899220
transform 1 0 436 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3013
timestamp 1710899220
transform 1 0 436 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3014
timestamp 1710899220
transform 1 0 636 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3015
timestamp 1710899220
transform 1 0 588 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3016
timestamp 1710899220
transform 1 0 620 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3017
timestamp 1710899220
transform 1 0 580 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3018
timestamp 1710899220
transform 1 0 532 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3019
timestamp 1710899220
transform 1 0 292 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3020
timestamp 1710899220
transform 1 0 364 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3021
timestamp 1710899220
transform 1 0 300 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3022
timestamp 1710899220
transform 1 0 428 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3023
timestamp 1710899220
transform 1 0 340 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3024
timestamp 1710899220
transform 1 0 356 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3025
timestamp 1710899220
transform 1 0 348 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3026
timestamp 1710899220
transform 1 0 548 0 1 1204
box -2 -2 2 2
use M2_M1  M2_M1_3027
timestamp 1710899220
transform 1 0 492 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3028
timestamp 1710899220
transform 1 0 564 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3029
timestamp 1710899220
transform 1 0 508 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3030
timestamp 1710899220
transform 1 0 244 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3031
timestamp 1710899220
transform 1 0 228 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3032
timestamp 1710899220
transform 1 0 524 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3033
timestamp 1710899220
transform 1 0 276 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3034
timestamp 1710899220
transform 1 0 332 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3035
timestamp 1710899220
transform 1 0 292 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3036
timestamp 1710899220
transform 1 0 428 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3037
timestamp 1710899220
transform 1 0 300 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3038
timestamp 1710899220
transform 1 0 372 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3039
timestamp 1710899220
transform 1 0 308 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3040
timestamp 1710899220
transform 1 0 500 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3041
timestamp 1710899220
transform 1 0 492 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3042
timestamp 1710899220
transform 1 0 508 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3043
timestamp 1710899220
transform 1 0 476 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3044
timestamp 1710899220
transform 1 0 164 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3045
timestamp 1710899220
transform 1 0 148 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3046
timestamp 1710899220
transform 1 0 212 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3047
timestamp 1710899220
transform 1 0 180 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3048
timestamp 1710899220
transform 1 0 252 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3049
timestamp 1710899220
transform 1 0 188 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3050
timestamp 1710899220
transform 1 0 276 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3051
timestamp 1710899220
transform 1 0 196 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3052
timestamp 1710899220
transform 1 0 308 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3053
timestamp 1710899220
transform 1 0 244 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3054
timestamp 1710899220
transform 1 0 308 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3055
timestamp 1710899220
transform 1 0 252 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3056
timestamp 1710899220
transform 1 0 468 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3057
timestamp 1710899220
transform 1 0 284 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3058
timestamp 1710899220
transform 1 0 364 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3059
timestamp 1710899220
transform 1 0 292 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3060
timestamp 1710899220
transform 1 0 404 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3061
timestamp 1710899220
transform 1 0 404 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3062
timestamp 1710899220
transform 1 0 380 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3063
timestamp 1710899220
transform 1 0 372 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3064
timestamp 1710899220
transform 1 0 356 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3065
timestamp 1710899220
transform 1 0 340 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3066
timestamp 1710899220
transform 1 0 340 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3067
timestamp 1710899220
transform 1 0 324 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3068
timestamp 1710899220
transform 1 0 420 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3069
timestamp 1710899220
transform 1 0 388 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3070
timestamp 1710899220
transform 1 0 380 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3071
timestamp 1710899220
transform 1 0 372 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3072
timestamp 1710899220
transform 1 0 356 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3073
timestamp 1710899220
transform 1 0 348 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3074
timestamp 1710899220
transform 1 0 340 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3075
timestamp 1710899220
transform 1 0 460 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3076
timestamp 1710899220
transform 1 0 460 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3077
timestamp 1710899220
transform 1 0 460 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3078
timestamp 1710899220
transform 1 0 460 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3079
timestamp 1710899220
transform 1 0 444 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3080
timestamp 1710899220
transform 1 0 444 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3081
timestamp 1710899220
transform 1 0 412 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3082
timestamp 1710899220
transform 1 0 412 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3083
timestamp 1710899220
transform 1 0 476 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3084
timestamp 1710899220
transform 1 0 476 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3085
timestamp 1710899220
transform 1 0 476 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3086
timestamp 1710899220
transform 1 0 476 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3087
timestamp 1710899220
transform 1 0 468 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3088
timestamp 1710899220
transform 1 0 428 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3089
timestamp 1710899220
transform 1 0 428 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3090
timestamp 1710899220
transform 1 0 468 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3091
timestamp 1710899220
transform 1 0 284 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3092
timestamp 1710899220
transform 1 0 380 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3093
timestamp 1710899220
transform 1 0 292 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3094
timestamp 1710899220
transform 1 0 308 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3095
timestamp 1710899220
transform 1 0 228 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3096
timestamp 1710899220
transform 1 0 260 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3097
timestamp 1710899220
transform 1 0 236 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3098
timestamp 1710899220
transform 1 0 420 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3099
timestamp 1710899220
transform 1 0 236 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3100
timestamp 1710899220
transform 1 0 348 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3101
timestamp 1710899220
transform 1 0 244 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3102
timestamp 1710899220
transform 1 0 468 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3103
timestamp 1710899220
transform 1 0 284 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3104
timestamp 1710899220
transform 1 0 412 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3105
timestamp 1710899220
transform 1 0 292 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3106
timestamp 1710899220
transform 1 0 132 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3107
timestamp 1710899220
transform 1 0 132 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3108
timestamp 1710899220
transform 1 0 300 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3109
timestamp 1710899220
transform 1 0 188 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3110
timestamp 1710899220
transform 1 0 236 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3111
timestamp 1710899220
transform 1 0 204 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3112
timestamp 1710899220
transform 1 0 420 0 1 1785
box -2 -2 2 2
use M2_M1  M2_M1_3113
timestamp 1710899220
transform 1 0 420 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3114
timestamp 1710899220
transform 1 0 212 0 1 1785
box -2 -2 2 2
use M2_M1  M2_M1_3115
timestamp 1710899220
transform 1 0 212 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3116
timestamp 1710899220
transform 1 0 332 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3117
timestamp 1710899220
transform 1 0 220 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3118
timestamp 1710899220
transform 1 0 460 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3119
timestamp 1710899220
transform 1 0 276 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3120
timestamp 1710899220
transform 1 0 372 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3121
timestamp 1710899220
transform 1 0 284 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3122
timestamp 1710899220
transform 1 0 196 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3123
timestamp 1710899220
transform 1 0 172 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3124
timestamp 1710899220
transform 1 0 228 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3125
timestamp 1710899220
transform 1 0 196 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3126
timestamp 1710899220
transform 1 0 252 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3127
timestamp 1710899220
transform 1 0 204 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3128
timestamp 1710899220
transform 1 0 276 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3129
timestamp 1710899220
transform 1 0 212 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3130
timestamp 1710899220
transform 1 0 532 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3131
timestamp 1710899220
transform 1 0 252 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3132
timestamp 1710899220
transform 1 0 308 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3133
timestamp 1710899220
transform 1 0 260 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3134
timestamp 1710899220
transform 1 0 484 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3135
timestamp 1710899220
transform 1 0 284 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3136
timestamp 1710899220
transform 1 0 404 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3137
timestamp 1710899220
transform 1 0 292 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3138
timestamp 1710899220
transform 1 0 636 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3139
timestamp 1710899220
transform 1 0 636 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3140
timestamp 1710899220
transform 1 0 580 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3141
timestamp 1710899220
transform 1 0 388 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3142
timestamp 1710899220
transform 1 0 364 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3143
timestamp 1710899220
transform 1 0 348 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3144
timestamp 1710899220
transform 1 0 332 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3145
timestamp 1710899220
transform 1 0 676 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3146
timestamp 1710899220
transform 1 0 652 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3147
timestamp 1710899220
transform 1 0 612 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3148
timestamp 1710899220
transform 1 0 412 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3149
timestamp 1710899220
transform 1 0 388 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3150
timestamp 1710899220
transform 1 0 372 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3151
timestamp 1710899220
transform 1 0 348 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3152
timestamp 1710899220
transform 1 0 580 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3153
timestamp 1710899220
transform 1 0 540 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3154
timestamp 1710899220
transform 1 0 532 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3155
timestamp 1710899220
transform 1 0 468 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3156
timestamp 1710899220
transform 1 0 444 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3157
timestamp 1710899220
transform 1 0 436 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3158
timestamp 1710899220
transform 1 0 412 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3159
timestamp 1710899220
transform 1 0 612 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3160
timestamp 1710899220
transform 1 0 564 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3161
timestamp 1710899220
transform 1 0 556 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3162
timestamp 1710899220
transform 1 0 492 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3163
timestamp 1710899220
transform 1 0 468 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3164
timestamp 1710899220
transform 1 0 452 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3165
timestamp 1710899220
transform 1 0 428 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3166
timestamp 1710899220
transform 1 0 556 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3167
timestamp 1710899220
transform 1 0 508 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3168
timestamp 1710899220
transform 1 0 644 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3169
timestamp 1710899220
transform 1 0 508 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3170
timestamp 1710899220
transform 1 0 524 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3171
timestamp 1710899220
transform 1 0 220 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3172
timestamp 1710899220
transform 1 0 340 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3173
timestamp 1710899220
transform 1 0 228 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3174
timestamp 1710899220
transform 1 0 444 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3175
timestamp 1710899220
transform 1 0 308 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3176
timestamp 1710899220
transform 1 0 364 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3177
timestamp 1710899220
transform 1 0 324 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3178
timestamp 1710899220
transform 1 0 548 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3179
timestamp 1710899220
transform 1 0 500 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3180
timestamp 1710899220
transform 1 0 604 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3181
timestamp 1710899220
transform 1 0 508 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3182
timestamp 1710899220
transform 1 0 188 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3183
timestamp 1710899220
transform 1 0 180 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3184
timestamp 1710899220
transform 1 0 260 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3185
timestamp 1710899220
transform 1 0 204 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3186
timestamp 1710899220
transform 1 0 308 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3187
timestamp 1710899220
transform 1 0 228 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3188
timestamp 1710899220
transform 1 0 420 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3189
timestamp 1710899220
transform 1 0 284 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3190
timestamp 1710899220
transform 1 0 340 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3191
timestamp 1710899220
transform 1 0 292 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3192
timestamp 1710899220
transform 1 0 460 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3193
timestamp 1710899220
transform 1 0 236 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3194
timestamp 1710899220
transform 1 0 380 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3195
timestamp 1710899220
transform 1 0 244 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3196
timestamp 1710899220
transform 1 0 2188 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3197
timestamp 1710899220
transform 1 0 2188 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3198
timestamp 1710899220
transform 1 0 2292 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3199
timestamp 1710899220
transform 1 0 2212 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3200
timestamp 1710899220
transform 1 0 1916 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3201
timestamp 1710899220
transform 1 0 1836 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3202
timestamp 1710899220
transform 1 0 1868 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3203
timestamp 1710899220
transform 1 0 1804 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3204
timestamp 1710899220
transform 1 0 1988 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3205
timestamp 1710899220
transform 1 0 1988 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3206
timestamp 1710899220
transform 1 0 700 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3207
timestamp 1710899220
transform 1 0 644 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3208
timestamp 1710899220
transform 1 0 356 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3209
timestamp 1710899220
transform 1 0 292 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3210
timestamp 1710899220
transform 1 0 324 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3211
timestamp 1710899220
transform 1 0 228 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3212
timestamp 1710899220
transform 1 0 292 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3213
timestamp 1710899220
transform 1 0 236 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3214
timestamp 1710899220
transform 1 0 1196 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3215
timestamp 1710899220
transform 1 0 1140 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3216
timestamp 1710899220
transform 1 0 1012 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3217
timestamp 1710899220
transform 1 0 972 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3218
timestamp 1710899220
transform 1 0 852 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3219
timestamp 1710899220
transform 1 0 796 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3220
timestamp 1710899220
transform 1 0 524 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3221
timestamp 1710899220
transform 1 0 500 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3222
timestamp 1710899220
transform 1 0 316 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3223
timestamp 1710899220
transform 1 0 228 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3224
timestamp 1710899220
transform 1 0 364 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3225
timestamp 1710899220
transform 1 0 292 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3226
timestamp 1710899220
transform 1 0 988 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3227
timestamp 1710899220
transform 1 0 988 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3228
timestamp 1710899220
transform 1 0 1108 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3229
timestamp 1710899220
transform 1 0 1108 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3230
timestamp 1710899220
transform 1 0 1180 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3231
timestamp 1710899220
transform 1 0 1164 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3232
timestamp 1710899220
transform 1 0 1748 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3233
timestamp 1710899220
transform 1 0 1676 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3234
timestamp 1710899220
transform 1 0 1596 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3235
timestamp 1710899220
transform 1 0 1596 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3236
timestamp 1710899220
transform 1 0 1700 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3237
timestamp 1710899220
transform 1 0 1676 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3238
timestamp 1710899220
transform 1 0 2076 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3239
timestamp 1710899220
transform 1 0 2004 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3240
timestamp 1710899220
transform 1 0 2068 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3241
timestamp 1710899220
transform 1 0 1996 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3242
timestamp 1710899220
transform 1 0 1980 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3243
timestamp 1710899220
transform 1 0 1972 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3244
timestamp 1710899220
transform 1 0 1644 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3245
timestamp 1710899220
transform 1 0 1612 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3246
timestamp 1710899220
transform 1 0 1828 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3247
timestamp 1710899220
transform 1 0 1724 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3248
timestamp 1710899220
transform 1 0 1940 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3249
timestamp 1710899220
transform 1 0 1868 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3250
timestamp 1710899220
transform 1 0 2044 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3251
timestamp 1710899220
transform 1 0 1972 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3252
timestamp 1710899220
transform 1 0 2068 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3253
timestamp 1710899220
transform 1 0 1980 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3254
timestamp 1710899220
transform 1 0 2092 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3255
timestamp 1710899220
transform 1 0 2020 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3256
timestamp 1710899220
transform 1 0 1492 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3257
timestamp 1710899220
transform 1 0 1452 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3258
timestamp 1710899220
transform 1 0 1996 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3259
timestamp 1710899220
transform 1 0 1836 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3260
timestamp 1710899220
transform 1 0 1868 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3261
timestamp 1710899220
transform 1 0 1788 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3262
timestamp 1710899220
transform 1 0 1588 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3263
timestamp 1710899220
transform 1 0 1548 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3264
timestamp 1710899220
transform 1 0 1460 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3265
timestamp 1710899220
transform 1 0 1420 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3266
timestamp 1710899220
transform 1 0 1460 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3267
timestamp 1710899220
transform 1 0 1420 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3268
timestamp 1710899220
transform 1 0 1876 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3269
timestamp 1710899220
transform 1 0 1780 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3270
timestamp 1710899220
transform 1 0 1884 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3271
timestamp 1710899220
transform 1 0 1836 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3272
timestamp 1710899220
transform 1 0 1804 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3273
timestamp 1710899220
transform 1 0 1788 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3274
timestamp 1710899220
transform 1 0 1388 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3275
timestamp 1710899220
transform 1 0 1388 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3276
timestamp 1710899220
transform 1 0 1548 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3277
timestamp 1710899220
transform 1 0 1508 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3278
timestamp 1710899220
transform 1 0 1492 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3279
timestamp 1710899220
transform 1 0 1452 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3280
timestamp 1710899220
transform 1 0 1332 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3281
timestamp 1710899220
transform 1 0 1316 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3282
timestamp 1710899220
transform 1 0 1188 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3283
timestamp 1710899220
transform 1 0 1124 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3284
timestamp 1710899220
transform 1 0 916 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3285
timestamp 1710899220
transform 1 0 916 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3286
timestamp 1710899220
transform 1 0 828 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3287
timestamp 1710899220
transform 1 0 812 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3288
timestamp 1710899220
transform 1 0 692 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3289
timestamp 1710899220
transform 1 0 676 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3290
timestamp 1710899220
transform 1 0 636 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3291
timestamp 1710899220
transform 1 0 612 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3292
timestamp 1710899220
transform 1 0 852 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3293
timestamp 1710899220
transform 1 0 796 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3294
timestamp 1710899220
transform 1 0 988 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3295
timestamp 1710899220
transform 1 0 900 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3296
timestamp 1710899220
transform 1 0 1188 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3297
timestamp 1710899220
transform 1 0 1116 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3298
timestamp 1710899220
transform 1 0 564 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3299
timestamp 1710899220
transform 1 0 500 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3300
timestamp 1710899220
transform 1 0 540 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3301
timestamp 1710899220
transform 1 0 460 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3302
timestamp 1710899220
transform 1 0 628 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3303
timestamp 1710899220
transform 1 0 604 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3304
timestamp 1710899220
transform 1 0 692 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3305
timestamp 1710899220
transform 1 0 628 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3306
timestamp 1710899220
transform 1 0 1172 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3307
timestamp 1710899220
transform 1 0 1164 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3308
timestamp 1710899220
transform 1 0 1172 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3309
timestamp 1710899220
transform 1 0 1156 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3310
timestamp 1710899220
transform 1 0 1348 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3311
timestamp 1710899220
transform 1 0 1276 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3312
timestamp 1710899220
transform 1 0 1476 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3313
timestamp 1710899220
transform 1 0 1412 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3314
timestamp 1710899220
transform 1 0 1324 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3315
timestamp 1710899220
transform 1 0 1260 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3316
timestamp 1710899220
transform 1 0 2348 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3317
timestamp 1710899220
transform 1 0 2340 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3318
timestamp 1710899220
transform 1 0 2364 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3319
timestamp 1710899220
transform 1 0 2364 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3320
timestamp 1710899220
transform 1 0 2428 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3321
timestamp 1710899220
transform 1 0 2428 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3322
timestamp 1710899220
transform 1 0 2476 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3323
timestamp 1710899220
transform 1 0 2468 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3324
timestamp 1710899220
transform 1 0 2356 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3325
timestamp 1710899220
transform 1 0 2148 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3326
timestamp 1710899220
transform 1 0 2564 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3327
timestamp 1710899220
transform 1 0 2540 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3328
timestamp 1710899220
transform 1 0 2556 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3329
timestamp 1710899220
transform 1 0 2524 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3330
timestamp 1710899220
transform 1 0 2508 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3331
timestamp 1710899220
transform 1 0 2508 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3332
timestamp 1710899220
transform 1 0 2428 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_3333
timestamp 1710899220
transform 1 0 2380 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3334
timestamp 1710899220
transform 1 0 2372 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_3335
timestamp 1710899220
transform 1 0 2620 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3336
timestamp 1710899220
transform 1 0 2556 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3337
timestamp 1710899220
transform 1 0 2548 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3338
timestamp 1710899220
transform 1 0 2324 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3339
timestamp 1710899220
transform 1 0 2212 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3340
timestamp 1710899220
transform 1 0 2308 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3341
timestamp 1710899220
transform 1 0 2260 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3342
timestamp 1710899220
transform 1 0 2252 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3343
timestamp 1710899220
transform 1 0 2276 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3344
timestamp 1710899220
transform 1 0 2252 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3345
timestamp 1710899220
transform 1 0 2204 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3346
timestamp 1710899220
transform 1 0 2492 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3347
timestamp 1710899220
transform 1 0 2284 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3348
timestamp 1710899220
transform 1 0 2284 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_3349
timestamp 1710899220
transform 1 0 2300 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3350
timestamp 1710899220
transform 1 0 2268 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3351
timestamp 1710899220
transform 1 0 2372 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3352
timestamp 1710899220
transform 1 0 2260 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_3353
timestamp 1710899220
transform 1 0 2388 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3354
timestamp 1710899220
transform 1 0 2388 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3355
timestamp 1710899220
transform 1 0 2372 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_3356
timestamp 1710899220
transform 1 0 2332 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3357
timestamp 1710899220
transform 1 0 2444 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3358
timestamp 1710899220
transform 1 0 2364 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3359
timestamp 1710899220
transform 1 0 2244 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3360
timestamp 1710899220
transform 1 0 2364 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3361
timestamp 1710899220
transform 1 0 2316 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3362
timestamp 1710899220
transform 1 0 2380 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3363
timestamp 1710899220
transform 1 0 2364 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_3364
timestamp 1710899220
transform 1 0 2444 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3365
timestamp 1710899220
transform 1 0 2436 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3366
timestamp 1710899220
transform 1 0 2548 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3367
timestamp 1710899220
transform 1 0 2452 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3368
timestamp 1710899220
transform 1 0 2492 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3369
timestamp 1710899220
transform 1 0 2484 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3370
timestamp 1710899220
transform 1 0 2532 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3371
timestamp 1710899220
transform 1 0 2484 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_3372
timestamp 1710899220
transform 1 0 2444 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3373
timestamp 1710899220
transform 1 0 2620 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3374
timestamp 1710899220
transform 1 0 2524 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3375
timestamp 1710899220
transform 1 0 2572 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3376
timestamp 1710899220
transform 1 0 2532 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3377
timestamp 1710899220
transform 1 0 2380 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3378
timestamp 1710899220
transform 1 0 2356 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3379
timestamp 1710899220
transform 1 0 2316 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3380
timestamp 1710899220
transform 1 0 2436 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3381
timestamp 1710899220
transform 1 0 2420 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3382
timestamp 1710899220
transform 1 0 2428 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3383
timestamp 1710899220
transform 1 0 2356 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3384
timestamp 1710899220
transform 1 0 2316 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3385
timestamp 1710899220
transform 1 0 2620 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3386
timestamp 1710899220
transform 1 0 2604 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3387
timestamp 1710899220
transform 1 0 2612 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3388
timestamp 1710899220
transform 1 0 2596 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3389
timestamp 1710899220
transform 1 0 2532 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3390
timestamp 1710899220
transform 1 0 2444 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3391
timestamp 1710899220
transform 1 0 2396 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3392
timestamp 1710899220
transform 1 0 2388 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3393
timestamp 1710899220
transform 1 0 2492 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3394
timestamp 1710899220
transform 1 0 2396 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_3395
timestamp 1710899220
transform 1 0 2564 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3396
timestamp 1710899220
transform 1 0 2476 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3397
timestamp 1710899220
transform 1 0 2492 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3398
timestamp 1710899220
transform 1 0 2436 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3399
timestamp 1710899220
transform 1 0 2364 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3400
timestamp 1710899220
transform 1 0 2324 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3401
timestamp 1710899220
transform 1 0 2300 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3402
timestamp 1710899220
transform 1 0 2356 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3403
timestamp 1710899220
transform 1 0 2324 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3404
timestamp 1710899220
transform 1 0 2380 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3405
timestamp 1710899220
transform 1 0 2324 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3406
timestamp 1710899220
transform 1 0 2644 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3407
timestamp 1710899220
transform 1 0 2524 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_3408
timestamp 1710899220
transform 1 0 2500 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3409
timestamp 1710899220
transform 1 0 2364 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_3410
timestamp 1710899220
transform 1 0 2580 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3411
timestamp 1710899220
transform 1 0 2476 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3412
timestamp 1710899220
transform 1 0 2476 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3413
timestamp 1710899220
transform 1 0 2468 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3414
timestamp 1710899220
transform 1 0 2524 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_3415
timestamp 1710899220
transform 1 0 2524 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3416
timestamp 1710899220
transform 1 0 2636 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3417
timestamp 1710899220
transform 1 0 2540 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3418
timestamp 1710899220
transform 1 0 2612 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_3419
timestamp 1710899220
transform 1 0 2596 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3420
timestamp 1710899220
transform 1 0 2612 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3421
timestamp 1710899220
transform 1 0 2556 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3422
timestamp 1710899220
transform 1 0 2236 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3423
timestamp 1710899220
transform 1 0 2132 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3424
timestamp 1710899220
transform 1 0 2300 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3425
timestamp 1710899220
transform 1 0 2188 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3426
timestamp 1710899220
transform 1 0 2332 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3427
timestamp 1710899220
transform 1 0 2252 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3428
timestamp 1710899220
transform 1 0 2036 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3429
timestamp 1710899220
transform 1 0 2020 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3430
timestamp 1710899220
transform 1 0 1988 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3431
timestamp 1710899220
transform 1 0 1980 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3432
timestamp 1710899220
transform 1 0 2124 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3433
timestamp 1710899220
transform 1 0 2060 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3434
timestamp 1710899220
transform 1 0 2036 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3435
timestamp 1710899220
transform 1 0 2260 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3436
timestamp 1710899220
transform 1 0 2220 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3437
timestamp 1710899220
transform 1 0 2116 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3438
timestamp 1710899220
transform 1 0 2260 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3439
timestamp 1710899220
transform 1 0 2156 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3440
timestamp 1710899220
transform 1 0 2124 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3441
timestamp 1710899220
transform 1 0 2172 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3442
timestamp 1710899220
transform 1 0 2116 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3443
timestamp 1710899220
transform 1 0 2028 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3444
timestamp 1710899220
transform 1 0 1492 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3445
timestamp 1710899220
transform 1 0 1380 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3446
timestamp 1710899220
transform 1 0 1380 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3447
timestamp 1710899220
transform 1 0 1684 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3448
timestamp 1710899220
transform 1 0 1524 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3449
timestamp 1710899220
transform 1 0 1508 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3450
timestamp 1710899220
transform 1 0 1764 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3451
timestamp 1710899220
transform 1 0 1620 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3452
timestamp 1710899220
transform 1 0 1156 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3453
timestamp 1710899220
transform 1 0 1324 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3454
timestamp 1710899220
transform 1 0 1324 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3455
timestamp 1710899220
transform 1 0 1012 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3456
timestamp 1710899220
transform 1 0 1284 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3457
timestamp 1710899220
transform 1 0 1140 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3458
timestamp 1710899220
transform 1 0 2468 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3459
timestamp 1710899220
transform 1 0 2412 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3460
timestamp 1710899220
transform 1 0 2332 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3461
timestamp 1710899220
transform 1 0 2220 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3462
timestamp 1710899220
transform 1 0 2668 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3463
timestamp 1710899220
transform 1 0 2572 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3464
timestamp 1710899220
transform 1 0 2324 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3465
timestamp 1710899220
transform 1 0 2148 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3466
timestamp 1710899220
transform 1 0 2044 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3467
timestamp 1710899220
transform 1 0 2124 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3468
timestamp 1710899220
transform 1 0 2004 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3469
timestamp 1710899220
transform 1 0 2100 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3470
timestamp 1710899220
transform 1 0 1996 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3471
timestamp 1710899220
transform 1 0 1572 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3472
timestamp 1710899220
transform 1 0 1996 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3473
timestamp 1710899220
transform 1 0 1892 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3474
timestamp 1710899220
transform 1 0 1652 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3475
timestamp 1710899220
transform 1 0 1588 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3476
timestamp 1710899220
transform 1 0 1556 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3477
timestamp 1710899220
transform 1 0 2036 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3478
timestamp 1710899220
transform 1 0 1996 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3479
timestamp 1710899220
transform 1 0 2124 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3480
timestamp 1710899220
transform 1 0 2020 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3481
timestamp 1710899220
transform 1 0 2132 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3482
timestamp 1710899220
transform 1 0 2028 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3483
timestamp 1710899220
transform 1 0 1756 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3484
timestamp 1710899220
transform 1 0 1700 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3485
timestamp 1710899220
transform 1 0 1644 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3486
timestamp 1710899220
transform 1 0 1620 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3487
timestamp 1710899220
transform 1 0 1612 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3488
timestamp 1710899220
transform 1 0 1556 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3489
timestamp 1710899220
transform 1 0 1804 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3490
timestamp 1710899220
transform 1 0 1700 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3491
timestamp 1710899220
transform 1 0 1588 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3492
timestamp 1710899220
transform 1 0 1236 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3493
timestamp 1710899220
transform 1 0 1188 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3494
timestamp 1710899220
transform 1 0 1044 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3495
timestamp 1710899220
transform 1 0 964 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3496
timestamp 1710899220
transform 1 0 1140 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3497
timestamp 1710899220
transform 1 0 1068 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3498
timestamp 1710899220
transform 1 0 892 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3499
timestamp 1710899220
transform 1 0 1044 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3500
timestamp 1710899220
transform 1 0 1012 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3501
timestamp 1710899220
transform 1 0 956 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3502
timestamp 1710899220
transform 1 0 924 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3503
timestamp 1710899220
transform 1 0 460 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3504
timestamp 1710899220
transform 1 0 340 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3505
timestamp 1710899220
transform 1 0 300 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3506
timestamp 1710899220
transform 1 0 532 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3507
timestamp 1710899220
transform 1 0 492 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3508
timestamp 1710899220
transform 1 0 492 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3509
timestamp 1710899220
transform 1 0 1004 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3510
timestamp 1710899220
transform 1 0 908 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3511
timestamp 1710899220
transform 1 0 844 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3512
timestamp 1710899220
transform 1 0 1012 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3513
timestamp 1710899220
transform 1 0 1012 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3514
timestamp 1710899220
transform 1 0 932 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3515
timestamp 1710899220
transform 1 0 1252 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3516
timestamp 1710899220
transform 1 0 1124 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3517
timestamp 1710899220
transform 1 0 1116 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3518
timestamp 1710899220
transform 1 0 964 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3519
timestamp 1710899220
transform 1 0 556 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3520
timestamp 1710899220
transform 1 0 316 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3521
timestamp 1710899220
transform 1 0 276 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3522
timestamp 1710899220
transform 1 0 388 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3523
timestamp 1710899220
transform 1 0 348 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3524
timestamp 1710899220
transform 1 0 300 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3525
timestamp 1710899220
transform 1 0 508 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3526
timestamp 1710899220
transform 1 0 428 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3527
timestamp 1710899220
transform 1 0 380 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3528
timestamp 1710899220
transform 1 0 332 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3529
timestamp 1710899220
transform 1 0 676 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3530
timestamp 1710899220
transform 1 0 676 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3531
timestamp 1710899220
transform 1 0 2052 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3532
timestamp 1710899220
transform 1 0 1948 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3533
timestamp 1710899220
transform 1 0 1924 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3534
timestamp 1710899220
transform 1 0 1820 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3535
timestamp 1710899220
transform 1 0 1796 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3536
timestamp 1710899220
transform 1 0 1644 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3537
timestamp 1710899220
transform 1 0 1620 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3538
timestamp 1710899220
transform 1 0 1564 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3539
timestamp 1710899220
transform 1 0 1596 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3540
timestamp 1710899220
transform 1 0 1524 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3541
timestamp 1710899220
transform 1 0 1452 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3542
timestamp 1710899220
transform 1 0 1396 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_3543
timestamp 1710899220
transform 1 0 1572 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_3544
timestamp 1710899220
transform 1 0 1548 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3545
timestamp 1710899220
transform 1 0 1516 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3546
timestamp 1710899220
transform 1 0 1372 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_3547
timestamp 1710899220
transform 1 0 1932 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3548
timestamp 1710899220
transform 1 0 1852 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3549
timestamp 1710899220
transform 1 0 1836 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3550
timestamp 1710899220
transform 1 0 1940 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3551
timestamp 1710899220
transform 1 0 1940 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3552
timestamp 1710899220
transform 1 0 1884 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3553
timestamp 1710899220
transform 1 0 1852 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3554
timestamp 1710899220
transform 1 0 1788 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3555
timestamp 1710899220
transform 1 0 1444 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3556
timestamp 1710899220
transform 1 0 1396 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3557
timestamp 1710899220
transform 1 0 1068 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_3558
timestamp 1710899220
transform 1 0 1604 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3559
timestamp 1710899220
transform 1 0 1596 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_3560
timestamp 1710899220
transform 1 0 1508 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3561
timestamp 1710899220
transform 1 0 1556 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3562
timestamp 1710899220
transform 1 0 1556 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3563
timestamp 1710899220
transform 1 0 1348 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3564
timestamp 1710899220
transform 1 0 1204 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_3565
timestamp 1710899220
transform 1 0 1028 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3566
timestamp 1710899220
transform 1 0 1028 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_3567
timestamp 1710899220
transform 1 0 1156 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3568
timestamp 1710899220
transform 1 0 1132 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3569
timestamp 1710899220
transform 1 0 1060 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3570
timestamp 1710899220
transform 1 0 1052 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_3571
timestamp 1710899220
transform 1 0 948 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3572
timestamp 1710899220
transform 1 0 940 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_3573
timestamp 1710899220
transform 1 0 924 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3574
timestamp 1710899220
transform 1 0 852 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3575
timestamp 1710899220
transform 1 0 780 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3576
timestamp 1710899220
transform 1 0 708 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3577
timestamp 1710899220
transform 1 0 748 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3578
timestamp 1710899220
transform 1 0 740 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3579
timestamp 1710899220
transform 1 0 684 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3580
timestamp 1710899220
transform 1 0 644 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3581
timestamp 1710899220
transform 1 0 596 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3582
timestamp 1710899220
transform 1 0 860 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3583
timestamp 1710899220
transform 1 0 836 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3584
timestamp 1710899220
transform 1 0 948 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3585
timestamp 1710899220
transform 1 0 900 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3586
timestamp 1710899220
transform 1 0 1388 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3587
timestamp 1710899220
transform 1 0 1244 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3588
timestamp 1710899220
transform 1 0 1140 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3589
timestamp 1710899220
transform 1 0 1100 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_3590
timestamp 1710899220
transform 1 0 532 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3591
timestamp 1710899220
transform 1 0 468 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3592
timestamp 1710899220
transform 1 0 436 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3593
timestamp 1710899220
transform 1 0 492 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3594
timestamp 1710899220
transform 1 0 476 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3595
timestamp 1710899220
transform 1 0 412 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3596
timestamp 1710899220
transform 1 0 636 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3597
timestamp 1710899220
transform 1 0 588 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3598
timestamp 1710899220
transform 1 0 540 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3599
timestamp 1710899220
transform 1 0 492 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_3600
timestamp 1710899220
transform 1 0 1084 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3601
timestamp 1710899220
transform 1 0 716 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3602
timestamp 1710899220
transform 1 0 660 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3603
timestamp 1710899220
transform 1 0 644 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_3604
timestamp 1710899220
transform 1 0 580 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3605
timestamp 1710899220
transform 1 0 1972 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3606
timestamp 1710899220
transform 1 0 1836 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3607
timestamp 1710899220
transform 1 0 1924 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3608
timestamp 1710899220
transform 1 0 1812 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3609
timestamp 1710899220
transform 1 0 2300 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3610
timestamp 1710899220
transform 1 0 2252 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3611
timestamp 1710899220
transform 1 0 2244 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3612
timestamp 1710899220
transform 1 0 2428 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3613
timestamp 1710899220
transform 1 0 2308 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3614
timestamp 1710899220
transform 1 0 2276 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3615
timestamp 1710899220
transform 1 0 2172 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3616
timestamp 1710899220
transform 1 0 2116 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3617
timestamp 1710899220
transform 1 0 2332 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3618
timestamp 1710899220
transform 1 0 2204 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3619
timestamp 1710899220
transform 1 0 2172 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3620
timestamp 1710899220
transform 1 0 2140 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3621
timestamp 1710899220
transform 1 0 2076 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_3622
timestamp 1710899220
transform 1 0 2076 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3623
timestamp 1710899220
transform 1 0 1964 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3624
timestamp 1710899220
transform 1 0 1908 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3625
timestamp 1710899220
transform 1 0 1924 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3626
timestamp 1710899220
transform 1 0 1852 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3627
timestamp 1710899220
transform 1 0 1964 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3628
timestamp 1710899220
transform 1 0 1908 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3629
timestamp 1710899220
transform 1 0 1964 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3630
timestamp 1710899220
transform 1 0 1908 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3631
timestamp 1710899220
transform 1 0 1988 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3632
timestamp 1710899220
transform 1 0 1924 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3633
timestamp 1710899220
transform 1 0 2292 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3634
timestamp 1710899220
transform 1 0 2180 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3635
timestamp 1710899220
transform 1 0 2068 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3636
timestamp 1710899220
transform 1 0 2148 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3637
timestamp 1710899220
transform 1 0 2060 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3638
timestamp 1710899220
transform 1 0 2044 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3639
timestamp 1710899220
transform 1 0 2412 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3640
timestamp 1710899220
transform 1 0 2284 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3641
timestamp 1710899220
transform 1 0 2156 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3642
timestamp 1710899220
transform 1 0 2388 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3643
timestamp 1710899220
transform 1 0 2316 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3644
timestamp 1710899220
transform 1 0 2204 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3645
timestamp 1710899220
transform 1 0 2516 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3646
timestamp 1710899220
transform 1 0 2404 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3647
timestamp 1710899220
transform 1 0 2644 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3648
timestamp 1710899220
transform 1 0 2596 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3649
timestamp 1710899220
transform 1 0 2484 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3650
timestamp 1710899220
transform 1 0 2668 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3651
timestamp 1710899220
transform 1 0 2556 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3652
timestamp 1710899220
transform 1 0 2444 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3653
timestamp 1710899220
transform 1 0 2500 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3654
timestamp 1710899220
transform 1 0 2364 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3655
timestamp 1710899220
transform 1 0 2652 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3656
timestamp 1710899220
transform 1 0 2556 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3657
timestamp 1710899220
transform 1 0 2444 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3658
timestamp 1710899220
transform 1 0 2668 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3659
timestamp 1710899220
transform 1 0 2556 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3660
timestamp 1710899220
transform 1 0 2444 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3661
timestamp 1710899220
transform 1 0 2652 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3662
timestamp 1710899220
transform 1 0 2540 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3663
timestamp 1710899220
transform 1 0 2428 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3664
timestamp 1710899220
transform 1 0 2668 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3665
timestamp 1710899220
transform 1 0 2572 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3666
timestamp 1710899220
transform 1 0 2460 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3667
timestamp 1710899220
transform 1 0 2372 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3668
timestamp 1710899220
transform 1 0 2316 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3669
timestamp 1710899220
transform 1 0 2372 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3670
timestamp 1710899220
transform 1 0 2316 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3671
timestamp 1710899220
transform 1 0 2668 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3672
timestamp 1710899220
transform 1 0 2572 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3673
timestamp 1710899220
transform 1 0 2460 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3674
timestamp 1710899220
transform 1 0 2660 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3675
timestamp 1710899220
transform 1 0 2620 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3676
timestamp 1710899220
transform 1 0 2548 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3677
timestamp 1710899220
transform 1 0 2540 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3678
timestamp 1710899220
transform 1 0 2500 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3679
timestamp 1710899220
transform 1 0 2428 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3680
timestamp 1710899220
transform 1 0 2364 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3681
timestamp 1710899220
transform 1 0 2348 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3682
timestamp 1710899220
transform 1 0 2324 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3683
timestamp 1710899220
transform 1 0 2372 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3684
timestamp 1710899220
transform 1 0 2372 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3685
timestamp 1710899220
transform 1 0 2556 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3686
timestamp 1710899220
transform 1 0 2492 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3687
timestamp 1710899220
transform 1 0 2380 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3688
timestamp 1710899220
transform 1 0 2668 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3689
timestamp 1710899220
transform 1 0 2540 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3690
timestamp 1710899220
transform 1 0 2500 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3691
timestamp 1710899220
transform 1 0 2652 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3692
timestamp 1710899220
transform 1 0 2652 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3693
timestamp 1710899220
transform 1 0 2612 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3694
timestamp 1710899220
transform 1 0 2052 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3695
timestamp 1710899220
transform 1 0 1996 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3696
timestamp 1710899220
transform 1 0 2284 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3697
timestamp 1710899220
transform 1 0 2284 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_3698
timestamp 1710899220
transform 1 0 2148 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3699
timestamp 1710899220
transform 1 0 2020 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3700
timestamp 1710899220
transform 1 0 2244 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3701
timestamp 1710899220
transform 1 0 2244 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_3702
timestamp 1710899220
transform 1 0 2244 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3703
timestamp 1710899220
transform 1 0 2196 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3704
timestamp 1710899220
transform 1 0 2196 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3705
timestamp 1710899220
transform 1 0 2172 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3706
timestamp 1710899220
transform 1 0 2164 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3707
timestamp 1710899220
transform 1 0 2148 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_3708
timestamp 1710899220
transform 1 0 2220 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3709
timestamp 1710899220
transform 1 0 2180 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3710
timestamp 1710899220
transform 1 0 2108 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3711
timestamp 1710899220
transform 1 0 1196 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3712
timestamp 1710899220
transform 1 0 1100 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3713
timestamp 1710899220
transform 1 0 1092 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3714
timestamp 1710899220
transform 1 0 1076 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3715
timestamp 1710899220
transform 1 0 1052 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3716
timestamp 1710899220
transform 1 0 940 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3717
timestamp 1710899220
transform 1 0 820 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3718
timestamp 1710899220
transform 1 0 820 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3719
timestamp 1710899220
transform 1 0 812 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_3720
timestamp 1710899220
transform 1 0 780 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3721
timestamp 1710899220
transform 1 0 764 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3722
timestamp 1710899220
transform 1 0 740 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_3723
timestamp 1710899220
transform 1 0 660 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3724
timestamp 1710899220
transform 1 0 620 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3725
timestamp 1710899220
transform 1 0 620 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3726
timestamp 1710899220
transform 1 0 604 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3727
timestamp 1710899220
transform 1 0 580 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3728
timestamp 1710899220
transform 1 0 580 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3729
timestamp 1710899220
transform 1 0 572 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3730
timestamp 1710899220
transform 1 0 564 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3731
timestamp 1710899220
transform 1 0 524 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3732
timestamp 1710899220
transform 1 0 516 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3733
timestamp 1710899220
transform 1 0 468 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3734
timestamp 1710899220
transform 1 0 356 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3735
timestamp 1710899220
transform 1 0 348 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3736
timestamp 1710899220
transform 1 0 324 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3737
timestamp 1710899220
transform 1 0 1188 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3738
timestamp 1710899220
transform 1 0 1132 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3739
timestamp 1710899220
transform 1 0 1092 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3740
timestamp 1710899220
transform 1 0 1084 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3741
timestamp 1710899220
transform 1 0 1060 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3742
timestamp 1710899220
transform 1 0 844 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3743
timestamp 1710899220
transform 1 0 828 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3744
timestamp 1710899220
transform 1 0 756 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3745
timestamp 1710899220
transform 1 0 668 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3746
timestamp 1710899220
transform 1 0 620 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3747
timestamp 1710899220
transform 1 0 596 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3748
timestamp 1710899220
transform 1 0 572 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3749
timestamp 1710899220
transform 1 0 556 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3750
timestamp 1710899220
transform 1 0 548 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_3751
timestamp 1710899220
transform 1 0 484 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3752
timestamp 1710899220
transform 1 0 396 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3753
timestamp 1710899220
transform 1 0 308 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_3754
timestamp 1710899220
transform 1 0 132 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3755
timestamp 1710899220
transform 1 0 100 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3756
timestamp 1710899220
transform 1 0 1308 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3757
timestamp 1710899220
transform 1 0 1252 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_3758
timestamp 1710899220
transform 1 0 1236 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_3759
timestamp 1710899220
transform 1 0 1140 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3760
timestamp 1710899220
transform 1 0 1092 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3761
timestamp 1710899220
transform 1 0 1036 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3762
timestamp 1710899220
transform 1 0 1028 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3763
timestamp 1710899220
transform 1 0 908 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3764
timestamp 1710899220
transform 1 0 900 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3765
timestamp 1710899220
transform 1 0 860 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3766
timestamp 1710899220
transform 1 0 396 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3767
timestamp 1710899220
transform 1 0 364 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3768
timestamp 1710899220
transform 1 0 324 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3769
timestamp 1710899220
transform 1 0 300 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3770
timestamp 1710899220
transform 1 0 228 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3771
timestamp 1710899220
transform 1 0 188 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3772
timestamp 1710899220
transform 1 0 140 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3773
timestamp 1710899220
transform 1 0 116 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3774
timestamp 1710899220
transform 1 0 108 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3775
timestamp 1710899220
transform 1 0 1444 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3776
timestamp 1710899220
transform 1 0 1308 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_3777
timestamp 1710899220
transform 1 0 1220 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3778
timestamp 1710899220
transform 1 0 1116 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3779
timestamp 1710899220
transform 1 0 1100 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3780
timestamp 1710899220
transform 1 0 1076 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3781
timestamp 1710899220
transform 1 0 716 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_3782
timestamp 1710899220
transform 1 0 668 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3783
timestamp 1710899220
transform 1 0 660 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3784
timestamp 1710899220
transform 1 0 212 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3785
timestamp 1710899220
transform 1 0 188 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3786
timestamp 1710899220
transform 1 0 132 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_3787
timestamp 1710899220
transform 1 0 132 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_3788
timestamp 1710899220
transform 1 0 124 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3789
timestamp 1710899220
transform 1 0 84 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_3790
timestamp 1710899220
transform 1 0 1292 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3791
timestamp 1710899220
transform 1 0 1188 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3792
timestamp 1710899220
transform 1 0 1172 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3793
timestamp 1710899220
transform 1 0 1076 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3794
timestamp 1710899220
transform 1 0 1044 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_3795
timestamp 1710899220
transform 1 0 1012 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_3796
timestamp 1710899220
transform 1 0 756 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3797
timestamp 1710899220
transform 1 0 716 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3798
timestamp 1710899220
transform 1 0 76 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3799
timestamp 1710899220
transform 1 0 76 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3800
timestamp 1710899220
transform 1 0 76 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3801
timestamp 1710899220
transform 1 0 2180 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3802
timestamp 1710899220
transform 1 0 2132 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3803
timestamp 1710899220
transform 1 0 2116 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_3804
timestamp 1710899220
transform 1 0 1884 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3805
timestamp 1710899220
transform 1 0 1828 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3806
timestamp 1710899220
transform 1 0 1732 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3807
timestamp 1710899220
transform 1 0 556 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3808
timestamp 1710899220
transform 1 0 548 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3809
timestamp 1710899220
transform 1 0 532 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_3810
timestamp 1710899220
transform 1 0 500 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3811
timestamp 1710899220
transform 1 0 500 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3812
timestamp 1710899220
transform 1 0 484 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3813
timestamp 1710899220
transform 1 0 1852 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3814
timestamp 1710899220
transform 1 0 1788 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3815
timestamp 1710899220
transform 1 0 1700 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3816
timestamp 1710899220
transform 1 0 924 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3817
timestamp 1710899220
transform 1 0 492 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_3818
timestamp 1710899220
transform 1 0 468 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3819
timestamp 1710899220
transform 1 0 452 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3820
timestamp 1710899220
transform 1 0 452 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3821
timestamp 1710899220
transform 1 0 1964 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3822
timestamp 1710899220
transform 1 0 1908 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3823
timestamp 1710899220
transform 1 0 1812 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_3824
timestamp 1710899220
transform 1 0 1788 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3825
timestamp 1710899220
transform 1 0 1580 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3826
timestamp 1710899220
transform 1 0 892 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3827
timestamp 1710899220
transform 1 0 668 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3828
timestamp 1710899220
transform 1 0 428 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3829
timestamp 1710899220
transform 1 0 420 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3830
timestamp 1710899220
transform 1 0 396 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3831
timestamp 1710899220
transform 1 0 1668 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3832
timestamp 1710899220
transform 1 0 1668 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3833
timestamp 1710899220
transform 1 0 1628 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3834
timestamp 1710899220
transform 1 0 1572 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3835
timestamp 1710899220
transform 1 0 1052 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3836
timestamp 1710899220
transform 1 0 636 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3837
timestamp 1710899220
transform 1 0 388 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_3838
timestamp 1710899220
transform 1 0 388 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3839
timestamp 1710899220
transform 1 0 348 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3840
timestamp 1710899220
transform 1 0 1724 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3841
timestamp 1710899220
transform 1 0 1684 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3842
timestamp 1710899220
transform 1 0 1588 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3843
timestamp 1710899220
transform 1 0 1564 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3844
timestamp 1710899220
transform 1 0 1540 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3845
timestamp 1710899220
transform 1 0 1012 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3846
timestamp 1710899220
transform 1 0 668 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3847
timestamp 1710899220
transform 1 0 652 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3848
timestamp 1710899220
transform 1 0 572 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3849
timestamp 1710899220
transform 1 0 484 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3850
timestamp 1710899220
transform 1 0 1532 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3851
timestamp 1710899220
transform 1 0 1524 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3852
timestamp 1710899220
transform 1 0 1492 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3853
timestamp 1710899220
transform 1 0 700 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3854
timestamp 1710899220
transform 1 0 636 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3855
timestamp 1710899220
transform 1 0 620 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3856
timestamp 1710899220
transform 1 0 540 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3857
timestamp 1710899220
transform 1 0 444 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3858
timestamp 1710899220
transform 1 0 1892 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3859
timestamp 1710899220
transform 1 0 1860 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3860
timestamp 1710899220
transform 1 0 1844 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3861
timestamp 1710899220
transform 1 0 1700 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3862
timestamp 1710899220
transform 1 0 716 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3863
timestamp 1710899220
transform 1 0 700 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3864
timestamp 1710899220
transform 1 0 660 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3865
timestamp 1710899220
transform 1 0 652 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_3866
timestamp 1710899220
transform 1 0 636 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3867
timestamp 1710899220
transform 1 0 396 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3868
timestamp 1710899220
transform 1 0 1932 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3869
timestamp 1710899220
transform 1 0 1924 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3870
timestamp 1710899220
transform 1 0 1924 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3871
timestamp 1710899220
transform 1 0 1884 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3872
timestamp 1710899220
transform 1 0 1876 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3873
timestamp 1710899220
transform 1 0 684 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3874
timestamp 1710899220
transform 1 0 684 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3875
timestamp 1710899220
transform 1 0 628 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3876
timestamp 1710899220
transform 1 0 604 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3877
timestamp 1710899220
transform 1 0 364 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3878
timestamp 1710899220
transform 1 0 1604 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3879
timestamp 1710899220
transform 1 0 1524 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3880
timestamp 1710899220
transform 1 0 1404 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3881
timestamp 1710899220
transform 1 0 692 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3882
timestamp 1710899220
transform 1 0 604 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3883
timestamp 1710899220
transform 1 0 460 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3884
timestamp 1710899220
transform 1 0 444 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3885
timestamp 1710899220
transform 1 0 436 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3886
timestamp 1710899220
transform 1 0 876 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3887
timestamp 1710899220
transform 1 0 876 0 1 1455
box -2 -2 2 2
use M2_M1  M2_M1_3888
timestamp 1710899220
transform 1 0 860 0 1 1455
box -2 -2 2 2
use M2_M1  M2_M1_3889
timestamp 1710899220
transform 1 0 852 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3890
timestamp 1710899220
transform 1 0 844 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3891
timestamp 1710899220
transform 1 0 836 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3892
timestamp 1710899220
transform 1 0 556 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3893
timestamp 1710899220
transform 1 0 428 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3894
timestamp 1710899220
transform 1 0 404 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3895
timestamp 1710899220
transform 1 0 404 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3896
timestamp 1710899220
transform 1 0 404 0 1 1185
box -2 -2 2 2
use M2_M1  M2_M1_3897
timestamp 1710899220
transform 1 0 1564 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3898
timestamp 1710899220
transform 1 0 1556 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3899
timestamp 1710899220
transform 1 0 1516 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3900
timestamp 1710899220
transform 1 0 1476 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3901
timestamp 1710899220
transform 1 0 1364 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3902
timestamp 1710899220
transform 1 0 900 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3903
timestamp 1710899220
transform 1 0 868 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3904
timestamp 1710899220
transform 1 0 692 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3905
timestamp 1710899220
transform 1 0 380 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3906
timestamp 1710899220
transform 1 0 380 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3907
timestamp 1710899220
transform 1 0 372 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3908
timestamp 1710899220
transform 1 0 1580 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3909
timestamp 1710899220
transform 1 0 1532 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3910
timestamp 1710899220
transform 1 0 1356 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3911
timestamp 1710899220
transform 1 0 1308 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3912
timestamp 1710899220
transform 1 0 1188 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3913
timestamp 1710899220
transform 1 0 1028 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3914
timestamp 1710899220
transform 1 0 660 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3915
timestamp 1710899220
transform 1 0 348 0 1 1055
box -2 -2 2 2
use M2_M1  M2_M1_3916
timestamp 1710899220
transform 1 0 348 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3917
timestamp 1710899220
transform 1 0 340 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3918
timestamp 1710899220
transform 1 0 332 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3919
timestamp 1710899220
transform 1 0 332 0 1 1055
box -2 -2 2 2
use M2_M1  M2_M1_3920
timestamp 1710899220
transform 1 0 1100 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3921
timestamp 1710899220
transform 1 0 1060 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3922
timestamp 1710899220
transform 1 0 1020 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3923
timestamp 1710899220
transform 1 0 988 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3924
timestamp 1710899220
transform 1 0 956 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3925
timestamp 1710899220
transform 1 0 564 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3926
timestamp 1710899220
transform 1 0 564 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3927
timestamp 1710899220
transform 1 0 548 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3928
timestamp 1710899220
transform 1 0 484 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3929
timestamp 1710899220
transform 1 0 1228 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3930
timestamp 1710899220
transform 1 0 1052 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3931
timestamp 1710899220
transform 1 0 972 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3932
timestamp 1710899220
transform 1 0 892 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3933
timestamp 1710899220
transform 1 0 868 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3934
timestamp 1710899220
transform 1 0 724 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3935
timestamp 1710899220
transform 1 0 532 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3936
timestamp 1710899220
transform 1 0 532 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3937
timestamp 1710899220
transform 1 0 492 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3938
timestamp 1710899220
transform 1 0 452 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3939
timestamp 1710899220
transform 1 0 1076 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3940
timestamp 1710899220
transform 1 0 916 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3941
timestamp 1710899220
transform 1 0 908 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3942
timestamp 1710899220
transform 1 0 716 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3943
timestamp 1710899220
transform 1 0 620 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3944
timestamp 1710899220
transform 1 0 604 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3945
timestamp 1710899220
transform 1 0 580 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3946
timestamp 1710899220
transform 1 0 428 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3947
timestamp 1710899220
transform 1 0 1116 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3948
timestamp 1710899220
transform 1 0 716 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3949
timestamp 1710899220
transform 1 0 700 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3950
timestamp 1710899220
transform 1 0 588 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3951
timestamp 1710899220
transform 1 0 572 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3952
timestamp 1710899220
transform 1 0 548 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3953
timestamp 1710899220
transform 1 0 452 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3954
timestamp 1710899220
transform 1 0 396 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3955
timestamp 1710899220
transform 1 0 796 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3956
timestamp 1710899220
transform 1 0 732 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3957
timestamp 1710899220
transform 1 0 708 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3958
timestamp 1710899220
transform 1 0 668 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3959
timestamp 1710899220
transform 1 0 460 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3960
timestamp 1710899220
transform 1 0 444 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3961
timestamp 1710899220
transform 1 0 436 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3962
timestamp 1710899220
transform 1 0 436 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3963
timestamp 1710899220
transform 1 0 396 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3964
timestamp 1710899220
transform 1 0 900 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3965
timestamp 1710899220
transform 1 0 892 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3966
timestamp 1710899220
transform 1 0 860 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3967
timestamp 1710899220
transform 1 0 636 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3968
timestamp 1710899220
transform 1 0 532 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3969
timestamp 1710899220
transform 1 0 484 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3970
timestamp 1710899220
transform 1 0 412 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3971
timestamp 1710899220
transform 1 0 404 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3972
timestamp 1710899220
transform 1 0 404 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3973
timestamp 1710899220
transform 1 0 1004 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3974
timestamp 1710899220
transform 1 0 996 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3975
timestamp 1710899220
transform 1 0 972 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3976
timestamp 1710899220
transform 1 0 924 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3977
timestamp 1710899220
transform 1 0 916 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3978
timestamp 1710899220
transform 1 0 868 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3979
timestamp 1710899220
transform 1 0 812 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3980
timestamp 1710899220
transform 1 0 708 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3981
timestamp 1710899220
transform 1 0 388 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3982
timestamp 1710899220
transform 1 0 356 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3983
timestamp 1710899220
transform 1 0 348 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3984
timestamp 1710899220
transform 1 0 1012 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3985
timestamp 1710899220
transform 1 0 964 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3986
timestamp 1710899220
transform 1 0 940 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3987
timestamp 1710899220
transform 1 0 924 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3988
timestamp 1710899220
transform 1 0 892 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3989
timestamp 1710899220
transform 1 0 828 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3990
timestamp 1710899220
transform 1 0 676 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3991
timestamp 1710899220
transform 1 0 340 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3992
timestamp 1710899220
transform 1 0 324 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3993
timestamp 1710899220
transform 1 0 316 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3994
timestamp 1710899220
transform 1 0 1068 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3995
timestamp 1710899220
transform 1 0 1036 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3996
timestamp 1710899220
transform 1 0 972 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3997
timestamp 1710899220
transform 1 0 972 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3998
timestamp 1710899220
transform 1 0 956 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3999
timestamp 1710899220
transform 1 0 540 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4000
timestamp 1710899220
transform 1 0 540 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4001
timestamp 1710899220
transform 1 0 516 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4002
timestamp 1710899220
transform 1 0 484 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4003
timestamp 1710899220
transform 1 0 476 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4004
timestamp 1710899220
transform 1 0 556 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4005
timestamp 1710899220
transform 1 0 548 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4006
timestamp 1710899220
transform 1 0 508 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4007
timestamp 1710899220
transform 1 0 484 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4008
timestamp 1710899220
transform 1 0 452 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4009
timestamp 1710899220
transform 1 0 444 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4010
timestamp 1710899220
transform 1 0 444 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4011
timestamp 1710899220
transform 1 0 444 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4012
timestamp 1710899220
transform 1 0 444 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4013
timestamp 1710899220
transform 1 0 908 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4014
timestamp 1710899220
transform 1 0 900 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4015
timestamp 1710899220
transform 1 0 676 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4016
timestamp 1710899220
transform 1 0 588 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4017
timestamp 1710899220
transform 1 0 492 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4018
timestamp 1710899220
transform 1 0 460 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4019
timestamp 1710899220
transform 1 0 404 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4020
timestamp 1710899220
transform 1 0 396 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4021
timestamp 1710899220
transform 1 0 388 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4022
timestamp 1710899220
transform 1 0 364 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4023
timestamp 1710899220
transform 1 0 620 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4024
timestamp 1710899220
transform 1 0 556 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4025
timestamp 1710899220
transform 1 0 556 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4026
timestamp 1710899220
transform 1 0 548 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4027
timestamp 1710899220
transform 1 0 452 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4028
timestamp 1710899220
transform 1 0 420 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4029
timestamp 1710899220
transform 1 0 364 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4030
timestamp 1710899220
transform 1 0 356 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4031
timestamp 1710899220
transform 1 0 932 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4032
timestamp 1710899220
transform 1 0 764 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4033
timestamp 1710899220
transform 1 0 572 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4034
timestamp 1710899220
transform 1 0 2428 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_4035
timestamp 1710899220
transform 1 0 2420 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4036
timestamp 1710899220
transform 1 0 2268 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_4037
timestamp 1710899220
transform 1 0 2284 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4038
timestamp 1710899220
transform 1 0 2268 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_4039
timestamp 1710899220
transform 1 0 2252 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4040
timestamp 1710899220
transform 1 0 2244 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_4041
timestamp 1710899220
transform 1 0 2244 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_4042
timestamp 1710899220
transform 1 0 2164 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4043
timestamp 1710899220
transform 1 0 2100 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4044
timestamp 1710899220
transform 1 0 2460 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4045
timestamp 1710899220
transform 1 0 2452 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4046
timestamp 1710899220
transform 1 0 2420 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4047
timestamp 1710899220
transform 1 0 2620 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4048
timestamp 1710899220
transform 1 0 2604 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4049
timestamp 1710899220
transform 1 0 2604 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4050
timestamp 1710899220
transform 1 0 2580 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4051
timestamp 1710899220
transform 1 0 2572 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4052
timestamp 1710899220
transform 1 0 2556 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4053
timestamp 1710899220
transform 1 0 2668 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4054
timestamp 1710899220
transform 1 0 2660 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4055
timestamp 1710899220
transform 1 0 2628 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4056
timestamp 1710899220
transform 1 0 2620 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4057
timestamp 1710899220
transform 1 0 2668 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4058
timestamp 1710899220
transform 1 0 2644 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_4059
timestamp 1710899220
transform 1 0 2620 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4060
timestamp 1710899220
transform 1 0 2612 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4061
timestamp 1710899220
transform 1 0 2596 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4062
timestamp 1710899220
transform 1 0 2596 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4063
timestamp 1710899220
transform 1 0 2564 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4064
timestamp 1710899220
transform 1 0 2636 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4065
timestamp 1710899220
transform 1 0 2588 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_4066
timestamp 1710899220
transform 1 0 2564 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_4067
timestamp 1710899220
transform 1 0 2500 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4068
timestamp 1710899220
transform 1 0 2492 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4069
timestamp 1710899220
transform 1 0 2468 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4070
timestamp 1710899220
transform 1 0 1324 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4071
timestamp 1710899220
transform 1 0 1292 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4072
timestamp 1710899220
transform 1 0 1964 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4073
timestamp 1710899220
transform 1 0 1916 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4074
timestamp 1710899220
transform 1 0 1852 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4075
timestamp 1710899220
transform 1 0 1828 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4076
timestamp 1710899220
transform 1 0 1804 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_0
timestamp 1710899220
transform 1 0 2300 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1
timestamp 1710899220
transform 1 0 2188 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2
timestamp 1710899220
transform 1 0 2196 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_3
timestamp 1710899220
transform 1 0 2092 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4
timestamp 1710899220
transform 1 0 2108 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_5
timestamp 1710899220
transform 1 0 1980 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_6
timestamp 1710899220
transform 1 0 1996 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_7
timestamp 1710899220
transform 1 0 1948 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_8
timestamp 1710899220
transform 1 0 2412 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_9
timestamp 1710899220
transform 1 0 2236 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_10
timestamp 1710899220
transform 1 0 2468 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_11
timestamp 1710899220
transform 1 0 2428 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_12
timestamp 1710899220
transform 1 0 2468 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_13
timestamp 1710899220
transform 1 0 2372 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_14
timestamp 1710899220
transform 1 0 2444 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_15
timestamp 1710899220
transform 1 0 2396 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_16
timestamp 1710899220
transform 1 0 2484 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_17
timestamp 1710899220
transform 1 0 2388 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_18
timestamp 1710899220
transform 1 0 2452 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_19
timestamp 1710899220
transform 1 0 2412 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_20
timestamp 1710899220
transform 1 0 2572 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_21
timestamp 1710899220
transform 1 0 2436 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_22
timestamp 1710899220
transform 1 0 2444 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_23
timestamp 1710899220
transform 1 0 2356 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_24
timestamp 1710899220
transform 1 0 2500 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_25
timestamp 1710899220
transform 1 0 2412 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_26
timestamp 1710899220
transform 1 0 2620 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_27
timestamp 1710899220
transform 1 0 2532 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_28
timestamp 1710899220
transform 1 0 1348 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_29
timestamp 1710899220
transform 1 0 1164 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_30
timestamp 1710899220
transform 1 0 1260 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_31
timestamp 1710899220
transform 1 0 1012 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_32
timestamp 1710899220
transform 1 0 1100 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_33
timestamp 1710899220
transform 1 0 804 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_34
timestamp 1710899220
transform 1 0 900 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_35
timestamp 1710899220
transform 1 0 500 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_36
timestamp 1710899220
transform 1 0 2132 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_37
timestamp 1710899220
transform 1 0 2116 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_38
timestamp 1710899220
transform 1 0 2156 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_39
timestamp 1710899220
transform 1 0 2060 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_40
timestamp 1710899220
transform 1 0 1732 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_41
timestamp 1710899220
transform 1 0 1652 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_42
timestamp 1710899220
transform 1 0 1652 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_43
timestamp 1710899220
transform 1 0 1604 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_44
timestamp 1710899220
transform 1 0 1604 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_45
timestamp 1710899220
transform 1 0 1524 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_46
timestamp 1710899220
transform 1 0 1388 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_47
timestamp 1710899220
transform 1 0 1756 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_48
timestamp 1710899220
transform 1 0 1684 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_49
timestamp 1710899220
transform 1 0 1668 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_50
timestamp 1710899220
transform 1 0 1596 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_51
timestamp 1710899220
transform 1 0 1548 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_52
timestamp 1710899220
transform 1 0 1468 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_53
timestamp 1710899220
transform 1 0 1564 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_54
timestamp 1710899220
transform 1 0 1492 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_55
timestamp 1710899220
transform 1 0 1444 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_56
timestamp 1710899220
transform 1 0 1436 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_57
timestamp 1710899220
transform 1 0 1380 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_58
timestamp 1710899220
transform 1 0 1356 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_59
timestamp 1710899220
transform 1 0 1340 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_60
timestamp 1710899220
transform 1 0 1244 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_61
timestamp 1710899220
transform 1 0 1164 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_62
timestamp 1710899220
transform 1 0 1092 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_63
timestamp 1710899220
transform 1 0 956 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_64
timestamp 1710899220
transform 1 0 900 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_65
timestamp 1710899220
transform 1 0 948 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_66
timestamp 1710899220
transform 1 0 892 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_67
timestamp 1710899220
transform 1 0 788 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_68
timestamp 1710899220
transform 1 0 764 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_69
timestamp 1710899220
transform 1 0 636 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_70
timestamp 1710899220
transform 1 0 564 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_71
timestamp 1710899220
transform 1 0 652 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_72
timestamp 1710899220
transform 1 0 572 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_73
timestamp 1710899220
transform 1 0 572 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_74
timestamp 1710899220
transform 1 0 460 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_75
timestamp 1710899220
transform 1 0 332 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_76
timestamp 1710899220
transform 1 0 268 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_77
timestamp 1710899220
transform 1 0 380 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_78
timestamp 1710899220
transform 1 0 300 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_79
timestamp 1710899220
transform 1 0 236 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_80
timestamp 1710899220
transform 1 0 204 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_81
timestamp 1710899220
transform 1 0 2516 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_82
timestamp 1710899220
transform 1 0 2492 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_83
timestamp 1710899220
transform 1 0 2484 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_84
timestamp 1710899220
transform 1 0 2460 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_85
timestamp 1710899220
transform 1 0 2380 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_86
timestamp 1710899220
transform 1 0 2356 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_87
timestamp 1710899220
transform 1 0 2276 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_88
timestamp 1710899220
transform 1 0 2612 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_89
timestamp 1710899220
transform 1 0 2540 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_90
timestamp 1710899220
transform 1 0 2444 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_91
timestamp 1710899220
transform 1 0 2636 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_92
timestamp 1710899220
transform 1 0 2612 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_93
timestamp 1710899220
transform 1 0 2476 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_94
timestamp 1710899220
transform 1 0 2460 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_95
timestamp 1710899220
transform 1 0 1724 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_96
timestamp 1710899220
transform 1 0 1596 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_97
timestamp 1710899220
transform 1 0 1540 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_98
timestamp 1710899220
transform 1 0 1452 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_99
timestamp 1710899220
transform 1 0 1220 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_100
timestamp 1710899220
transform 1 0 1148 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_101
timestamp 1710899220
transform 1 0 1068 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_102
timestamp 1710899220
transform 1 0 852 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_103
timestamp 1710899220
transform 1 0 756 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_104
timestamp 1710899220
transform 1 0 684 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_105
timestamp 1710899220
transform 1 0 484 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_106
timestamp 1710899220
transform 1 0 404 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_107
timestamp 1710899220
transform 1 0 276 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_108
timestamp 1710899220
transform 1 0 196 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_109
timestamp 1710899220
transform 1 0 124 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_110
timestamp 1710899220
transform 1 0 148 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_111
timestamp 1710899220
transform 1 0 76 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_112
timestamp 1710899220
transform 1 0 516 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_113
timestamp 1710899220
transform 1 0 420 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_114
timestamp 1710899220
transform 1 0 492 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_115
timestamp 1710899220
transform 1 0 388 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_116
timestamp 1710899220
transform 1 0 644 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_117
timestamp 1710899220
transform 1 0 588 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_118
timestamp 1710899220
transform 1 0 772 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_119
timestamp 1710899220
transform 1 0 700 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_120
timestamp 1710899220
transform 1 0 628 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_121
timestamp 1710899220
transform 1 0 828 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_122
timestamp 1710899220
transform 1 0 692 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_123
timestamp 1710899220
transform 1 0 1228 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_124
timestamp 1710899220
transform 1 0 1172 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_125
timestamp 1710899220
transform 1 0 1164 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_126
timestamp 1710899220
transform 1 0 932 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_127
timestamp 1710899220
transform 1 0 1292 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_128
timestamp 1710899220
transform 1 0 1012 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_129
timestamp 1710899220
transform 1 0 1308 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_130
timestamp 1710899220
transform 1 0 1140 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_131
timestamp 1710899220
transform 1 0 1444 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_132
timestamp 1710899220
transform 1 0 1372 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_133
timestamp 1710899220
transform 1 0 1204 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_134
timestamp 1710899220
transform 1 0 1628 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_135
timestamp 1710899220
transform 1 0 1492 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_136
timestamp 1710899220
transform 1 0 1564 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_137
timestamp 1710899220
transform 1 0 1460 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_138
timestamp 1710899220
transform 1 0 1388 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_139
timestamp 1710899220
transform 1 0 1748 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_140
timestamp 1710899220
transform 1 0 1668 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_141
timestamp 1710899220
transform 1 0 1708 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_142
timestamp 1710899220
transform 1 0 1460 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_143
timestamp 1710899220
transform 1 0 1436 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_144
timestamp 1710899220
transform 1 0 1396 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_145
timestamp 1710899220
transform 1 0 1332 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_146
timestamp 1710899220
transform 1 0 1676 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_147
timestamp 1710899220
transform 1 0 1460 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_148
timestamp 1710899220
transform 1 0 1420 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_149
timestamp 1710899220
transform 1 0 1372 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_150
timestamp 1710899220
transform 1 0 1356 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_151
timestamp 1710899220
transform 1 0 1652 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_152
timestamp 1710899220
transform 1 0 1636 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_153
timestamp 1710899220
transform 1 0 1556 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_154
timestamp 1710899220
transform 1 0 1556 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_155
timestamp 1710899220
transform 1 0 1540 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_156
timestamp 1710899220
transform 1 0 1588 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_157
timestamp 1710899220
transform 1 0 1548 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_158
timestamp 1710899220
transform 1 0 1524 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_159
timestamp 1710899220
transform 1 0 1508 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_160
timestamp 1710899220
transform 1 0 1444 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_161
timestamp 1710899220
transform 1 0 1436 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_162
timestamp 1710899220
transform 1 0 1420 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_163
timestamp 1710899220
transform 1 0 1364 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_164
timestamp 1710899220
transform 1 0 1364 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_165
timestamp 1710899220
transform 1 0 1324 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_166
timestamp 1710899220
transform 1 0 1324 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_167
timestamp 1710899220
transform 1 0 804 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_168
timestamp 1710899220
transform 1 0 740 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_169
timestamp 1710899220
transform 1 0 732 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_170
timestamp 1710899220
transform 1 0 660 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_171
timestamp 1710899220
transform 1 0 628 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_172
timestamp 1710899220
transform 1 0 596 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_173
timestamp 1710899220
transform 1 0 596 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_174
timestamp 1710899220
transform 1 0 572 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_175
timestamp 1710899220
transform 1 0 1196 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_176
timestamp 1710899220
transform 1 0 1172 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_177
timestamp 1710899220
transform 1 0 1332 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_178
timestamp 1710899220
transform 1 0 1324 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_179
timestamp 1710899220
transform 1 0 1220 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_180
timestamp 1710899220
transform 1 0 1092 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_181
timestamp 1710899220
transform 1 0 1092 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_182
timestamp 1710899220
transform 1 0 732 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_183
timestamp 1710899220
transform 1 0 1356 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_184
timestamp 1710899220
transform 1 0 1300 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_185
timestamp 1710899220
transform 1 0 1340 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_186
timestamp 1710899220
transform 1 0 1292 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_187
timestamp 1710899220
transform 1 0 1332 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_188
timestamp 1710899220
transform 1 0 1324 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_189
timestamp 1710899220
transform 1 0 1292 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_190
timestamp 1710899220
transform 1 0 1292 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_191
timestamp 1710899220
transform 1 0 1252 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_192
timestamp 1710899220
transform 1 0 1244 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_193
timestamp 1710899220
transform 1 0 1100 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_194
timestamp 1710899220
transform 1 0 964 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_195
timestamp 1710899220
transform 1 0 764 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_196
timestamp 1710899220
transform 1 0 1364 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_197
timestamp 1710899220
transform 1 0 1356 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_198
timestamp 1710899220
transform 1 0 1196 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_199
timestamp 1710899220
transform 1 0 1188 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_200
timestamp 1710899220
transform 1 0 1068 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_201
timestamp 1710899220
transform 1 0 884 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_202
timestamp 1710899220
transform 1 0 788 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_203
timestamp 1710899220
transform 1 0 1380 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_204
timestamp 1710899220
transform 1 0 1348 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_205
timestamp 1710899220
transform 1 0 1308 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_206
timestamp 1710899220
transform 1 0 1140 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_207
timestamp 1710899220
transform 1 0 1100 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_208
timestamp 1710899220
transform 1 0 1052 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_209
timestamp 1710899220
transform 1 0 788 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_210
timestamp 1710899220
transform 1 0 1028 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_211
timestamp 1710899220
transform 1 0 980 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_212
timestamp 1710899220
transform 1 0 956 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_213
timestamp 1710899220
transform 1 0 956 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_214
timestamp 1710899220
transform 1 0 900 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_215
timestamp 1710899220
transform 1 0 796 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_216
timestamp 1710899220
transform 1 0 780 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_217
timestamp 1710899220
transform 1 0 732 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_218
timestamp 1710899220
transform 1 0 1260 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_219
timestamp 1710899220
transform 1 0 1236 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_220
timestamp 1710899220
transform 1 0 804 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_221
timestamp 1710899220
transform 1 0 2124 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_222
timestamp 1710899220
transform 1 0 2092 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_223
timestamp 1710899220
transform 1 0 1380 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_224
timestamp 1710899220
transform 1 0 1268 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_225
timestamp 1710899220
transform 1 0 1212 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_226
timestamp 1710899220
transform 1 0 1052 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_227
timestamp 1710899220
transform 1 0 732 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_228
timestamp 1710899220
transform 1 0 1500 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_229
timestamp 1710899220
transform 1 0 1180 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_230
timestamp 1710899220
transform 1 0 1140 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_231
timestamp 1710899220
transform 1 0 684 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_232
timestamp 1710899220
transform 1 0 684 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_233
timestamp 1710899220
transform 1 0 660 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_234
timestamp 1710899220
transform 1 0 1132 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_235
timestamp 1710899220
transform 1 0 1052 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_236
timestamp 1710899220
transform 1 0 980 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_237
timestamp 1710899220
transform 1 0 828 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_238
timestamp 1710899220
transform 1 0 508 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_239
timestamp 1710899220
transform 1 0 996 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_240
timestamp 1710899220
transform 1 0 836 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_241
timestamp 1710899220
transform 1 0 652 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_242
timestamp 1710899220
transform 1 0 428 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_243
timestamp 1710899220
transform 1 0 252 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_244
timestamp 1710899220
transform 1 0 1676 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_245
timestamp 1710899220
transform 1 0 1644 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_246
timestamp 1710899220
transform 1 0 1604 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_247
timestamp 1710899220
transform 1 0 1540 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_248
timestamp 1710899220
transform 1 0 2020 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_249
timestamp 1710899220
transform 1 0 1972 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_250
timestamp 1710899220
transform 1 0 1900 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_251
timestamp 1710899220
transform 1 0 1748 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_252
timestamp 1710899220
transform 1 0 1548 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_253
timestamp 1710899220
transform 1 0 1068 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_254
timestamp 1710899220
transform 1 0 1916 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_255
timestamp 1710899220
transform 1 0 1828 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_256
timestamp 1710899220
transform 1 0 1796 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_257
timestamp 1710899220
transform 1 0 1956 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_258
timestamp 1710899220
transform 1 0 1956 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_259
timestamp 1710899220
transform 1 0 1932 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_260
timestamp 1710899220
transform 1 0 1932 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_261
timestamp 1710899220
transform 1 0 1932 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_262
timestamp 1710899220
transform 1 0 1924 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_263
timestamp 1710899220
transform 1 0 1884 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_264
timestamp 1710899220
transform 1 0 1884 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_265
timestamp 1710899220
transform 1 0 1812 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_266
timestamp 1710899220
transform 1 0 1804 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_267
timestamp 1710899220
transform 1 0 1012 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_268
timestamp 1710899220
transform 1 0 980 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_269
timestamp 1710899220
transform 1 0 1004 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_270
timestamp 1710899220
transform 1 0 932 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_271
timestamp 1710899220
transform 1 0 1148 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_272
timestamp 1710899220
transform 1 0 1148 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_273
timestamp 1710899220
transform 1 0 1100 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_274
timestamp 1710899220
transform 1 0 1100 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_275
timestamp 1710899220
transform 1 0 1052 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_276
timestamp 1710899220
transform 1 0 1044 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_277
timestamp 1710899220
transform 1 0 1044 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_278
timestamp 1710899220
transform 1 0 1044 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_279
timestamp 1710899220
transform 1 0 996 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_280
timestamp 1710899220
transform 1 0 972 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_281
timestamp 1710899220
transform 1 0 1948 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_282
timestamp 1710899220
transform 1 0 1884 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_283
timestamp 1710899220
transform 1 0 1868 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_284
timestamp 1710899220
transform 1 0 1620 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_285
timestamp 1710899220
transform 1 0 1652 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_286
timestamp 1710899220
transform 1 0 1620 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_287
timestamp 1710899220
transform 1 0 1620 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_288
timestamp 1710899220
transform 1 0 1476 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_289
timestamp 1710899220
transform 1 0 1308 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_290
timestamp 1710899220
transform 1 0 1308 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_291
timestamp 1710899220
transform 1 0 836 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_292
timestamp 1710899220
transform 1 0 788 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_293
timestamp 1710899220
transform 1 0 788 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_294
timestamp 1710899220
transform 1 0 780 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_295
timestamp 1710899220
transform 1 0 764 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_296
timestamp 1710899220
transform 1 0 1148 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_297
timestamp 1710899220
transform 1 0 924 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_298
timestamp 1710899220
transform 1 0 884 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_299
timestamp 1710899220
transform 1 0 876 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_300
timestamp 1710899220
transform 1 0 868 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_301
timestamp 1710899220
transform 1 0 484 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_302
timestamp 1710899220
transform 1 0 276 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_303
timestamp 1710899220
transform 1 0 220 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_304
timestamp 1710899220
transform 1 0 732 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_305
timestamp 1710899220
transform 1 0 572 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_306
timestamp 1710899220
transform 1 0 796 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_307
timestamp 1710899220
transform 1 0 772 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_308
timestamp 1710899220
transform 1 0 756 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_309
timestamp 1710899220
transform 1 0 732 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_310
timestamp 1710899220
transform 1 0 692 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_311
timestamp 1710899220
transform 1 0 692 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_312
timestamp 1710899220
transform 1 0 516 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_313
timestamp 1710899220
transform 1 0 708 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_314
timestamp 1710899220
transform 1 0 684 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_315
timestamp 1710899220
transform 1 0 1020 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_316
timestamp 1710899220
transform 1 0 1012 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_317
timestamp 1710899220
transform 1 0 988 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_318
timestamp 1710899220
transform 1 0 980 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_319
timestamp 1710899220
transform 1 0 948 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_320
timestamp 1710899220
transform 1 0 940 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_321
timestamp 1710899220
transform 1 0 796 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_322
timestamp 1710899220
transform 1 0 748 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_323
timestamp 1710899220
transform 1 0 628 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_324
timestamp 1710899220
transform 1 0 628 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_325
timestamp 1710899220
transform 1 0 548 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_326
timestamp 1710899220
transform 1 0 804 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_327
timestamp 1710899220
transform 1 0 772 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_328
timestamp 1710899220
transform 1 0 740 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_329
timestamp 1710899220
transform 1 0 740 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_330
timestamp 1710899220
transform 1 0 724 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_331
timestamp 1710899220
transform 1 0 508 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_332
timestamp 1710899220
transform 1 0 252 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_333
timestamp 1710899220
transform 1 0 204 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_334
timestamp 1710899220
transform 1 0 196 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_335
timestamp 1710899220
transform 1 0 180 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_336
timestamp 1710899220
transform 1 0 156 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_337
timestamp 1710899220
transform 1 0 148 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_338
timestamp 1710899220
transform 1 0 812 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_339
timestamp 1710899220
transform 1 0 764 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_340
timestamp 1710899220
transform 1 0 1636 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_341
timestamp 1710899220
transform 1 0 1180 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_342
timestamp 1710899220
transform 1 0 1132 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_343
timestamp 1710899220
transform 1 0 908 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_344
timestamp 1710899220
transform 1 0 884 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_345
timestamp 1710899220
transform 1 0 876 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_346
timestamp 1710899220
transform 1 0 1780 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_347
timestamp 1710899220
transform 1 0 1716 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_348
timestamp 1710899220
transform 1 0 1708 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_349
timestamp 1710899220
transform 1 0 1684 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_350
timestamp 1710899220
transform 1 0 2020 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_351
timestamp 1710899220
transform 1 0 1988 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_352
timestamp 1710899220
transform 1 0 1332 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_353
timestamp 1710899220
transform 1 0 1268 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_354
timestamp 1710899220
transform 1 0 1228 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_355
timestamp 1710899220
transform 1 0 1180 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_356
timestamp 1710899220
transform 1 0 1140 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_357
timestamp 1710899220
transform 1 0 1004 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_358
timestamp 1710899220
transform 1 0 964 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_359
timestamp 1710899220
transform 1 0 948 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_360
timestamp 1710899220
transform 1 0 948 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_361
timestamp 1710899220
transform 1 0 932 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_362
timestamp 1710899220
transform 1 0 932 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_363
timestamp 1710899220
transform 1 0 780 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_364
timestamp 1710899220
transform 1 0 740 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_365
timestamp 1710899220
transform 1 0 724 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_366
timestamp 1710899220
transform 1 0 716 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_367
timestamp 1710899220
transform 1 0 980 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_368
timestamp 1710899220
transform 1 0 980 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_369
timestamp 1710899220
transform 1 0 932 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_370
timestamp 1710899220
transform 1 0 932 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_371
timestamp 1710899220
transform 1 0 892 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_372
timestamp 1710899220
transform 1 0 804 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_373
timestamp 1710899220
transform 1 0 692 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_374
timestamp 1710899220
transform 1 0 1340 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_375
timestamp 1710899220
transform 1 0 1324 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_376
timestamp 1710899220
transform 1 0 1292 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_377
timestamp 1710899220
transform 1 0 1180 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_378
timestamp 1710899220
transform 1 0 1164 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_379
timestamp 1710899220
transform 1 0 1132 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_380
timestamp 1710899220
transform 1 0 1116 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_381
timestamp 1710899220
transform 1 0 1100 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_382
timestamp 1710899220
transform 1 0 1084 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_383
timestamp 1710899220
transform 1 0 1076 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_384
timestamp 1710899220
transform 1 0 1012 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_385
timestamp 1710899220
transform 1 0 1004 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_386
timestamp 1710899220
transform 1 0 1004 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_387
timestamp 1710899220
transform 1 0 996 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_388
timestamp 1710899220
transform 1 0 964 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_389
timestamp 1710899220
transform 1 0 684 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_390
timestamp 1710899220
transform 1 0 644 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_391
timestamp 1710899220
transform 1 0 612 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_392
timestamp 1710899220
transform 1 0 524 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_393
timestamp 1710899220
transform 1 0 1156 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_394
timestamp 1710899220
transform 1 0 1092 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_395
timestamp 1710899220
transform 1 0 1084 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_396
timestamp 1710899220
transform 1 0 1060 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_397
timestamp 1710899220
transform 1 0 892 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_398
timestamp 1710899220
transform 1 0 788 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_399
timestamp 1710899220
transform 1 0 788 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_400
timestamp 1710899220
transform 1 0 668 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_401
timestamp 1710899220
transform 1 0 660 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_402
timestamp 1710899220
transform 1 0 636 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_403
timestamp 1710899220
transform 1 0 628 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_404
timestamp 1710899220
transform 1 0 340 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_405
timestamp 1710899220
transform 1 0 308 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_406
timestamp 1710899220
transform 1 0 244 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_407
timestamp 1710899220
transform 1 0 188 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_408
timestamp 1710899220
transform 1 0 476 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_409
timestamp 1710899220
transform 1 0 444 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_410
timestamp 1710899220
transform 1 0 244 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_411
timestamp 1710899220
transform 1 0 196 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_412
timestamp 1710899220
transform 1 0 148 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_413
timestamp 1710899220
transform 1 0 1020 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_414
timestamp 1710899220
transform 1 0 940 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_415
timestamp 1710899220
transform 1 0 940 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_416
timestamp 1710899220
transform 1 0 900 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_417
timestamp 1710899220
transform 1 0 1076 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_418
timestamp 1710899220
transform 1 0 1052 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_419
timestamp 1710899220
transform 1 0 1724 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_420
timestamp 1710899220
transform 1 0 1676 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_421
timestamp 1710899220
transform 1 0 1676 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_422
timestamp 1710899220
transform 1 0 1644 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_423
timestamp 1710899220
transform 1 0 1596 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_424
timestamp 1710899220
transform 1 0 1348 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_425
timestamp 1710899220
transform 1 0 1228 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_426
timestamp 1710899220
transform 1 0 1196 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_427
timestamp 1710899220
transform 1 0 1308 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_428
timestamp 1710899220
transform 1 0 1276 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_429
timestamp 1710899220
transform 1 0 1252 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_430
timestamp 1710899220
transform 1 0 1244 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_431
timestamp 1710899220
transform 1 0 1084 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_432
timestamp 1710899220
transform 1 0 1084 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_433
timestamp 1710899220
transform 1 0 732 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_434
timestamp 1710899220
transform 1 0 732 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_435
timestamp 1710899220
transform 1 0 692 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_436
timestamp 1710899220
transform 1 0 708 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_437
timestamp 1710899220
transform 1 0 668 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_438
timestamp 1710899220
transform 1 0 548 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_439
timestamp 1710899220
transform 1 0 372 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_440
timestamp 1710899220
transform 1 0 548 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_441
timestamp 1710899220
transform 1 0 500 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_442
timestamp 1710899220
transform 1 0 396 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_443
timestamp 1710899220
transform 1 0 332 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_444
timestamp 1710899220
transform 1 0 556 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_445
timestamp 1710899220
transform 1 0 548 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_446
timestamp 1710899220
transform 1 0 524 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_447
timestamp 1710899220
transform 1 0 500 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_448
timestamp 1710899220
transform 1 0 340 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_449
timestamp 1710899220
transform 1 0 300 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_450
timestamp 1710899220
transform 1 0 1148 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_451
timestamp 1710899220
transform 1 0 1084 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_452
timestamp 1710899220
transform 1 0 1020 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_453
timestamp 1710899220
transform 1 0 1020 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_454
timestamp 1710899220
transform 1 0 964 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_455
timestamp 1710899220
transform 1 0 844 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_456
timestamp 1710899220
transform 1 0 804 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_457
timestamp 1710899220
transform 1 0 756 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_458
timestamp 1710899220
transform 1 0 836 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_459
timestamp 1710899220
transform 1 0 756 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_460
timestamp 1710899220
transform 1 0 580 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_461
timestamp 1710899220
transform 1 0 836 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_462
timestamp 1710899220
transform 1 0 652 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_463
timestamp 1710899220
transform 1 0 372 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_464
timestamp 1710899220
transform 1 0 1388 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_465
timestamp 1710899220
transform 1 0 1140 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_466
timestamp 1710899220
transform 1 0 1140 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_467
timestamp 1710899220
transform 1 0 1060 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_468
timestamp 1710899220
transform 1 0 1060 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_469
timestamp 1710899220
transform 1 0 796 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_470
timestamp 1710899220
transform 1 0 396 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_471
timestamp 1710899220
transform 1 0 1036 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_472
timestamp 1710899220
transform 1 0 988 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_473
timestamp 1710899220
transform 1 0 972 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_474
timestamp 1710899220
transform 1 0 972 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_475
timestamp 1710899220
transform 1 0 908 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_476
timestamp 1710899220
transform 1 0 1276 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_477
timestamp 1710899220
transform 1 0 1140 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_478
timestamp 1710899220
transform 1 0 1300 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_479
timestamp 1710899220
transform 1 0 1268 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_480
timestamp 1710899220
transform 1 0 1196 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_481
timestamp 1710899220
transform 1 0 1180 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_482
timestamp 1710899220
transform 1 0 1684 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_483
timestamp 1710899220
transform 1 0 1636 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_484
timestamp 1710899220
transform 1 0 1564 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_485
timestamp 1710899220
transform 1 0 1564 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_486
timestamp 1710899220
transform 1 0 1412 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_487
timestamp 1710899220
transform 1 0 1284 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_488
timestamp 1710899220
transform 1 0 1620 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_489
timestamp 1710899220
transform 1 0 1620 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_490
timestamp 1710899220
transform 1 0 1604 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_491
timestamp 1710899220
transform 1 0 1484 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_492
timestamp 1710899220
transform 1 0 1484 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_493
timestamp 1710899220
transform 1 0 1380 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_494
timestamp 1710899220
transform 1 0 1684 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_495
timestamp 1710899220
transform 1 0 1660 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_496
timestamp 1710899220
transform 1 0 1452 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_497
timestamp 1710899220
transform 1 0 1396 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_498
timestamp 1710899220
transform 1 0 1380 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_499
timestamp 1710899220
transform 1 0 2012 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_500
timestamp 1710899220
transform 1 0 1956 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_501
timestamp 1710899220
transform 1 0 1844 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_502
timestamp 1710899220
transform 1 0 1844 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_503
timestamp 1710899220
transform 1 0 1804 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_504
timestamp 1710899220
transform 1 0 1788 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_505
timestamp 1710899220
transform 1 0 1772 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_506
timestamp 1710899220
transform 1 0 2004 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_507
timestamp 1710899220
transform 1 0 1964 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_508
timestamp 1710899220
transform 1 0 1948 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_509
timestamp 1710899220
transform 1 0 1812 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_510
timestamp 1710899220
transform 1 0 1836 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_511
timestamp 1710899220
transform 1 0 1724 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_512
timestamp 1710899220
transform 1 0 1716 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_513
timestamp 1710899220
transform 1 0 1676 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_514
timestamp 1710899220
transform 1 0 2012 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_515
timestamp 1710899220
transform 1 0 1980 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_516
timestamp 1710899220
transform 1 0 1820 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_517
timestamp 1710899220
transform 1 0 1820 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_518
timestamp 1710899220
transform 1 0 1788 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_519
timestamp 1710899220
transform 1 0 1644 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_520
timestamp 1710899220
transform 1 0 1556 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_521
timestamp 1710899220
transform 1 0 1556 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_522
timestamp 1710899220
transform 1 0 1508 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_523
timestamp 1710899220
transform 1 0 1508 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_524
timestamp 1710899220
transform 1 0 1396 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_525
timestamp 1710899220
transform 1 0 1804 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_526
timestamp 1710899220
transform 1 0 1516 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_527
timestamp 1710899220
transform 1 0 1460 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_528
timestamp 1710899220
transform 1 0 1460 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_529
timestamp 1710899220
transform 1 0 1396 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_530
timestamp 1710899220
transform 1 0 1684 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_531
timestamp 1710899220
transform 1 0 1660 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_532
timestamp 1710899220
transform 1 0 1644 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_533
timestamp 1710899220
transform 1 0 1876 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_534
timestamp 1710899220
transform 1 0 1820 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_535
timestamp 1710899220
transform 1 0 1820 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_536
timestamp 1710899220
transform 1 0 1772 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_537
timestamp 1710899220
transform 1 0 1772 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_538
timestamp 1710899220
transform 1 0 1748 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_539
timestamp 1710899220
transform 1 0 1628 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_540
timestamp 1710899220
transform 1 0 1524 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_541
timestamp 1710899220
transform 1 0 1980 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_542
timestamp 1710899220
transform 1 0 1948 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_543
timestamp 1710899220
transform 1 0 1828 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_544
timestamp 1710899220
transform 1 0 1828 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_545
timestamp 1710899220
transform 1 0 1764 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_546
timestamp 1710899220
transform 1 0 1764 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_547
timestamp 1710899220
transform 1 0 1988 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_548
timestamp 1710899220
transform 1 0 1956 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_549
timestamp 1710899220
transform 1 0 1932 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_550
timestamp 1710899220
transform 1 0 1820 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_551
timestamp 1710899220
transform 1 0 1796 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_552
timestamp 1710899220
transform 1 0 1740 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_553
timestamp 1710899220
transform 1 0 1516 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_554
timestamp 1710899220
transform 1 0 1436 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_555
timestamp 1710899220
transform 1 0 2028 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_556
timestamp 1710899220
transform 1 0 1860 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_557
timestamp 1710899220
transform 1 0 1788 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_558
timestamp 1710899220
transform 1 0 1780 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_559
timestamp 1710899220
transform 1 0 1564 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_560
timestamp 1710899220
transform 1 0 1564 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_561
timestamp 1710899220
transform 1 0 1524 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_562
timestamp 1710899220
transform 1 0 1500 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_563
timestamp 1710899220
transform 1 0 1500 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_564
timestamp 1710899220
transform 1 0 1500 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_565
timestamp 1710899220
transform 1 0 1420 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_566
timestamp 1710899220
transform 1 0 1596 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_567
timestamp 1710899220
transform 1 0 1532 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_568
timestamp 1710899220
transform 1 0 1556 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_569
timestamp 1710899220
transform 1 0 1492 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_570
timestamp 1710899220
transform 1 0 740 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_571
timestamp 1710899220
transform 1 0 692 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_572
timestamp 1710899220
transform 1 0 348 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_573
timestamp 1710899220
transform 1 0 308 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_574
timestamp 1710899220
transform 1 0 324 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_575
timestamp 1710899220
transform 1 0 284 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_576
timestamp 1710899220
transform 1 0 844 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_577
timestamp 1710899220
transform 1 0 788 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_578
timestamp 1710899220
transform 1 0 348 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_579
timestamp 1710899220
transform 1 0 308 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_580
timestamp 1710899220
transform 1 0 412 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_581
timestamp 1710899220
transform 1 0 388 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_582
timestamp 1710899220
transform 1 0 364 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_583
timestamp 1710899220
transform 1 0 1012 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_584
timestamp 1710899220
transform 1 0 980 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_585
timestamp 1710899220
transform 1 0 1700 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_586
timestamp 1710899220
transform 1 0 1660 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_587
timestamp 1710899220
transform 1 0 1700 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_588
timestamp 1710899220
transform 1 0 1628 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_589
timestamp 1710899220
transform 1 0 2028 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_590
timestamp 1710899220
transform 1 0 1940 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_591
timestamp 1710899220
transform 1 0 1892 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_592
timestamp 1710899220
transform 1 0 2028 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_593
timestamp 1710899220
transform 1 0 2028 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_594
timestamp 1710899220
transform 1 0 1988 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_595
timestamp 1710899220
transform 1 0 1956 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_596
timestamp 1710899220
transform 1 0 1916 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_597
timestamp 1710899220
transform 1 0 2004 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_598
timestamp 1710899220
transform 1 0 1980 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_599
timestamp 1710899220
transform 1 0 1676 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_600
timestamp 1710899220
transform 1 0 1628 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_601
timestamp 1710899220
transform 1 0 1572 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_602
timestamp 1710899220
transform 1 0 1892 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_603
timestamp 1710899220
transform 1 0 1852 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_604
timestamp 1710899220
transform 1 0 1772 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_605
timestamp 1710899220
transform 1 0 1724 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_606
timestamp 1710899220
transform 1 0 1996 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_607
timestamp 1710899220
transform 1 0 1956 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_608
timestamp 1710899220
transform 1 0 2004 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_609
timestamp 1710899220
transform 1 0 1956 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_610
timestamp 1710899220
transform 1 0 1924 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_611
timestamp 1710899220
transform 1 0 2052 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_612
timestamp 1710899220
transform 1 0 2012 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_613
timestamp 1710899220
transform 1 0 2012 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_614
timestamp 1710899220
transform 1 0 1908 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_615
timestamp 1710899220
transform 1 0 1852 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_616
timestamp 1710899220
transform 1 0 2316 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_617
timestamp 1710899220
transform 1 0 2268 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_618
timestamp 1710899220
transform 1 0 2532 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_619
timestamp 1710899220
transform 1 0 2476 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_620
timestamp 1710899220
transform 1 0 2476 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_621
timestamp 1710899220
transform 1 0 2396 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_622
timestamp 1710899220
transform 1 0 2348 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_623
timestamp 1710899220
transform 1 0 2508 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_624
timestamp 1710899220
transform 1 0 2412 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_625
timestamp 1710899220
transform 1 0 2484 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_626
timestamp 1710899220
transform 1 0 2396 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_627
timestamp 1710899220
transform 1 0 2316 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_628
timestamp 1710899220
transform 1 0 2572 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_629
timestamp 1710899220
transform 1 0 2532 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_630
timestamp 1710899220
transform 1 0 2500 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_631
timestamp 1710899220
transform 1 0 2468 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_632
timestamp 1710899220
transform 1 0 2572 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_633
timestamp 1710899220
transform 1 0 2516 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_634
timestamp 1710899220
transform 1 0 2548 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_635
timestamp 1710899220
transform 1 0 2436 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_636
timestamp 1710899220
transform 1 0 2372 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_637
timestamp 1710899220
transform 1 0 2332 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_638
timestamp 1710899220
transform 1 0 2276 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_639
timestamp 1710899220
transform 1 0 2548 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_640
timestamp 1710899220
transform 1 0 2404 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_641
timestamp 1710899220
transform 1 0 2628 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_642
timestamp 1710899220
transform 1 0 2404 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_643
timestamp 1710899220
transform 1 0 2468 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_644
timestamp 1710899220
transform 1 0 2412 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_645
timestamp 1710899220
transform 1 0 2340 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_646
timestamp 1710899220
transform 1 0 2292 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_647
timestamp 1710899220
transform 1 0 2324 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_648
timestamp 1710899220
transform 1 0 2324 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_649
timestamp 1710899220
transform 1 0 2292 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_650
timestamp 1710899220
transform 1 0 2260 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_651
timestamp 1710899220
transform 1 0 2252 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_652
timestamp 1710899220
transform 1 0 2236 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_653
timestamp 1710899220
transform 1 0 2060 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_654
timestamp 1710899220
transform 1 0 2276 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_655
timestamp 1710899220
transform 1 0 2236 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_656
timestamp 1710899220
transform 1 0 2188 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_657
timestamp 1710899220
transform 1 0 2132 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_658
timestamp 1710899220
transform 1 0 2196 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_659
timestamp 1710899220
transform 1 0 2180 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_660
timestamp 1710899220
transform 1 0 2484 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_661
timestamp 1710899220
transform 1 0 2460 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_662
timestamp 1710899220
transform 1 0 1260 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_663
timestamp 1710899220
transform 1 0 1156 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_664
timestamp 1710899220
transform 1 0 1028 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_665
timestamp 1710899220
transform 1 0 948 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_666
timestamp 1710899220
transform 1 0 1156 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_667
timestamp 1710899220
transform 1 0 1004 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_668
timestamp 1710899220
transform 1 0 900 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_669
timestamp 1710899220
transform 1 0 1092 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_670
timestamp 1710899220
transform 1 0 940 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_671
timestamp 1710899220
transform 1 0 852 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_672
timestamp 1710899220
transform 1 0 852 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_673
timestamp 1710899220
transform 1 0 668 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_674
timestamp 1710899220
transform 1 0 668 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_675
timestamp 1710899220
transform 1 0 516 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_676
timestamp 1710899220
transform 1 0 716 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_677
timestamp 1710899220
transform 1 0 524 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_678
timestamp 1710899220
transform 1 0 524 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_679
timestamp 1710899220
transform 1 0 444 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_680
timestamp 1710899220
transform 1 0 292 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_681
timestamp 1710899220
transform 1 0 756 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_682
timestamp 1710899220
transform 1 0 700 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_683
timestamp 1710899220
transform 1 0 484 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_684
timestamp 1710899220
transform 1 0 268 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_685
timestamp 1710899220
transform 1 0 228 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_686
timestamp 1710899220
transform 1 0 148 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_687
timestamp 1710899220
transform 1 0 356 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_688
timestamp 1710899220
transform 1 0 268 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_689
timestamp 1710899220
transform 1 0 484 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_690
timestamp 1710899220
transform 1 0 396 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_691
timestamp 1710899220
transform 1 0 396 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_692
timestamp 1710899220
transform 1 0 292 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_693
timestamp 1710899220
transform 1 0 588 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_694
timestamp 1710899220
transform 1 0 476 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_695
timestamp 1710899220
transform 1 0 660 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_696
timestamp 1710899220
transform 1 0 572 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_697
timestamp 1710899220
transform 1 0 908 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_698
timestamp 1710899220
transform 1 0 860 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_699
timestamp 1710899220
transform 1 0 780 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_700
timestamp 1710899220
transform 1 0 788 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_701
timestamp 1710899220
transform 1 0 700 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_702
timestamp 1710899220
transform 1 0 980 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_703
timestamp 1710899220
transform 1 0 892 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_704
timestamp 1710899220
transform 1 0 1164 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_705
timestamp 1710899220
transform 1 0 1076 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_706
timestamp 1710899220
transform 1 0 1116 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_707
timestamp 1710899220
transform 1 0 1020 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_708
timestamp 1710899220
transform 1 0 1020 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_709
timestamp 1710899220
transform 1 0 860 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_710
timestamp 1710899220
transform 1 0 1460 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_711
timestamp 1710899220
transform 1 0 1372 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_712
timestamp 1710899220
transform 1 0 1356 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_713
timestamp 1710899220
transform 1 0 1316 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_714
timestamp 1710899220
transform 1 0 1588 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_715
timestamp 1710899220
transform 1 0 1500 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_716
timestamp 1710899220
transform 1 0 1332 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_717
timestamp 1710899220
transform 1 0 1780 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_718
timestamp 1710899220
transform 1 0 1692 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_719
timestamp 1710899220
transform 1 0 1580 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_720
timestamp 1710899220
transform 1 0 1420 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_721
timestamp 1710899220
transform 1 0 1692 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_722
timestamp 1710899220
transform 1 0 1604 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_723
timestamp 1710899220
transform 1 0 1812 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_724
timestamp 1710899220
transform 1 0 1708 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_725
timestamp 1710899220
transform 1 0 1740 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_726
timestamp 1710899220
transform 1 0 1668 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_727
timestamp 1710899220
transform 1 0 1644 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_728
timestamp 1710899220
transform 1 0 1612 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_729
timestamp 1710899220
transform 1 0 1564 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_730
timestamp 1710899220
transform 1 0 1532 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_731
timestamp 1710899220
transform 1 0 1468 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_732
timestamp 1710899220
transform 1 0 1660 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_733
timestamp 1710899220
transform 1 0 1644 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_734
timestamp 1710899220
transform 1 0 1468 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_735
timestamp 1710899220
transform 1 0 1428 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_736
timestamp 1710899220
transform 1 0 1348 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_737
timestamp 1710899220
transform 1 0 1268 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_738
timestamp 1710899220
transform 1 0 1516 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_739
timestamp 1710899220
transform 1 0 1500 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_740
timestamp 1710899220
transform 1 0 1316 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_741
timestamp 1710899220
transform 1 0 1316 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_742
timestamp 1710899220
transform 1 0 1316 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_743
timestamp 1710899220
transform 1 0 1292 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_744
timestamp 1710899220
transform 1 0 2236 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_745
timestamp 1710899220
transform 1 0 2212 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_746
timestamp 1710899220
transform 1 0 2508 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_747
timestamp 1710899220
transform 1 0 2468 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_748
timestamp 1710899220
transform 1 0 2628 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_749
timestamp 1710899220
transform 1 0 2588 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_750
timestamp 1710899220
transform 1 0 2324 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_751
timestamp 1710899220
transform 1 0 2284 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_752
timestamp 1710899220
transform 1 0 2324 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_753
timestamp 1710899220
transform 1 0 2284 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_754
timestamp 1710899220
transform 1 0 2596 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_755
timestamp 1710899220
transform 1 0 2556 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_756
timestamp 1710899220
transform 1 0 2612 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_757
timestamp 1710899220
transform 1 0 2572 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_758
timestamp 1710899220
transform 1 0 2460 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_759
timestamp 1710899220
transform 1 0 2420 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_760
timestamp 1710899220
transform 1 0 1916 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_761
timestamp 1710899220
transform 1 0 1876 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_762
timestamp 1710899220
transform 1 0 1924 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_763
timestamp 1710899220
transform 1 0 1876 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_764
timestamp 1710899220
transform 1 0 1916 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_765
timestamp 1710899220
transform 1 0 1876 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_766
timestamp 1710899220
transform 1 0 2284 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_767
timestamp 1710899220
transform 1 0 2236 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_768
timestamp 1710899220
transform 1 0 2132 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_769
timestamp 1710899220
transform 1 0 2084 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_770
timestamp 1710899220
transform 1 0 2260 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_771
timestamp 1710899220
transform 1 0 2212 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_772
timestamp 1710899220
transform 1 0 1812 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_773
timestamp 1710899220
transform 1 0 1796 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_774
timestamp 1710899220
transform 1 0 1460 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_775
timestamp 1710899220
transform 1 0 1308 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_776
timestamp 1710899220
transform 1 0 1156 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_777
timestamp 1710899220
transform 1 0 2092 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_778
timestamp 1710899220
transform 1 0 2052 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_779
timestamp 1710899220
transform 1 0 2268 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_780
timestamp 1710899220
transform 1 0 2172 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_781
timestamp 1710899220
transform 1 0 2116 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_782
timestamp 1710899220
transform 1 0 2116 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_783
timestamp 1710899220
transform 1 0 2052 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_784
timestamp 1710899220
transform 1 0 1180 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_785
timestamp 1710899220
transform 1 0 916 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_786
timestamp 1710899220
transform 1 0 868 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_787
timestamp 1710899220
transform 1 0 1092 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_788
timestamp 1710899220
transform 1 0 892 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_789
timestamp 1710899220
transform 1 0 1044 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_790
timestamp 1710899220
transform 1 0 948 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_791
timestamp 1710899220
transform 1 0 1748 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_792
timestamp 1710899220
transform 1 0 1732 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_793
timestamp 1710899220
transform 1 0 1068 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_794
timestamp 1710899220
transform 1 0 924 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_795
timestamp 1710899220
transform 1 0 1148 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_796
timestamp 1710899220
transform 1 0 1116 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_797
timestamp 1710899220
transform 1 0 1900 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_798
timestamp 1710899220
transform 1 0 1852 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_799
timestamp 1710899220
transform 1 0 1852 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_800
timestamp 1710899220
transform 1 0 1804 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_801
timestamp 1710899220
transform 1 0 1196 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_802
timestamp 1710899220
transform 1 0 1124 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_803
timestamp 1710899220
transform 1 0 1060 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_804
timestamp 1710899220
transform 1 0 988 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_805
timestamp 1710899220
transform 1 0 1836 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_806
timestamp 1710899220
transform 1 0 1796 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_807
timestamp 1710899220
transform 1 0 2588 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_808
timestamp 1710899220
transform 1 0 2572 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_809
timestamp 1710899220
transform 1 0 2540 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_810
timestamp 1710899220
transform 1 0 2476 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_811
timestamp 1710899220
transform 1 0 2444 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_812
timestamp 1710899220
transform 1 0 2420 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_813
timestamp 1710899220
transform 1 0 2396 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_814
timestamp 1710899220
transform 1 0 2340 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_815
timestamp 1710899220
transform 1 0 2292 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_816
timestamp 1710899220
transform 1 0 2284 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_817
timestamp 1710899220
transform 1 0 1980 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_818
timestamp 1710899220
transform 1 0 1892 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_819
timestamp 1710899220
transform 1 0 1844 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_820
timestamp 1710899220
transform 1 0 2588 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_821
timestamp 1710899220
transform 1 0 2572 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_822
timestamp 1710899220
transform 1 0 2564 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_823
timestamp 1710899220
transform 1 0 2436 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_824
timestamp 1710899220
transform 1 0 2420 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_825
timestamp 1710899220
transform 1 0 2308 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_826
timestamp 1710899220
transform 1 0 2284 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_827
timestamp 1710899220
transform 1 0 2236 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_828
timestamp 1710899220
transform 1 0 2236 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_829
timestamp 1710899220
transform 1 0 2348 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_830
timestamp 1710899220
transform 1 0 2252 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_831
timestamp 1710899220
transform 1 0 2212 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_832
timestamp 1710899220
transform 1 0 2164 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_833
timestamp 1710899220
transform 1 0 2124 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_834
timestamp 1710899220
transform 1 0 2068 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_835
timestamp 1710899220
transform 1 0 2036 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_836
timestamp 1710899220
transform 1 0 1996 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_837
timestamp 1710899220
transform 1 0 1964 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_838
timestamp 1710899220
transform 1 0 1844 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_839
timestamp 1710899220
transform 1 0 1828 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_840
timestamp 1710899220
transform 1 0 2068 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_841
timestamp 1710899220
transform 1 0 2044 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_842
timestamp 1710899220
transform 1 0 1956 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_843
timestamp 1710899220
transform 1 0 1916 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_844
timestamp 1710899220
transform 1 0 1724 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_845
timestamp 1710899220
transform 1 0 1676 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_846
timestamp 1710899220
transform 1 0 1676 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_847
timestamp 1710899220
transform 1 0 1572 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_848
timestamp 1710899220
transform 1 0 1564 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_849
timestamp 1710899220
transform 1 0 1236 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_850
timestamp 1710899220
transform 1 0 1172 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_851
timestamp 1710899220
transform 1 0 1172 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_852
timestamp 1710899220
transform 1 0 1156 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_853
timestamp 1710899220
transform 1 0 1060 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_854
timestamp 1710899220
transform 1 0 964 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_855
timestamp 1710899220
transform 1 0 964 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_856
timestamp 1710899220
transform 1 0 924 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_857
timestamp 1710899220
transform 1 0 924 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_858
timestamp 1710899220
transform 1 0 828 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_859
timestamp 1710899220
transform 1 0 596 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_860
timestamp 1710899220
transform 1 0 588 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_861
timestamp 1710899220
transform 1 0 452 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_862
timestamp 1710899220
transform 1 0 244 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_863
timestamp 1710899220
transform 1 0 244 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_864
timestamp 1710899220
transform 1 0 188 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_865
timestamp 1710899220
transform 1 0 180 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_866
timestamp 1710899220
transform 1 0 1972 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_867
timestamp 1710899220
transform 1 0 1860 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_868
timestamp 1710899220
transform 1 0 1844 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_869
timestamp 1710899220
transform 1 0 1772 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_870
timestamp 1710899220
transform 1 0 1564 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_871
timestamp 1710899220
transform 1 0 1524 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_872
timestamp 1710899220
transform 1 0 1516 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_873
timestamp 1710899220
transform 1 0 1468 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_874
timestamp 1710899220
transform 1 0 1468 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_875
timestamp 1710899220
transform 1 0 1460 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_876
timestamp 1710899220
transform 1 0 1436 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_877
timestamp 1710899220
transform 1 0 1436 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_878
timestamp 1710899220
transform 1 0 1364 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_879
timestamp 1710899220
transform 1 0 1364 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_880
timestamp 1710899220
transform 1 0 1324 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_881
timestamp 1710899220
transform 1 0 1268 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_882
timestamp 1710899220
transform 1 0 1260 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_883
timestamp 1710899220
transform 1 0 1212 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_884
timestamp 1710899220
transform 1 0 1212 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_885
timestamp 1710899220
transform 1 0 1172 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_886
timestamp 1710899220
transform 1 0 1164 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_887
timestamp 1710899220
transform 1 0 1164 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_888
timestamp 1710899220
transform 1 0 1116 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_889
timestamp 1710899220
transform 1 0 1076 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_890
timestamp 1710899220
transform 1 0 868 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_891
timestamp 1710899220
transform 1 0 860 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_892
timestamp 1710899220
transform 1 0 764 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_893
timestamp 1710899220
transform 1 0 748 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_894
timestamp 1710899220
transform 1 0 668 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_895
timestamp 1710899220
transform 1 0 588 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_896
timestamp 1710899220
transform 1 0 580 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_897
timestamp 1710899220
transform 1 0 564 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_898
timestamp 1710899220
transform 1 0 556 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_899
timestamp 1710899220
transform 1 0 452 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_900
timestamp 1710899220
transform 1 0 412 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_901
timestamp 1710899220
transform 1 0 2180 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_902
timestamp 1710899220
transform 1 0 2140 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_903
timestamp 1710899220
transform 1 0 2044 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_904
timestamp 1710899220
transform 1 0 1948 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_905
timestamp 1710899220
transform 1 0 1948 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_906
timestamp 1710899220
transform 1 0 1900 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_907
timestamp 1710899220
transform 1 0 1884 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_908
timestamp 1710899220
transform 1 0 1804 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_909
timestamp 1710899220
transform 1 0 1588 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_910
timestamp 1710899220
transform 1 0 1396 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_911
timestamp 1710899220
transform 1 0 1364 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_912
timestamp 1710899220
transform 1 0 1228 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_913
timestamp 1710899220
transform 1 0 1228 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_914
timestamp 1710899220
transform 1 0 1228 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_915
timestamp 1710899220
transform 1 0 1228 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_916
timestamp 1710899220
transform 1 0 1108 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_917
timestamp 1710899220
transform 1 0 1060 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_918
timestamp 1710899220
transform 1 0 1060 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_919
timestamp 1710899220
transform 1 0 1740 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_920
timestamp 1710899220
transform 1 0 1444 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_921
timestamp 1710899220
transform 1 0 1444 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_922
timestamp 1710899220
transform 1 0 1204 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_923
timestamp 1710899220
transform 1 0 1020 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_924
timestamp 1710899220
transform 1 0 940 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_925
timestamp 1710899220
transform 1 0 924 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_926
timestamp 1710899220
transform 1 0 884 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_927
timestamp 1710899220
transform 1 0 820 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_928
timestamp 1710899220
transform 1 0 804 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_929
timestamp 1710899220
transform 1 0 780 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_930
timestamp 1710899220
transform 1 0 756 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_931
timestamp 1710899220
transform 1 0 692 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_932
timestamp 1710899220
transform 1 0 540 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_933
timestamp 1710899220
transform 1 0 476 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_934
timestamp 1710899220
transform 1 0 1852 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_935
timestamp 1710899220
transform 1 0 1820 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_936
timestamp 1710899220
transform 1 0 1772 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_937
timestamp 1710899220
transform 1 0 1764 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_938
timestamp 1710899220
transform 1 0 1684 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_939
timestamp 1710899220
transform 1 0 1644 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_940
timestamp 1710899220
transform 1 0 1604 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_941
timestamp 1710899220
transform 1 0 1444 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_942
timestamp 1710899220
transform 1 0 1412 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_943
timestamp 1710899220
transform 1 0 1236 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_944
timestamp 1710899220
transform 1 0 1140 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_945
timestamp 1710899220
transform 1 0 1036 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_946
timestamp 1710899220
transform 1 0 996 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_947
timestamp 1710899220
transform 1 0 2268 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_948
timestamp 1710899220
transform 1 0 2060 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_949
timestamp 1710899220
transform 1 0 2028 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_950
timestamp 1710899220
transform 1 0 1772 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_951
timestamp 1710899220
transform 1 0 1316 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_952
timestamp 1710899220
transform 1 0 1300 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_953
timestamp 1710899220
transform 1 0 1244 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_954
timestamp 1710899220
transform 1 0 1220 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_955
timestamp 1710899220
transform 1 0 1844 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_956
timestamp 1710899220
transform 1 0 1804 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_957
timestamp 1710899220
transform 1 0 1476 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_958
timestamp 1710899220
transform 1 0 1452 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_959
timestamp 1710899220
transform 1 0 1452 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_960
timestamp 1710899220
transform 1 0 1428 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_961
timestamp 1710899220
transform 1 0 1428 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_962
timestamp 1710899220
transform 1 0 1428 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_963
timestamp 1710899220
transform 1 0 1420 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_964
timestamp 1710899220
transform 1 0 1420 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_965
timestamp 1710899220
transform 1 0 1404 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_966
timestamp 1710899220
transform 1 0 1396 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_967
timestamp 1710899220
transform 1 0 1364 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_968
timestamp 1710899220
transform 1 0 1332 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_969
timestamp 1710899220
transform 1 0 1324 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_970
timestamp 1710899220
transform 1 0 1284 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_971
timestamp 1710899220
transform 1 0 1260 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_972
timestamp 1710899220
transform 1 0 1220 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_973
timestamp 1710899220
transform 1 0 1124 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_974
timestamp 1710899220
transform 1 0 1004 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_975
timestamp 1710899220
transform 1 0 876 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_976
timestamp 1710899220
transform 1 0 836 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_977
timestamp 1710899220
transform 1 0 756 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_978
timestamp 1710899220
transform 1 0 724 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_979
timestamp 1710899220
transform 1 0 700 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_980
timestamp 1710899220
transform 1 0 684 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_981
timestamp 1710899220
transform 1 0 676 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_982
timestamp 1710899220
transform 1 0 660 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_983
timestamp 1710899220
transform 1 0 1812 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_984
timestamp 1710899220
transform 1 0 1812 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_985
timestamp 1710899220
transform 1 0 1772 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_986
timestamp 1710899220
transform 1 0 1764 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_987
timestamp 1710899220
transform 1 0 1764 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_988
timestamp 1710899220
transform 1 0 1548 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_989
timestamp 1710899220
transform 1 0 1548 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_990
timestamp 1710899220
transform 1 0 1532 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_991
timestamp 1710899220
transform 1 0 1492 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_992
timestamp 1710899220
transform 1 0 1492 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_993
timestamp 1710899220
transform 1 0 1484 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_994
timestamp 1710899220
transform 1 0 1420 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_995
timestamp 1710899220
transform 1 0 1404 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_996
timestamp 1710899220
transform 1 0 1396 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_997
timestamp 1710899220
transform 1 0 1324 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_998
timestamp 1710899220
transform 1 0 1260 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_999
timestamp 1710899220
transform 1 0 1172 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_1000
timestamp 1710899220
transform 1 0 1100 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1001
timestamp 1710899220
transform 1 0 972 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1002
timestamp 1710899220
transform 1 0 972 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_1003
timestamp 1710899220
transform 1 0 868 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1004
timestamp 1710899220
transform 1 0 812 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_1005
timestamp 1710899220
transform 1 0 812 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1006
timestamp 1710899220
transform 1 0 668 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_1007
timestamp 1710899220
transform 1 0 668 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_1008
timestamp 1710899220
transform 1 0 612 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_1009
timestamp 1710899220
transform 1 0 540 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_1010
timestamp 1710899220
transform 1 0 1148 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_1011
timestamp 1710899220
transform 1 0 1124 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1012
timestamp 1710899220
transform 1 0 1092 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_1013
timestamp 1710899220
transform 1 0 996 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1014
timestamp 1710899220
transform 1 0 964 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1015
timestamp 1710899220
transform 1 0 964 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_1016
timestamp 1710899220
transform 1 0 956 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_1017
timestamp 1710899220
transform 1 0 772 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_1018
timestamp 1710899220
transform 1 0 748 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_1019
timestamp 1710899220
transform 1 0 740 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_1020
timestamp 1710899220
transform 1 0 508 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_1021
timestamp 1710899220
transform 1 0 348 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1022
timestamp 1710899220
transform 1 0 348 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_1023
timestamp 1710899220
transform 1 0 340 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1024
timestamp 1710899220
transform 1 0 284 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1025
timestamp 1710899220
transform 1 0 276 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_1026
timestamp 1710899220
transform 1 0 276 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1027
timestamp 1710899220
transform 1 0 2004 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1028
timestamp 1710899220
transform 1 0 1988 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_1029
timestamp 1710899220
transform 1 0 1988 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_1030
timestamp 1710899220
transform 1 0 1980 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1031
timestamp 1710899220
transform 1 0 1964 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1032
timestamp 1710899220
transform 1 0 1964 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1033
timestamp 1710899220
transform 1 0 1964 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1034
timestamp 1710899220
transform 1 0 1948 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_1035
timestamp 1710899220
transform 1 0 1924 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_1036
timestamp 1710899220
transform 1 0 1924 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_1037
timestamp 1710899220
transform 1 0 1860 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1038
timestamp 1710899220
transform 1 0 1860 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1039
timestamp 1710899220
transform 1 0 1852 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1040
timestamp 1710899220
transform 1 0 1812 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1041
timestamp 1710899220
transform 1 0 1652 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1042
timestamp 1710899220
transform 1 0 1636 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_1043
timestamp 1710899220
transform 1 0 1580 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1044
timestamp 1710899220
transform 1 0 2620 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1045
timestamp 1710899220
transform 1 0 2556 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1046
timestamp 1710899220
transform 1 0 2532 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1047
timestamp 1710899220
transform 1 0 2532 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1048
timestamp 1710899220
transform 1 0 2516 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1049
timestamp 1710899220
transform 1 0 2444 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1050
timestamp 1710899220
transform 1 0 2348 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1051
timestamp 1710899220
transform 1 0 2340 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1052
timestamp 1710899220
transform 1 0 2316 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1053
timestamp 1710899220
transform 1 0 2292 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1054
timestamp 1710899220
transform 1 0 2564 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1055
timestamp 1710899220
transform 1 0 2460 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1056
timestamp 1710899220
transform 1 0 2452 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1057
timestamp 1710899220
transform 1 0 2300 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_1058
timestamp 1710899220
transform 1 0 2276 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_1059
timestamp 1710899220
transform 1 0 2268 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1060
timestamp 1710899220
transform 1 0 2252 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_1061
timestamp 1710899220
transform 1 0 2252 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1062
timestamp 1710899220
transform 1 0 2236 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1063
timestamp 1710899220
transform 1 0 2140 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1064
timestamp 1710899220
transform 1 0 2140 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1065
timestamp 1710899220
transform 1 0 2116 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1066
timestamp 1710899220
transform 1 0 1956 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1067
timestamp 1710899220
transform 1 0 1940 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1068
timestamp 1710899220
transform 1 0 1932 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1069
timestamp 1710899220
transform 1 0 1884 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1070
timestamp 1710899220
transform 1 0 1844 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1071
timestamp 1710899220
transform 1 0 1820 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1072
timestamp 1710899220
transform 1 0 2180 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1073
timestamp 1710899220
transform 1 0 2076 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_1074
timestamp 1710899220
transform 1 0 2076 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_1075
timestamp 1710899220
transform 1 0 2068 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_1076
timestamp 1710899220
transform 1 0 2036 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_1077
timestamp 1710899220
transform 1 0 2036 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1078
timestamp 1710899220
transform 1 0 2020 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1079
timestamp 1710899220
transform 1 0 2020 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_1080
timestamp 1710899220
transform 1 0 2004 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_1081
timestamp 1710899220
transform 1 0 1988 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_1082
timestamp 1710899220
transform 1 0 1964 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1083
timestamp 1710899220
transform 1 0 1940 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1084
timestamp 1710899220
transform 1 0 1932 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_1085
timestamp 1710899220
transform 1 0 1932 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1086
timestamp 1710899220
transform 1 0 1844 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1087
timestamp 1710899220
transform 1 0 1612 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_1088
timestamp 1710899220
transform 1 0 1612 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_1089
timestamp 1710899220
transform 1 0 1188 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_1090
timestamp 1710899220
transform 1 0 1180 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_1091
timestamp 1710899220
transform 1 0 1156 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1092
timestamp 1710899220
transform 1 0 1076 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_1093
timestamp 1710899220
transform 1 0 1060 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1094
timestamp 1710899220
transform 1 0 1052 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_1095
timestamp 1710899220
transform 1 0 1028 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_1096
timestamp 1710899220
transform 1 0 1004 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_1097
timestamp 1710899220
transform 1 0 996 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1098
timestamp 1710899220
transform 1 0 940 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1099
timestamp 1710899220
transform 1 0 940 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_1100
timestamp 1710899220
transform 1 0 812 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1101
timestamp 1710899220
transform 1 0 812 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1102
timestamp 1710899220
transform 1 0 716 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1103
timestamp 1710899220
transform 1 0 348 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1104
timestamp 1710899220
transform 1 0 1148 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1105
timestamp 1710899220
transform 1 0 1020 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1106
timestamp 1710899220
transform 1 0 972 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1107
timestamp 1710899220
transform 1 0 972 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1108
timestamp 1710899220
transform 1 0 924 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1109
timestamp 1710899220
transform 1 0 852 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1110
timestamp 1710899220
transform 1 0 828 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1111
timestamp 1710899220
transform 1 0 828 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1112
timestamp 1710899220
transform 1 0 796 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1113
timestamp 1710899220
transform 1 0 684 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1114
timestamp 1710899220
transform 1 0 644 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1115
timestamp 1710899220
transform 1 0 644 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1116
timestamp 1710899220
transform 1 0 596 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1117
timestamp 1710899220
transform 1 0 596 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1118
timestamp 1710899220
transform 1 0 596 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1119
timestamp 1710899220
transform 1 0 556 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1120
timestamp 1710899220
transform 1 0 492 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1121
timestamp 1710899220
transform 1 0 492 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1122
timestamp 1710899220
transform 1 0 444 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1123
timestamp 1710899220
transform 1 0 1748 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1124
timestamp 1710899220
transform 1 0 1716 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1125
timestamp 1710899220
transform 1 0 1684 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1126
timestamp 1710899220
transform 1 0 1668 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1127
timestamp 1710899220
transform 1 0 1612 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1128
timestamp 1710899220
transform 1 0 1588 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1129
timestamp 1710899220
transform 1 0 1556 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1130
timestamp 1710899220
transform 1 0 1404 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1131
timestamp 1710899220
transform 1 0 1348 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1132
timestamp 1710899220
transform 1 0 1316 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1133
timestamp 1710899220
transform 1 0 1452 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_1134
timestamp 1710899220
transform 1 0 1356 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_1135
timestamp 1710899220
transform 1 0 1348 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1136
timestamp 1710899220
transform 1 0 1252 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1137
timestamp 1710899220
transform 1 0 1220 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1138
timestamp 1710899220
transform 1 0 1220 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1139
timestamp 1710899220
transform 1 0 1188 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1140
timestamp 1710899220
transform 1 0 1180 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1141
timestamp 1710899220
transform 1 0 1156 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1142
timestamp 1710899220
transform 1 0 1148 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1143
timestamp 1710899220
transform 1 0 1124 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1144
timestamp 1710899220
transform 1 0 1116 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1145
timestamp 1710899220
transform 1 0 2012 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1146
timestamp 1710899220
transform 1 0 1948 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1147
timestamp 1710899220
transform 1 0 1876 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1148
timestamp 1710899220
transform 1 0 2228 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1149
timestamp 1710899220
transform 1 0 2044 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1150
timestamp 1710899220
transform 1 0 1932 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1151
timestamp 1710899220
transform 1 0 1916 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1152
timestamp 1710899220
transform 1 0 1644 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1153
timestamp 1710899220
transform 1 0 1860 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1154
timestamp 1710899220
transform 1 0 1732 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1155
timestamp 1710899220
transform 1 0 1612 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1156
timestamp 1710899220
transform 1 0 1612 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1157
timestamp 1710899220
transform 1 0 1524 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1158
timestamp 1710899220
transform 1 0 1380 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1159
timestamp 1710899220
transform 1 0 1340 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1160
timestamp 1710899220
transform 1 0 1332 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1161
timestamp 1710899220
transform 1 0 1316 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1162
timestamp 1710899220
transform 1 0 1044 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1163
timestamp 1710899220
transform 1 0 1004 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1164
timestamp 1710899220
transform 1 0 964 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1165
timestamp 1710899220
transform 1 0 964 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1166
timestamp 1710899220
transform 1 0 940 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1167
timestamp 1710899220
transform 1 0 940 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1168
timestamp 1710899220
transform 1 0 876 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1169
timestamp 1710899220
transform 1 0 852 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1170
timestamp 1710899220
transform 1 0 828 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1171
timestamp 1710899220
transform 1 0 676 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1172
timestamp 1710899220
transform 1 0 676 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1173
timestamp 1710899220
transform 1 0 636 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1174
timestamp 1710899220
transform 1 0 2572 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1175
timestamp 1710899220
transform 1 0 2548 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1176
timestamp 1710899220
transform 1 0 2388 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1177
timestamp 1710899220
transform 1 0 2348 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1178
timestamp 1710899220
transform 1 0 2308 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1179
timestamp 1710899220
transform 1 0 2308 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1180
timestamp 1710899220
transform 1 0 2292 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1181
timestamp 1710899220
transform 1 0 2284 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1182
timestamp 1710899220
transform 1 0 2276 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1183
timestamp 1710899220
transform 1 0 2180 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1184
timestamp 1710899220
transform 1 0 2180 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1185
timestamp 1710899220
transform 1 0 2172 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_1186
timestamp 1710899220
transform 1 0 2156 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1187
timestamp 1710899220
transform 1 0 2132 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1188
timestamp 1710899220
transform 1 0 2116 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1189
timestamp 1710899220
transform 1 0 2028 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1190
timestamp 1710899220
transform 1 0 1972 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_1191
timestamp 1710899220
transform 1 0 1956 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1192
timestamp 1710899220
transform 1 0 1940 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1193
timestamp 1710899220
transform 1 0 2652 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1194
timestamp 1710899220
transform 1 0 2604 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1195
timestamp 1710899220
transform 1 0 2564 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1196
timestamp 1710899220
transform 1 0 2564 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1197
timestamp 1710899220
transform 1 0 2532 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1198
timestamp 1710899220
transform 1 0 2532 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1199
timestamp 1710899220
transform 1 0 2524 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1200
timestamp 1710899220
transform 1 0 2484 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1201
timestamp 1710899220
transform 1 0 2484 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1202
timestamp 1710899220
transform 1 0 2484 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1203
timestamp 1710899220
transform 1 0 2364 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1204
timestamp 1710899220
transform 1 0 2364 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1205
timestamp 1710899220
transform 1 0 2332 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1206
timestamp 1710899220
transform 1 0 2292 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1207
timestamp 1710899220
transform 1 0 2188 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1208
timestamp 1710899220
transform 1 0 2052 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1209
timestamp 1710899220
transform 1 0 1964 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1210
timestamp 1710899220
transform 1 0 1452 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_1211
timestamp 1710899220
transform 1 0 1324 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1212
timestamp 1710899220
transform 1 0 1260 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1213
timestamp 1710899220
transform 1 0 1260 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1214
timestamp 1710899220
transform 1 0 1124 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1215
timestamp 1710899220
transform 1 0 1108 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1216
timestamp 1710899220
transform 1 0 1092 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1217
timestamp 1710899220
transform 1 0 2476 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1218
timestamp 1710899220
transform 1 0 2404 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1219
timestamp 1710899220
transform 1 0 2348 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1220
timestamp 1710899220
transform 1 0 2324 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1221
timestamp 1710899220
transform 1 0 2316 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1222
timestamp 1710899220
transform 1 0 2268 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1223
timestamp 1710899220
transform 1 0 2172 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1224
timestamp 1710899220
transform 1 0 2172 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1225
timestamp 1710899220
transform 1 0 2148 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1226
timestamp 1710899220
transform 1 0 2148 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1227
timestamp 1710899220
transform 1 0 1956 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_1228
timestamp 1710899220
transform 1 0 1956 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1229
timestamp 1710899220
transform 1 0 1924 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_1230
timestamp 1710899220
transform 1 0 2268 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1231
timestamp 1710899220
transform 1 0 2236 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1232
timestamp 1710899220
transform 1 0 2180 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1233
timestamp 1710899220
transform 1 0 2588 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1234
timestamp 1710899220
transform 1 0 2588 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1235
timestamp 1710899220
transform 1 0 2540 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1236
timestamp 1710899220
transform 1 0 2492 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1237
timestamp 1710899220
transform 1 0 2492 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1238
timestamp 1710899220
transform 1 0 2492 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1239
timestamp 1710899220
transform 1 0 2340 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_1240
timestamp 1710899220
transform 1 0 2284 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_1241
timestamp 1710899220
transform 1 0 2284 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1242
timestamp 1710899220
transform 1 0 2252 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1243
timestamp 1710899220
transform 1 0 2236 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1244
timestamp 1710899220
transform 1 0 2204 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1245
timestamp 1710899220
transform 1 0 2164 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1246
timestamp 1710899220
transform 1 0 2140 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1247
timestamp 1710899220
transform 1 0 220 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1248
timestamp 1710899220
transform 1 0 100 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1249
timestamp 1710899220
transform 1 0 100 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1250
timestamp 1710899220
transform 1 0 228 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_1251
timestamp 1710899220
transform 1 0 180 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_1252
timestamp 1710899220
transform 1 0 836 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1253
timestamp 1710899220
transform 1 0 804 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1254
timestamp 1710899220
transform 1 0 300 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1255
timestamp 1710899220
transform 1 0 196 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1256
timestamp 1710899220
transform 1 0 404 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1257
timestamp 1710899220
transform 1 0 308 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1258
timestamp 1710899220
transform 1 0 516 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1259
timestamp 1710899220
transform 1 0 412 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1260
timestamp 1710899220
transform 1 0 244 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1261
timestamp 1710899220
transform 1 0 156 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1262
timestamp 1710899220
transform 1 0 140 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1263
timestamp 1710899220
transform 1 0 132 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1264
timestamp 1710899220
transform 1 0 76 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1265
timestamp 1710899220
transform 1 0 1260 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1266
timestamp 1710899220
transform 1 0 1212 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1267
timestamp 1710899220
transform 1 0 196 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1268
timestamp 1710899220
transform 1 0 132 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1269
timestamp 1710899220
transform 1 0 132 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1270
timestamp 1710899220
transform 1 0 76 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1271
timestamp 1710899220
transform 1 0 148 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1272
timestamp 1710899220
transform 1 0 132 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1273
timestamp 1710899220
transform 1 0 100 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1274
timestamp 1710899220
transform 1 0 100 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1275
timestamp 1710899220
transform 1 0 164 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1276
timestamp 1710899220
transform 1 0 132 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1277
timestamp 1710899220
transform 1 0 340 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1278
timestamp 1710899220
transform 1 0 252 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1279
timestamp 1710899220
transform 1 0 252 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1280
timestamp 1710899220
transform 1 0 220 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1281
timestamp 1710899220
transform 1 0 348 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1282
timestamp 1710899220
transform 1 0 124 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1283
timestamp 1710899220
transform 1 0 492 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1284
timestamp 1710899220
transform 1 0 252 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1285
timestamp 1710899220
transform 1 0 644 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1286
timestamp 1710899220
transform 1 0 396 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1287
timestamp 1710899220
transform 1 0 964 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1288
timestamp 1710899220
transform 1 0 548 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1289
timestamp 1710899220
transform 1 0 1084 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1290
timestamp 1710899220
transform 1 0 868 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1291
timestamp 1710899220
transform 1 0 1204 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1292
timestamp 1710899220
transform 1 0 988 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1293
timestamp 1710899220
transform 1 0 1156 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1294
timestamp 1710899220
transform 1 0 1100 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1295
timestamp 1710899220
transform 1 0 244 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1296
timestamp 1710899220
transform 1 0 116 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1297
timestamp 1710899220
transform 1 0 420 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1298
timestamp 1710899220
transform 1 0 244 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1299
timestamp 1710899220
transform 1 0 420 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1300
timestamp 1710899220
transform 1 0 148 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1301
timestamp 1710899220
transform 1 0 412 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1302
timestamp 1710899220
transform 1 0 316 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1303
timestamp 1710899220
transform 1 0 636 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1304
timestamp 1710899220
transform 1 0 380 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1305
timestamp 1710899220
transform 1 0 628 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1306
timestamp 1710899220
transform 1 0 540 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1307
timestamp 1710899220
transform 1 0 652 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1308
timestamp 1710899220
transform 1 0 324 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1309
timestamp 1710899220
transform 1 0 644 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1310
timestamp 1710899220
transform 1 0 540 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1311
timestamp 1710899220
transform 1 0 452 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1312
timestamp 1710899220
transform 1 0 308 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1313
timestamp 1710899220
transform 1 0 844 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1314
timestamp 1710899220
transform 1 0 532 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1315
timestamp 1710899220
transform 1 0 892 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1316
timestamp 1710899220
transform 1 0 532 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1317
timestamp 1710899220
transform 1 0 884 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1318
timestamp 1710899220
transform 1 0 748 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1319
timestamp 1710899220
transform 1 0 772 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1320
timestamp 1710899220
transform 1 0 548 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1321
timestamp 1710899220
transform 1 0 812 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_1322
timestamp 1710899220
transform 1 0 740 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_1323
timestamp 1710899220
transform 1 0 1044 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1324
timestamp 1710899220
transform 1 0 852 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1325
timestamp 1710899220
transform 1 0 972 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1326
timestamp 1710899220
transform 1 0 724 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1327
timestamp 1710899220
transform 1 0 1084 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1328
timestamp 1710899220
transform 1 0 948 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1329
timestamp 1710899220
transform 1 0 252 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1330
timestamp 1710899220
transform 1 0 140 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1331
timestamp 1710899220
transform 1 0 452 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1332
timestamp 1710899220
transform 1 0 316 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1333
timestamp 1710899220
transform 1 0 676 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_1334
timestamp 1710899220
transform 1 0 436 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_1335
timestamp 1710899220
transform 1 0 276 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1336
timestamp 1710899220
transform 1 0 132 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1337
timestamp 1710899220
transform 1 0 428 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1338
timestamp 1710899220
transform 1 0 324 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1339
timestamp 1710899220
transform 1 0 492 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1340
timestamp 1710899220
transform 1 0 436 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1341
timestamp 1710899220
transform 1 0 476 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1342
timestamp 1710899220
transform 1 0 308 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1343
timestamp 1710899220
transform 1 0 660 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1344
timestamp 1710899220
transform 1 0 540 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1345
timestamp 1710899220
transform 1 0 884 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1346
timestamp 1710899220
transform 1 0 532 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1347
timestamp 1710899220
transform 1 0 1132 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1348
timestamp 1710899220
transform 1 0 1068 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1349
timestamp 1710899220
transform 1 0 1196 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1350
timestamp 1710899220
transform 1 0 1124 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1351
timestamp 1710899220
transform 1 0 908 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1352
timestamp 1710899220
transform 1 0 780 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1353
timestamp 1710899220
transform 1 0 1700 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1354
timestamp 1710899220
transform 1 0 1628 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1355
timestamp 1710899220
transform 1 0 1788 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1356
timestamp 1710899220
transform 1 0 1724 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1357
timestamp 1710899220
transform 1 0 1820 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1358
timestamp 1710899220
transform 1 0 1700 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1359
timestamp 1710899220
transform 1 0 1596 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1360
timestamp 1710899220
transform 1 0 1396 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1361
timestamp 1710899220
transform 1 0 1628 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1362
timestamp 1710899220
transform 1 0 1548 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1363
timestamp 1710899220
transform 1 0 1524 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1364
timestamp 1710899220
transform 1 0 1428 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1365
timestamp 1710899220
transform 1 0 820 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1366
timestamp 1710899220
transform 1 0 764 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1367
timestamp 1710899220
transform 1 0 564 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1368
timestamp 1710899220
transform 1 0 500 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1369
timestamp 1710899220
transform 1 0 220 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1370
timestamp 1710899220
transform 1 0 132 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1371
timestamp 1710899220
transform 1 0 204 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1372
timestamp 1710899220
transform 1 0 124 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1373
timestamp 1710899220
transform 1 0 428 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_1374
timestamp 1710899220
transform 1 0 276 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_1375
timestamp 1710899220
transform 1 0 732 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_1376
timestamp 1710899220
transform 1 0 580 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_1377
timestamp 1710899220
transform 1 0 1140 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1378
timestamp 1710899220
transform 1 0 1028 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1379
timestamp 1710899220
transform 1 0 1044 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_1380
timestamp 1710899220
transform 1 0 900 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_1381
timestamp 1710899220
transform 1 0 1532 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_1382
timestamp 1710899220
transform 1 0 1380 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_1383
timestamp 1710899220
transform 1 0 1692 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1384
timestamp 1710899220
transform 1 0 1628 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1385
timestamp 1710899220
transform 1 0 1708 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1386
timestamp 1710899220
transform 1 0 1668 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1387
timestamp 1710899220
transform 1 0 1788 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1388
timestamp 1710899220
transform 1 0 1716 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1389
timestamp 1710899220
transform 1 0 2236 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1390
timestamp 1710899220
transform 1 0 2220 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1391
timestamp 1710899220
transform 1 0 2084 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1392
timestamp 1710899220
transform 1 0 1588 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1393
timestamp 1710899220
transform 1 0 1516 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1394
timestamp 1710899220
transform 1 0 1436 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1395
timestamp 1710899220
transform 1 0 1524 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1396
timestamp 1710899220
transform 1 0 1460 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1397
timestamp 1710899220
transform 1 0 1420 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1398
timestamp 1710899220
transform 1 0 1348 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1399
timestamp 1710899220
transform 1 0 1436 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1400
timestamp 1710899220
transform 1 0 1404 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1401
timestamp 1710899220
transform 1 0 1356 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1402
timestamp 1710899220
transform 1 0 1332 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1403
timestamp 1710899220
transform 1 0 1252 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1404
timestamp 1710899220
transform 1 0 1220 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1405
timestamp 1710899220
transform 1 0 1140 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1406
timestamp 1710899220
transform 1 0 996 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1407
timestamp 1710899220
transform 1 0 956 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1408
timestamp 1710899220
transform 1 0 884 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1409
timestamp 1710899220
transform 1 0 700 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1410
timestamp 1710899220
transform 1 0 660 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1411
timestamp 1710899220
transform 1 0 636 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1412
timestamp 1710899220
transform 1 0 532 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1413
timestamp 1710899220
transform 1 0 364 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1414
timestamp 1710899220
transform 1 0 292 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1415
timestamp 1710899220
transform 1 0 196 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1416
timestamp 1710899220
transform 1 0 132 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1417
timestamp 1710899220
transform 1 0 180 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1418
timestamp 1710899220
transform 1 0 132 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1419
timestamp 1710899220
transform 1 0 76 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1420
timestamp 1710899220
transform 1 0 2124 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1421
timestamp 1710899220
transform 1 0 2004 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1422
timestamp 1710899220
transform 1 0 2092 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1423
timestamp 1710899220
transform 1 0 2036 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1424
timestamp 1710899220
transform 1 0 2012 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1425
timestamp 1710899220
transform 1 0 1948 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1426
timestamp 1710899220
transform 1 0 2052 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1427
timestamp 1710899220
transform 1 0 1988 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1428
timestamp 1710899220
transform 1 0 212 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1429
timestamp 1710899220
transform 1 0 148 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1430
timestamp 1710899220
transform 1 0 252 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1431
timestamp 1710899220
transform 1 0 188 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1432
timestamp 1710899220
transform 1 0 364 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1433
timestamp 1710899220
transform 1 0 284 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1434
timestamp 1710899220
transform 1 0 460 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1435
timestamp 1710899220
transform 1 0 396 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1436
timestamp 1710899220
transform 1 0 636 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1437
timestamp 1710899220
transform 1 0 532 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1438
timestamp 1710899220
transform 1 0 964 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1439
timestamp 1710899220
transform 1 0 788 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1440
timestamp 1710899220
transform 1 0 1084 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1441
timestamp 1710899220
transform 1 0 996 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1442
timestamp 1710899220
transform 1 0 1188 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1443
timestamp 1710899220
transform 1 0 1148 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1444
timestamp 1710899220
transform 1 0 1372 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1445
timestamp 1710899220
transform 1 0 1292 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1446
timestamp 1710899220
transform 1 0 2308 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1447
timestamp 1710899220
transform 1 0 2204 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1448
timestamp 1710899220
transform 1 0 2156 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1449
timestamp 1710899220
transform 1 0 2068 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1450
timestamp 1710899220
transform 1 0 1996 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1451
timestamp 1710899220
transform 1 0 1996 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1452
timestamp 1710899220
transform 1 0 1964 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1453
timestamp 1710899220
transform 1 0 1964 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1454
timestamp 1710899220
transform 1 0 1884 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1455
timestamp 1710899220
transform 1 0 1764 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1456
timestamp 1710899220
transform 1 0 1596 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1457
timestamp 1710899220
transform 1 0 1548 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1458
timestamp 1710899220
transform 1 0 1532 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1459
timestamp 1710899220
transform 1 0 1532 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1460
timestamp 1710899220
transform 1 0 1508 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1461
timestamp 1710899220
transform 1 0 1500 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1462
timestamp 1710899220
transform 1 0 1428 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1463
timestamp 1710899220
transform 1 0 1428 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1464
timestamp 1710899220
transform 1 0 1420 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1465
timestamp 1710899220
transform 1 0 1340 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1466
timestamp 1710899220
transform 1 0 1268 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1467
timestamp 1710899220
transform 1 0 1188 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1468
timestamp 1710899220
transform 1 0 1188 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1469
timestamp 1710899220
transform 1 0 1140 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1470
timestamp 1710899220
transform 1 0 972 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1471
timestamp 1710899220
transform 1 0 940 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1472
timestamp 1710899220
transform 1 0 828 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1473
timestamp 1710899220
transform 1 0 828 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1474
timestamp 1710899220
transform 1 0 1356 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1475
timestamp 1710899220
transform 1 0 1036 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1476
timestamp 1710899220
transform 1 0 1388 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1477
timestamp 1710899220
transform 1 0 1340 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1478
timestamp 1710899220
transform 1 0 2004 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1479
timestamp 1710899220
transform 1 0 1676 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1480
timestamp 1710899220
transform 1 0 1580 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1481
timestamp 1710899220
transform 1 0 1444 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1482
timestamp 1710899220
transform 1 0 1548 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1483
timestamp 1710899220
transform 1 0 1380 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1484
timestamp 1710899220
transform 1 0 1236 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1485
timestamp 1710899220
transform 1 0 684 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1486
timestamp 1710899220
transform 1 0 668 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1487
timestamp 1710899220
transform 1 0 1084 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1488
timestamp 1710899220
transform 1 0 708 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1489
timestamp 1710899220
transform 1 0 1284 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1490
timestamp 1710899220
transform 1 0 1164 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1491
timestamp 1710899220
transform 1 0 1076 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1492
timestamp 1710899220
transform 1 0 1700 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1493
timestamp 1710899220
transform 1 0 1668 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1494
timestamp 1710899220
transform 1 0 1660 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_1495
timestamp 1710899220
transform 1 0 1196 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_1496
timestamp 1710899220
transform 1 0 1108 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1497
timestamp 1710899220
transform 1 0 1108 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_1498
timestamp 1710899220
transform 1 0 1060 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1499
timestamp 1710899220
transform 1 0 956 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1500
timestamp 1710899220
transform 1 0 932 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1501
timestamp 1710899220
transform 1 0 1148 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1502
timestamp 1710899220
transform 1 0 1076 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1503
timestamp 1710899220
transform 1 0 1308 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1504
timestamp 1710899220
transform 1 0 1156 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1505
timestamp 1710899220
transform 1 0 1124 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1506
timestamp 1710899220
transform 1 0 660 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1507
timestamp 1710899220
transform 1 0 1564 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1508
timestamp 1710899220
transform 1 0 1532 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1509
timestamp 1710899220
transform 1 0 1260 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1510
timestamp 1710899220
transform 1 0 1204 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1511
timestamp 1710899220
transform 1 0 1188 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1512
timestamp 1710899220
transform 1 0 1188 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1513
timestamp 1710899220
transform 1 0 1164 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1514
timestamp 1710899220
transform 1 0 1140 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1515
timestamp 1710899220
transform 1 0 1108 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1516
timestamp 1710899220
transform 1 0 1188 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1517
timestamp 1710899220
transform 1 0 1036 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1518
timestamp 1710899220
transform 1 0 1724 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1519
timestamp 1710899220
transform 1 0 1684 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1520
timestamp 1710899220
transform 1 0 1636 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1521
timestamp 1710899220
transform 1 0 1332 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1522
timestamp 1710899220
transform 1 0 1300 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1523
timestamp 1710899220
transform 1 0 1164 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1524
timestamp 1710899220
transform 1 0 1404 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1525
timestamp 1710899220
transform 1 0 1300 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1526
timestamp 1710899220
transform 1 0 1180 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1527
timestamp 1710899220
transform 1 0 1060 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1528
timestamp 1710899220
transform 1 0 1588 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1529
timestamp 1710899220
transform 1 0 1252 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1530
timestamp 1710899220
transform 1 0 1252 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1531
timestamp 1710899220
transform 1 0 1180 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1532
timestamp 1710899220
transform 1 0 836 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1533
timestamp 1710899220
transform 1 0 820 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1534
timestamp 1710899220
transform 1 0 1260 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1535
timestamp 1710899220
transform 1 0 916 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1536
timestamp 1710899220
transform 1 0 916 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1537
timestamp 1710899220
transform 1 0 852 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1538
timestamp 1710899220
transform 1 0 1252 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1539
timestamp 1710899220
transform 1 0 1180 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1540
timestamp 1710899220
transform 1 0 1220 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1541
timestamp 1710899220
transform 1 0 1164 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1542
timestamp 1710899220
transform 1 0 1324 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1543
timestamp 1710899220
transform 1 0 1204 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1544
timestamp 1710899220
transform 1 0 1412 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1545
timestamp 1710899220
transform 1 0 1340 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1546
timestamp 1710899220
transform 1 0 1276 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1547
timestamp 1710899220
transform 1 0 1100 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1548
timestamp 1710899220
transform 1 0 1788 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1549
timestamp 1710899220
transform 1 0 1684 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1550
timestamp 1710899220
transform 1 0 1652 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1551
timestamp 1710899220
transform 1 0 1508 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1552
timestamp 1710899220
transform 1 0 1692 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1553
timestamp 1710899220
transform 1 0 1548 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1554
timestamp 1710899220
transform 1 0 1628 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1555
timestamp 1710899220
transform 1 0 1572 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1556
timestamp 1710899220
transform 1 0 1540 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1557
timestamp 1710899220
transform 1 0 1516 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1558
timestamp 1710899220
transform 1 0 1604 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1559
timestamp 1710899220
transform 1 0 1572 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1560
timestamp 1710899220
transform 1 0 1668 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1561
timestamp 1710899220
transform 1 0 1628 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1562
timestamp 1710899220
transform 1 0 1860 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1563
timestamp 1710899220
transform 1 0 1820 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1564
timestamp 1710899220
transform 1 0 1676 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1565
timestamp 1710899220
transform 1 0 1620 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1566
timestamp 1710899220
transform 1 0 1716 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1567
timestamp 1710899220
transform 1 0 1580 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1568
timestamp 1710899220
transform 1 0 2148 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_1569
timestamp 1710899220
transform 1 0 2108 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_1570
timestamp 1710899220
transform 1 0 2028 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_1571
timestamp 1710899220
transform 1 0 1380 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1572
timestamp 1710899220
transform 1 0 1340 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1573
timestamp 1710899220
transform 1 0 1900 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1574
timestamp 1710899220
transform 1 0 1604 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1575
timestamp 1710899220
transform 1 0 1532 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1576
timestamp 1710899220
transform 1 0 1420 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1577
timestamp 1710899220
transform 1 0 1332 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1578
timestamp 1710899220
transform 1 0 2236 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1579
timestamp 1710899220
transform 1 0 2180 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1580
timestamp 1710899220
transform 1 0 2148 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1581
timestamp 1710899220
transform 1 0 2036 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1582
timestamp 1710899220
transform 1 0 2244 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1583
timestamp 1710899220
transform 1 0 2156 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1584
timestamp 1710899220
transform 1 0 2292 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1585
timestamp 1710899220
transform 1 0 2268 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1586
timestamp 1710899220
transform 1 0 2244 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1587
timestamp 1710899220
transform 1 0 2220 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1588
timestamp 1710899220
transform 1 0 972 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1589
timestamp 1710899220
transform 1 0 892 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1590
timestamp 1710899220
transform 1 0 692 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1591
timestamp 1710899220
transform 1 0 588 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1592
timestamp 1710899220
transform 1 0 964 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1593
timestamp 1710899220
transform 1 0 868 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1594
timestamp 1710899220
transform 1 0 652 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1595
timestamp 1710899220
transform 1 0 524 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1596
timestamp 1710899220
transform 1 0 1052 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1597
timestamp 1710899220
transform 1 0 996 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1598
timestamp 1710899220
transform 1 0 1004 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1599
timestamp 1710899220
transform 1 0 932 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1600
timestamp 1710899220
transform 1 0 1028 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1601
timestamp 1710899220
transform 1 0 972 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1602
timestamp 1710899220
transform 1 0 884 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1603
timestamp 1710899220
transform 1 0 828 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1604
timestamp 1710899220
transform 1 0 844 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1605
timestamp 1710899220
transform 1 0 748 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1606
timestamp 1710899220
transform 1 0 1180 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1607
timestamp 1710899220
transform 1 0 1084 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1608
timestamp 1710899220
transform 1 0 1124 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1609
timestamp 1710899220
transform 1 0 1044 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1610
timestamp 1710899220
transform 1 0 1284 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1611
timestamp 1710899220
transform 1 0 1196 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1612
timestamp 1710899220
transform 1 0 1156 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1613
timestamp 1710899220
transform 1 0 1084 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1614
timestamp 1710899220
transform 1 0 1348 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1615
timestamp 1710899220
transform 1 0 1276 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1616
timestamp 1710899220
transform 1 0 1420 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1617
timestamp 1710899220
transform 1 0 1356 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1618
timestamp 1710899220
transform 1 0 868 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1619
timestamp 1710899220
transform 1 0 804 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1620
timestamp 1710899220
transform 1 0 1468 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1621
timestamp 1710899220
transform 1 0 1396 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1622
timestamp 1710899220
transform 1 0 1540 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1623
timestamp 1710899220
transform 1 0 1468 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1624
timestamp 1710899220
transform 1 0 1908 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1625
timestamp 1710899220
transform 1 0 1868 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1626
timestamp 1710899220
transform 1 0 1796 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1627
timestamp 1710899220
transform 1 0 1756 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1628
timestamp 1710899220
transform 1 0 1828 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1629
timestamp 1710899220
transform 1 0 1788 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1630
timestamp 1710899220
transform 1 0 1372 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1631
timestamp 1710899220
transform 1 0 1252 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1632
timestamp 1710899220
transform 1 0 1372 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1633
timestamp 1710899220
transform 1 0 1284 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1634
timestamp 1710899220
transform 1 0 1372 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1635
timestamp 1710899220
transform 1 0 1356 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1636
timestamp 1710899220
transform 1 0 1348 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1637
timestamp 1710899220
transform 1 0 1284 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1638
timestamp 1710899220
transform 1 0 1428 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1639
timestamp 1710899220
transform 1 0 1340 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1640
timestamp 1710899220
transform 1 0 1444 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_1641
timestamp 1710899220
transform 1 0 1324 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_1642
timestamp 1710899220
transform 1 0 1380 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1643
timestamp 1710899220
transform 1 0 1356 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1644
timestamp 1710899220
transform 1 0 1428 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1645
timestamp 1710899220
transform 1 0 1372 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1646
timestamp 1710899220
transform 1 0 1404 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1647
timestamp 1710899220
transform 1 0 1340 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1648
timestamp 1710899220
transform 1 0 708 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1649
timestamp 1710899220
transform 1 0 644 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1650
timestamp 1710899220
transform 1 0 724 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1651
timestamp 1710899220
transform 1 0 684 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1652
timestamp 1710899220
transform 1 0 780 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1653
timestamp 1710899220
transform 1 0 660 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1654
timestamp 1710899220
transform 1 0 748 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1655
timestamp 1710899220
transform 1 0 716 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1656
timestamp 1710899220
transform 1 0 532 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1657
timestamp 1710899220
transform 1 0 396 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1658
timestamp 1710899220
transform 1 0 396 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_1659
timestamp 1710899220
transform 1 0 260 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_1660
timestamp 1710899220
transform 1 0 172 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_1661
timestamp 1710899220
transform 1 0 284 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_1662
timestamp 1710899220
transform 1 0 228 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1663
timestamp 1710899220
transform 1 0 212 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1664
timestamp 1710899220
transform 1 0 164 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1665
timestamp 1710899220
transform 1 0 124 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1666
timestamp 1710899220
transform 1 0 404 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1667
timestamp 1710899220
transform 1 0 340 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1668
timestamp 1710899220
transform 1 0 324 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1669
timestamp 1710899220
transform 1 0 308 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_1670
timestamp 1710899220
transform 1 0 308 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1671
timestamp 1710899220
transform 1 0 300 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1672
timestamp 1710899220
transform 1 0 236 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_1673
timestamp 1710899220
transform 1 0 188 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_1674
timestamp 1710899220
transform 1 0 284 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1675
timestamp 1710899220
transform 1 0 260 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1676
timestamp 1710899220
transform 1 0 204 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1677
timestamp 1710899220
transform 1 0 756 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1678
timestamp 1710899220
transform 1 0 716 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1679
timestamp 1710899220
transform 1 0 652 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1680
timestamp 1710899220
transform 1 0 644 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1681
timestamp 1710899220
transform 1 0 628 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1682
timestamp 1710899220
transform 1 0 620 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1683
timestamp 1710899220
transform 1 0 820 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1684
timestamp 1710899220
transform 1 0 716 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1685
timestamp 1710899220
transform 1 0 1460 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1686
timestamp 1710899220
transform 1 0 1460 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1687
timestamp 1710899220
transform 1 0 1404 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1688
timestamp 1710899220
transform 1 0 1300 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1689
timestamp 1710899220
transform 1 0 1116 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1690
timestamp 1710899220
transform 1 0 1580 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1691
timestamp 1710899220
transform 1 0 1428 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1692
timestamp 1710899220
transform 1 0 1412 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1693
timestamp 1710899220
transform 1 0 1156 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1694
timestamp 1710899220
transform 1 0 1652 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1695
timestamp 1710899220
transform 1 0 1444 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1696
timestamp 1710899220
transform 1 0 1420 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1697
timestamp 1710899220
transform 1 0 1076 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1698
timestamp 1710899220
transform 1 0 1548 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_1699
timestamp 1710899220
transform 1 0 1516 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_1700
timestamp 1710899220
transform 1 0 1604 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1701
timestamp 1710899220
transform 1 0 1484 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1702
timestamp 1710899220
transform 1 0 2340 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_1703
timestamp 1710899220
transform 1 0 2276 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_1704
timestamp 1710899220
transform 1 0 2236 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1705
timestamp 1710899220
transform 1 0 2148 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1706
timestamp 1710899220
transform 1 0 2236 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1707
timestamp 1710899220
transform 1 0 2164 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1708
timestamp 1710899220
transform 1 0 2036 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1709
timestamp 1710899220
transform 1 0 1932 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1710
timestamp 1710899220
transform 1 0 2004 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1711
timestamp 1710899220
transform 1 0 1900 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1712
timestamp 1710899220
transform 1 0 2036 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1713
timestamp 1710899220
transform 1 0 1940 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1714
timestamp 1710899220
transform 1 0 2036 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1715
timestamp 1710899220
transform 1 0 1932 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1716
timestamp 1710899220
transform 1 0 2052 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1717
timestamp 1710899220
transform 1 0 1948 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1718
timestamp 1710899220
transform 1 0 2124 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1719
timestamp 1710899220
transform 1 0 2004 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1720
timestamp 1710899220
transform 1 0 2460 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1721
timestamp 1710899220
transform 1 0 2364 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1722
timestamp 1710899220
transform 1 0 2428 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1723
timestamp 1710899220
transform 1 0 2332 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1724
timestamp 1710899220
transform 1 0 2444 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1725
timestamp 1710899220
transform 1 0 2348 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1726
timestamp 1710899220
transform 1 0 2444 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1727
timestamp 1710899220
transform 1 0 2348 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1728
timestamp 1710899220
transform 1 0 2412 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1729
timestamp 1710899220
transform 1 0 2292 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1730
timestamp 1710899220
transform 1 0 2436 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1731
timestamp 1710899220
transform 1 0 2324 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1732
timestamp 1710899220
transform 1 0 2564 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_1733
timestamp 1710899220
transform 1 0 2508 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_1734
timestamp 1710899220
transform 1 0 2644 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1735
timestamp 1710899220
transform 1 0 2580 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1736
timestamp 1710899220
transform 1 0 1460 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_1737
timestamp 1710899220
transform 1 0 1276 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_1738
timestamp 1710899220
transform 1 0 1452 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1739
timestamp 1710899220
transform 1 0 1364 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1740
timestamp 1710899220
transform 1 0 1780 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1741
timestamp 1710899220
transform 1 0 1284 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1742
timestamp 1710899220
transform 1 0 1556 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_1743
timestamp 1710899220
transform 1 0 1492 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_1744
timestamp 1710899220
transform 1 0 1628 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1745
timestamp 1710899220
transform 1 0 1556 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1746
timestamp 1710899220
transform 1 0 1532 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1747
timestamp 1710899220
transform 1 0 1372 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1748
timestamp 1710899220
transform 1 0 1612 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1749
timestamp 1710899220
transform 1 0 1556 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1750
timestamp 1710899220
transform 1 0 1476 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1751
timestamp 1710899220
transform 1 0 1452 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1752
timestamp 1710899220
transform 1 0 1284 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1753
timestamp 1710899220
transform 1 0 1452 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_1754
timestamp 1710899220
transform 1 0 1364 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_1755
timestamp 1710899220
transform 1 0 2156 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1756
timestamp 1710899220
transform 1 0 2084 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1757
timestamp 1710899220
transform 1 0 2084 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1758
timestamp 1710899220
transform 1 0 2012 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1759
timestamp 1710899220
transform 1 0 2012 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_1760
timestamp 1710899220
transform 1 0 1996 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_1761
timestamp 1710899220
transform 1 0 1988 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1762
timestamp 1710899220
transform 1 0 1884 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_1763
timestamp 1710899220
transform 1 0 1772 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_1764
timestamp 1710899220
transform 1 0 1772 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1765
timestamp 1710899220
transform 1 0 1692 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_1766
timestamp 1710899220
transform 1 0 1692 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_1767
timestamp 1710899220
transform 1 0 1660 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1768
timestamp 1710899220
transform 1 0 1124 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_1769
timestamp 1710899220
transform 1 0 540 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_1770
timestamp 1710899220
transform 1 0 532 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_1771
timestamp 1710899220
transform 1 0 388 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_1772
timestamp 1710899220
transform 1 0 2252 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1773
timestamp 1710899220
transform 1 0 2196 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1774
timestamp 1710899220
transform 1 0 2292 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1775
timestamp 1710899220
transform 1 0 2164 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1776
timestamp 1710899220
transform 1 0 2212 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1777
timestamp 1710899220
transform 1 0 2132 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1778
timestamp 1710899220
transform 1 0 2108 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1779
timestamp 1710899220
transform 1 0 2268 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1780
timestamp 1710899220
transform 1 0 2220 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1781
timestamp 1710899220
transform 1 0 2012 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_1782
timestamp 1710899220
transform 1 0 1876 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_1783
timestamp 1710899220
transform 1 0 1820 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_1784
timestamp 1710899220
transform 1 0 1980 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1785
timestamp 1710899220
transform 1 0 1972 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1786
timestamp 1710899220
transform 1 0 1940 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1787
timestamp 1710899220
transform 1 0 1940 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1788
timestamp 1710899220
transform 1 0 1772 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1789
timestamp 1710899220
transform 1 0 1708 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1790
timestamp 1710899220
transform 1 0 1708 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1791
timestamp 1710899220
transform 1 0 1700 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1792
timestamp 1710899220
transform 1 0 1732 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1793
timestamp 1710899220
transform 1 0 1692 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1794
timestamp 1710899220
transform 1 0 1692 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_1795
timestamp 1710899220
transform 1 0 1524 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_1796
timestamp 1710899220
transform 1 0 1716 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1797
timestamp 1710899220
transform 1 0 1580 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1798
timestamp 1710899220
transform 1 0 1980 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1799
timestamp 1710899220
transform 1 0 1972 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1800
timestamp 1710899220
transform 1 0 1804 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1801
timestamp 1710899220
transform 1 0 1716 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_1802
timestamp 1710899220
transform 1 0 1732 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1803
timestamp 1710899220
transform 1 0 1540 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1804
timestamp 1710899220
transform 1 0 1548 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1805
timestamp 1710899220
transform 1 0 1540 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1806
timestamp 1710899220
transform 1 0 1492 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1807
timestamp 1710899220
transform 1 0 1484 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1808
timestamp 1710899220
transform 1 0 1516 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1809
timestamp 1710899220
transform 1 0 1428 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1810
timestamp 1710899220
transform 1 0 1404 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1811
timestamp 1710899220
transform 1 0 1284 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1812
timestamp 1710899220
transform 1 0 1524 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1813
timestamp 1710899220
transform 1 0 1484 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1814
timestamp 1710899220
transform 1 0 1500 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1815
timestamp 1710899220
transform 1 0 1468 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1816
timestamp 1710899220
transform 1 0 1404 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1817
timestamp 1710899220
transform 1 0 1372 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1818
timestamp 1710899220
transform 1 0 1492 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1819
timestamp 1710899220
transform 1 0 1444 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1820
timestamp 1710899220
transform 1 0 1532 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_1821
timestamp 1710899220
transform 1 0 1484 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_1822
timestamp 1710899220
transform 1 0 1508 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1823
timestamp 1710899220
transform 1 0 1396 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1824
timestamp 1710899220
transform 1 0 1412 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1825
timestamp 1710899220
transform 1 0 1388 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1826
timestamp 1710899220
transform 1 0 1204 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1827
timestamp 1710899220
transform 1 0 1204 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1828
timestamp 1710899220
transform 1 0 1060 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1829
timestamp 1710899220
transform 1 0 1788 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1830
timestamp 1710899220
transform 1 0 1740 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1831
timestamp 1710899220
transform 1 0 1268 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1832
timestamp 1710899220
transform 1 0 1244 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1833
timestamp 1710899220
transform 1 0 1268 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_1834
timestamp 1710899220
transform 1 0 1236 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_1835
timestamp 1710899220
transform 1 0 1812 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1836
timestamp 1710899220
transform 1 0 1228 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_1837
timestamp 1710899220
transform 1 0 1252 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_1838
timestamp 1710899220
transform 1 0 580 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_1839
timestamp 1710899220
transform 1 0 1244 0 1 75
box -3 -3 3 3
use M3_M2  M3_M2_1840
timestamp 1710899220
transform 1 0 892 0 1 75
box -3 -3 3 3
use M3_M2  M3_M2_1841
timestamp 1710899220
transform 1 0 2660 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1842
timestamp 1710899220
transform 1 0 2596 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_1843
timestamp 1710899220
transform 1 0 2524 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1844
timestamp 1710899220
transform 1 0 2508 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1845
timestamp 1710899220
transform 1 0 2668 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1846
timestamp 1710899220
transform 1 0 2556 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1847
timestamp 1710899220
transform 1 0 2548 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1848
timestamp 1710899220
transform 1 0 2524 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1849
timestamp 1710899220
transform 1 0 2556 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1850
timestamp 1710899220
transform 1 0 2540 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1851
timestamp 1710899220
transform 1 0 2652 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1852
timestamp 1710899220
transform 1 0 2540 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1853
timestamp 1710899220
transform 1 0 2316 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_1854
timestamp 1710899220
transform 1 0 2300 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_1855
timestamp 1710899220
transform 1 0 1948 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1856
timestamp 1710899220
transform 1 0 1916 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1857
timestamp 1710899220
transform 1 0 1948 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1858
timestamp 1710899220
transform 1 0 1924 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1859
timestamp 1710899220
transform 1 0 2284 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1860
timestamp 1710899220
transform 1 0 2252 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1861
timestamp 1710899220
transform 1 0 2060 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1862
timestamp 1710899220
transform 1 0 2036 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1863
timestamp 1710899220
transform 1 0 1964 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1864
timestamp 1710899220
transform 1 0 1948 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1865
timestamp 1710899220
transform 1 0 1892 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_1866
timestamp 1710899220
transform 1 0 1892 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1867
timestamp 1710899220
transform 1 0 1756 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1868
timestamp 1710899220
transform 1 0 1756 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1869
timestamp 1710899220
transform 1 0 1724 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1870
timestamp 1710899220
transform 1 0 1708 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1871
timestamp 1710899220
transform 1 0 1636 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1872
timestamp 1710899220
transform 1 0 1724 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1873
timestamp 1710899220
transform 1 0 1700 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1874
timestamp 1710899220
transform 1 0 1636 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_1875
timestamp 1710899220
transform 1 0 1500 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_1876
timestamp 1710899220
transform 1 0 1700 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1877
timestamp 1710899220
transform 1 0 1532 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_1878
timestamp 1710899220
transform 1 0 1532 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1879
timestamp 1710899220
transform 1 0 596 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1880
timestamp 1710899220
transform 1 0 1812 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1881
timestamp 1710899220
transform 1 0 1652 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1882
timestamp 1710899220
transform 1 0 1612 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1883
timestamp 1710899220
transform 1 0 1804 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_1884
timestamp 1710899220
transform 1 0 1612 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_1885
timestamp 1710899220
transform 1 0 1460 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_1886
timestamp 1710899220
transform 1 0 1460 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_1887
timestamp 1710899220
transform 1 0 1068 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_1888
timestamp 1710899220
transform 1 0 1620 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1889
timestamp 1710899220
transform 1 0 1620 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1890
timestamp 1710899220
transform 1 0 1572 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1891
timestamp 1710899220
transform 1 0 1436 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1892
timestamp 1710899220
transform 1 0 1436 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_1893
timestamp 1710899220
transform 1 0 764 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_1894
timestamp 1710899220
transform 1 0 1604 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_1895
timestamp 1710899220
transform 1 0 1044 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1896
timestamp 1710899220
transform 1 0 1660 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1897
timestamp 1710899220
transform 1 0 1076 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1898
timestamp 1710899220
transform 1 0 1668 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1899
timestamp 1710899220
transform 1 0 1556 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1900
timestamp 1710899220
transform 1 0 1556 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1901
timestamp 1710899220
transform 1 0 1348 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1902
timestamp 1710899220
transform 1 0 1348 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1903
timestamp 1710899220
transform 1 0 844 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_1904
timestamp 1710899220
transform 1 0 1876 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_1905
timestamp 1710899220
transform 1 0 1876 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_1906
timestamp 1710899220
transform 1 0 1788 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_1907
timestamp 1710899220
transform 1 0 1700 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_1908
timestamp 1710899220
transform 1 0 1908 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_1909
timestamp 1710899220
transform 1 0 1780 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_1910
timestamp 1710899220
transform 1 0 1740 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1911
timestamp 1710899220
transform 1 0 1668 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1912
timestamp 1710899220
transform 1 0 604 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_1913
timestamp 1710899220
transform 1 0 452 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_1914
timestamp 1710899220
transform 1 0 1036 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1915
timestamp 1710899220
transform 1 0 884 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1916
timestamp 1710899220
transform 1 0 772 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1917
timestamp 1710899220
transform 1 0 724 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1918
timestamp 1710899220
transform 1 0 1804 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1919
timestamp 1710899220
transform 1 0 1780 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1920
timestamp 1710899220
transform 1 0 1668 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1921
timestamp 1710899220
transform 1 0 1580 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1922
timestamp 1710899220
transform 1 0 1924 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1923
timestamp 1710899220
transform 1 0 1908 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1924
timestamp 1710899220
transform 1 0 1996 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_1925
timestamp 1710899220
transform 1 0 1932 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_1926
timestamp 1710899220
transform 1 0 2028 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1927
timestamp 1710899220
transform 1 0 1964 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1928
timestamp 1710899220
transform 1 0 1900 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_1929
timestamp 1710899220
transform 1 0 1828 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_1930
timestamp 1710899220
transform 1 0 1076 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1931
timestamp 1710899220
transform 1 0 1044 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1932
timestamp 1710899220
transform 1 0 1868 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1933
timestamp 1710899220
transform 1 0 1724 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1934
timestamp 1710899220
transform 1 0 1740 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_1935
timestamp 1710899220
transform 1 0 1644 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_1936
timestamp 1710899220
transform 1 0 1644 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1937
timestamp 1710899220
transform 1 0 1572 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1938
timestamp 1710899220
transform 1 0 1708 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1939
timestamp 1710899220
transform 1 0 1652 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1940
timestamp 1710899220
transform 1 0 1684 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_1941
timestamp 1710899220
transform 1 0 1588 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_1942
timestamp 1710899220
transform 1 0 1764 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1943
timestamp 1710899220
transform 1 0 1716 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1944
timestamp 1710899220
transform 1 0 1876 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1945
timestamp 1710899220
transform 1 0 1708 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1946
timestamp 1710899220
transform 1 0 1932 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1947
timestamp 1710899220
transform 1 0 1892 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1948
timestamp 1710899220
transform 1 0 836 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_1949
timestamp 1710899220
transform 1 0 524 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_1950
timestamp 1710899220
transform 1 0 900 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1951
timestamp 1710899220
transform 1 0 860 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1952
timestamp 1710899220
transform 1 0 932 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1953
timestamp 1710899220
transform 1 0 868 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1954
timestamp 1710899220
transform 1 0 876 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1955
timestamp 1710899220
transform 1 0 652 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1956
timestamp 1710899220
transform 1 0 636 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1957
timestamp 1710899220
transform 1 0 540 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1958
timestamp 1710899220
transform 1 0 540 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1959
timestamp 1710899220
transform 1 0 396 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_1960
timestamp 1710899220
transform 1 0 1004 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1961
timestamp 1710899220
transform 1 0 508 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_1962
timestamp 1710899220
transform 1 0 500 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1963
timestamp 1710899220
transform 1 0 452 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1964
timestamp 1710899220
transform 1 0 460 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_1965
timestamp 1710899220
transform 1 0 444 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_1966
timestamp 1710899220
transform 1 0 572 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_1967
timestamp 1710899220
transform 1 0 452 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1968
timestamp 1710899220
transform 1 0 1028 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1969
timestamp 1710899220
transform 1 0 988 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1970
timestamp 1710899220
transform 1 0 1052 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1971
timestamp 1710899220
transform 1 0 1020 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1972
timestamp 1710899220
transform 1 0 1060 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1973
timestamp 1710899220
transform 1 0 636 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1974
timestamp 1710899220
transform 1 0 1044 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1975
timestamp 1710899220
transform 1 0 948 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1976
timestamp 1710899220
transform 1 0 1036 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1977
timestamp 1710899220
transform 1 0 988 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1978
timestamp 1710899220
transform 1 0 1620 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_1979
timestamp 1710899220
transform 1 0 1364 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1980
timestamp 1710899220
transform 1 0 1364 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1981
timestamp 1710899220
transform 1 0 1044 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1982
timestamp 1710899220
transform 1 0 1692 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_1983
timestamp 1710899220
transform 1 0 1652 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_1984
timestamp 1710899220
transform 1 0 1788 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1985
timestamp 1710899220
transform 1 0 1692 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1986
timestamp 1710899220
transform 1 0 1100 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_1987
timestamp 1710899220
transform 1 0 972 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_1988
timestamp 1710899220
transform 1 0 612 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1989
timestamp 1710899220
transform 1 0 412 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1990
timestamp 1710899220
transform 1 0 620 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1991
timestamp 1710899220
transform 1 0 540 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1992
timestamp 1710899220
transform 1 0 804 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1993
timestamp 1710899220
transform 1 0 628 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1994
timestamp 1710899220
transform 1 0 932 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1995
timestamp 1710899220
transform 1 0 772 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1996
timestamp 1710899220
transform 1 0 804 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1997
timestamp 1710899220
transform 1 0 780 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1998
timestamp 1710899220
transform 1 0 652 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1999
timestamp 1710899220
transform 1 0 596 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2000
timestamp 1710899220
transform 1 0 596 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2001
timestamp 1710899220
transform 1 0 524 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2002
timestamp 1710899220
transform 1 0 1860 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2003
timestamp 1710899220
transform 1 0 1844 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2004
timestamp 1710899220
transform 1 0 1836 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2005
timestamp 1710899220
transform 1 0 1316 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_2006
timestamp 1710899220
transform 1 0 1316 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2007
timestamp 1710899220
transform 1 0 1028 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2008
timestamp 1710899220
transform 1 0 1028 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2009
timestamp 1710899220
transform 1 0 724 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2010
timestamp 1710899220
transform 1 0 724 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2011
timestamp 1710899220
transform 1 0 684 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2012
timestamp 1710899220
transform 1 0 1732 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2013
timestamp 1710899220
transform 1 0 1524 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2014
timestamp 1710899220
transform 1 0 1524 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2015
timestamp 1710899220
transform 1 0 1436 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2016
timestamp 1710899220
transform 1 0 1276 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2017
timestamp 1710899220
transform 1 0 1452 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_2018
timestamp 1710899220
transform 1 0 1332 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_2019
timestamp 1710899220
transform 1 0 1324 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_2020
timestamp 1710899220
transform 1 0 1300 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_2021
timestamp 1710899220
transform 1 0 1300 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2022
timestamp 1710899220
transform 1 0 1252 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2023
timestamp 1710899220
transform 1 0 1820 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_2024
timestamp 1710899220
transform 1 0 1404 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_2025
timestamp 1710899220
transform 1 0 1780 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2026
timestamp 1710899220
transform 1 0 1444 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2027
timestamp 1710899220
transform 1 0 1548 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2028
timestamp 1710899220
transform 1 0 1404 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2029
timestamp 1710899220
transform 1 0 1420 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_2030
timestamp 1710899220
transform 1 0 1364 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_2031
timestamp 1710899220
transform 1 0 1420 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2032
timestamp 1710899220
transform 1 0 1380 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2033
timestamp 1710899220
transform 1 0 1772 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_2034
timestamp 1710899220
transform 1 0 1420 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2035
timestamp 1710899220
transform 1 0 1828 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_2036
timestamp 1710899220
transform 1 0 1436 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_2037
timestamp 1710899220
transform 1 0 1788 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_2038
timestamp 1710899220
transform 1 0 1484 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_2039
timestamp 1710899220
transform 1 0 1508 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2040
timestamp 1710899220
transform 1 0 1468 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2041
timestamp 1710899220
transform 1 0 1452 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2042
timestamp 1710899220
transform 1 0 1420 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2043
timestamp 1710899220
transform 1 0 1332 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2044
timestamp 1710899220
transform 1 0 1292 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2045
timestamp 1710899220
transform 1 0 908 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2046
timestamp 1710899220
transform 1 0 820 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2047
timestamp 1710899220
transform 1 0 828 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_2048
timestamp 1710899220
transform 1 0 764 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_2049
timestamp 1710899220
transform 1 0 684 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2050
timestamp 1710899220
transform 1 0 564 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2051
timestamp 1710899220
transform 1 0 628 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2052
timestamp 1710899220
transform 1 0 540 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2053
timestamp 1710899220
transform 1 0 708 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2054
timestamp 1710899220
transform 1 0 660 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2055
timestamp 1710899220
transform 1 0 2116 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2056
timestamp 1710899220
transform 1 0 1740 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2057
timestamp 1710899220
transform 1 0 1284 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2058
timestamp 1710899220
transform 1 0 2164 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2059
timestamp 1710899220
transform 1 0 1972 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2060
timestamp 1710899220
transform 1 0 1500 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2061
timestamp 1710899220
transform 1 0 1372 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2062
timestamp 1710899220
transform 1 0 1348 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2063
timestamp 1710899220
transform 1 0 1196 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2064
timestamp 1710899220
transform 1 0 1516 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2065
timestamp 1710899220
transform 1 0 1436 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2066
timestamp 1710899220
transform 1 0 1356 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2067
timestamp 1710899220
transform 1 0 1260 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2068
timestamp 1710899220
transform 1 0 1268 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_2069
timestamp 1710899220
transform 1 0 188 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_2070
timestamp 1710899220
transform 1 0 1460 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2071
timestamp 1710899220
transform 1 0 1380 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2072
timestamp 1710899220
transform 1 0 1292 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2073
timestamp 1710899220
transform 1 0 1260 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2074
timestamp 1710899220
transform 1 0 1252 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2075
timestamp 1710899220
transform 1 0 1004 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2076
timestamp 1710899220
transform 1 0 1292 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_2077
timestamp 1710899220
transform 1 0 1292 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2078
timestamp 1710899220
transform 1 0 1236 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2079
timestamp 1710899220
transform 1 0 172 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_2080
timestamp 1710899220
transform 1 0 1284 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2081
timestamp 1710899220
transform 1 0 1268 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2082
timestamp 1710899220
transform 1 0 1228 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2083
timestamp 1710899220
transform 1 0 1108 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2084
timestamp 1710899220
transform 1 0 252 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2085
timestamp 1710899220
transform 1 0 1284 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2086
timestamp 1710899220
transform 1 0 1188 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2087
timestamp 1710899220
transform 1 0 1668 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2088
timestamp 1710899220
transform 1 0 1596 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2089
timestamp 1710899220
transform 1 0 1220 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2090
timestamp 1710899220
transform 1 0 1716 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_2091
timestamp 1710899220
transform 1 0 1676 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_2092
timestamp 1710899220
transform 1 0 1508 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2093
timestamp 1710899220
transform 1 0 1436 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2094
timestamp 1710899220
transform 1 0 1588 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2095
timestamp 1710899220
transform 1 0 1420 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2096
timestamp 1710899220
transform 1 0 1348 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2097
timestamp 1710899220
transform 1 0 1252 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2098
timestamp 1710899220
transform 1 0 1236 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2099
timestamp 1710899220
transform 1 0 1532 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2100
timestamp 1710899220
transform 1 0 1484 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2101
timestamp 1710899220
transform 1 0 1412 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2102
timestamp 1710899220
transform 1 0 1356 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2103
timestamp 1710899220
transform 1 0 1084 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2104
timestamp 1710899220
transform 1 0 924 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2105
timestamp 1710899220
transform 1 0 908 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2106
timestamp 1710899220
transform 1 0 844 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2107
timestamp 1710899220
transform 1 0 956 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2108
timestamp 1710899220
transform 1 0 844 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2109
timestamp 1710899220
transform 1 0 908 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2110
timestamp 1710899220
transform 1 0 892 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2111
timestamp 1710899220
transform 1 0 796 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2112
timestamp 1710899220
transform 1 0 772 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2113
timestamp 1710899220
transform 1 0 1100 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2114
timestamp 1710899220
transform 1 0 1036 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2115
timestamp 1710899220
transform 1 0 948 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2116
timestamp 1710899220
transform 1 0 1116 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2117
timestamp 1710899220
transform 1 0 1060 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2118
timestamp 1710899220
transform 1 0 1044 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_2119
timestamp 1710899220
transform 1 0 1044 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2120
timestamp 1710899220
transform 1 0 988 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_2121
timestamp 1710899220
transform 1 0 964 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2122
timestamp 1710899220
transform 1 0 1156 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2123
timestamp 1710899220
transform 1 0 1092 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2124
timestamp 1710899220
transform 1 0 1092 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2125
timestamp 1710899220
transform 1 0 884 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2126
timestamp 1710899220
transform 1 0 1172 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2127
timestamp 1710899220
transform 1 0 988 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2128
timestamp 1710899220
transform 1 0 1004 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2129
timestamp 1710899220
transform 1 0 980 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2130
timestamp 1710899220
transform 1 0 980 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2131
timestamp 1710899220
transform 1 0 940 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2132
timestamp 1710899220
transform 1 0 1124 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2133
timestamp 1710899220
transform 1 0 1012 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2134
timestamp 1710899220
transform 1 0 900 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2135
timestamp 1710899220
transform 1 0 852 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2136
timestamp 1710899220
transform 1 0 876 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2137
timestamp 1710899220
transform 1 0 836 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2138
timestamp 1710899220
transform 1 0 796 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2139
timestamp 1710899220
transform 1 0 852 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_2140
timestamp 1710899220
transform 1 0 828 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_2141
timestamp 1710899220
transform 1 0 828 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2142
timestamp 1710899220
transform 1 0 788 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2143
timestamp 1710899220
transform 1 0 1052 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2144
timestamp 1710899220
transform 1 0 988 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2145
timestamp 1710899220
transform 1 0 1084 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2146
timestamp 1710899220
transform 1 0 1052 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2147
timestamp 1710899220
transform 1 0 1028 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2148
timestamp 1710899220
transform 1 0 740 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2149
timestamp 1710899220
transform 1 0 948 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_2150
timestamp 1710899220
transform 1 0 780 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_2151
timestamp 1710899220
transform 1 0 1036 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_2152
timestamp 1710899220
transform 1 0 892 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_2153
timestamp 1710899220
transform 1 0 860 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2154
timestamp 1710899220
transform 1 0 804 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2155
timestamp 1710899220
transform 1 0 892 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2156
timestamp 1710899220
transform 1 0 876 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2157
timestamp 1710899220
transform 1 0 924 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2158
timestamp 1710899220
transform 1 0 876 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2159
timestamp 1710899220
transform 1 0 812 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2160
timestamp 1710899220
transform 1 0 764 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2161
timestamp 1710899220
transform 1 0 828 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2162
timestamp 1710899220
transform 1 0 812 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_2163
timestamp 1710899220
transform 1 0 804 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2164
timestamp 1710899220
transform 1 0 756 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_2165
timestamp 1710899220
transform 1 0 1028 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2166
timestamp 1710899220
transform 1 0 964 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2167
timestamp 1710899220
transform 1 0 1036 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2168
timestamp 1710899220
transform 1 0 964 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2169
timestamp 1710899220
transform 1 0 1068 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2170
timestamp 1710899220
transform 1 0 1012 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2171
timestamp 1710899220
transform 1 0 1004 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2172
timestamp 1710899220
transform 1 0 972 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2173
timestamp 1710899220
transform 1 0 916 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2174
timestamp 1710899220
transform 1 0 1044 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2175
timestamp 1710899220
transform 1 0 1020 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2176
timestamp 1710899220
transform 1 0 932 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2177
timestamp 1710899220
transform 1 0 844 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2178
timestamp 1710899220
transform 1 0 916 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2179
timestamp 1710899220
transform 1 0 876 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2180
timestamp 1710899220
transform 1 0 932 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2181
timestamp 1710899220
transform 1 0 876 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2182
timestamp 1710899220
transform 1 0 844 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2183
timestamp 1710899220
transform 1 0 836 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2184
timestamp 1710899220
transform 1 0 788 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2185
timestamp 1710899220
transform 1 0 1052 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2186
timestamp 1710899220
transform 1 0 1004 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2187
timestamp 1710899220
transform 1 0 1020 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_2188
timestamp 1710899220
transform 1 0 860 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_2189
timestamp 1710899220
transform 1 0 988 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2190
timestamp 1710899220
transform 1 0 900 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2191
timestamp 1710899220
transform 1 0 868 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2192
timestamp 1710899220
transform 1 0 804 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2193
timestamp 1710899220
transform 1 0 756 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2194
timestamp 1710899220
transform 1 0 708 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2195
timestamp 1710899220
transform 1 0 764 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2196
timestamp 1710899220
transform 1 0 724 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2197
timestamp 1710899220
transform 1 0 764 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2198
timestamp 1710899220
transform 1 0 700 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2199
timestamp 1710899220
transform 1 0 756 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2200
timestamp 1710899220
transform 1 0 708 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2201
timestamp 1710899220
transform 1 0 868 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2202
timestamp 1710899220
transform 1 0 796 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2203
timestamp 1710899220
transform 1 0 908 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2204
timestamp 1710899220
transform 1 0 876 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2205
timestamp 1710899220
transform 1 0 788 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2206
timestamp 1710899220
transform 1 0 708 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2207
timestamp 1710899220
transform 1 0 676 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2208
timestamp 1710899220
transform 1 0 532 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2209
timestamp 1710899220
transform 1 0 676 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2210
timestamp 1710899220
transform 1 0 652 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2211
timestamp 1710899220
transform 1 0 724 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2212
timestamp 1710899220
transform 1 0 708 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2213
timestamp 1710899220
transform 1 0 684 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2214
timestamp 1710899220
transform 1 0 660 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2215
timestamp 1710899220
transform 1 0 620 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2216
timestamp 1710899220
transform 1 0 612 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2217
timestamp 1710899220
transform 1 0 588 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2218
timestamp 1710899220
transform 1 0 628 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_2219
timestamp 1710899220
transform 1 0 628 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2220
timestamp 1710899220
transform 1 0 556 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_2221
timestamp 1710899220
transform 1 0 516 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_2222
timestamp 1710899220
transform 1 0 516 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2223
timestamp 1710899220
transform 1 0 660 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2224
timestamp 1710899220
transform 1 0 660 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2225
timestamp 1710899220
transform 1 0 596 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2226
timestamp 1710899220
transform 1 0 540 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2227
timestamp 1710899220
transform 1 0 524 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2228
timestamp 1710899220
transform 1 0 732 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2229
timestamp 1710899220
transform 1 0 652 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2230
timestamp 1710899220
transform 1 0 716 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2231
timestamp 1710899220
transform 1 0 700 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2232
timestamp 1710899220
transform 1 0 724 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2233
timestamp 1710899220
transform 1 0 628 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2234
timestamp 1710899220
transform 1 0 700 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2235
timestamp 1710899220
transform 1 0 588 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2236
timestamp 1710899220
transform 1 0 612 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2237
timestamp 1710899220
transform 1 0 532 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2238
timestamp 1710899220
transform 1 0 612 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2239
timestamp 1710899220
transform 1 0 572 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2240
timestamp 1710899220
transform 1 0 556 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2241
timestamp 1710899220
transform 1 0 548 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2242
timestamp 1710899220
transform 1 0 764 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2243
timestamp 1710899220
transform 1 0 628 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2244
timestamp 1710899220
transform 1 0 716 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2245
timestamp 1710899220
transform 1 0 652 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2246
timestamp 1710899220
transform 1 0 596 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2247
timestamp 1710899220
transform 1 0 524 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2248
timestamp 1710899220
transform 1 0 228 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2249
timestamp 1710899220
transform 1 0 212 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2250
timestamp 1710899220
transform 1 0 324 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_2251
timestamp 1710899220
transform 1 0 180 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_2252
timestamp 1710899220
transform 1 0 284 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2253
timestamp 1710899220
transform 1 0 188 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2254
timestamp 1710899220
transform 1 0 604 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_2255
timestamp 1710899220
transform 1 0 268 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_2256
timestamp 1710899220
transform 1 0 396 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2257
timestamp 1710899220
transform 1 0 268 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2258
timestamp 1710899220
transform 1 0 468 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2259
timestamp 1710899220
transform 1 0 372 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2260
timestamp 1710899220
transform 1 0 588 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2261
timestamp 1710899220
transform 1 0 548 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2262
timestamp 1710899220
transform 1 0 548 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_2263
timestamp 1710899220
transform 1 0 452 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_2264
timestamp 1710899220
transform 1 0 380 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2265
timestamp 1710899220
transform 1 0 356 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_2266
timestamp 1710899220
transform 1 0 348 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2267
timestamp 1710899220
transform 1 0 628 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2268
timestamp 1710899220
transform 1 0 572 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2269
timestamp 1710899220
transform 1 0 484 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2270
timestamp 1710899220
transform 1 0 420 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2271
timestamp 1710899220
transform 1 0 380 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2272
timestamp 1710899220
transform 1 0 364 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2273
timestamp 1710899220
transform 1 0 628 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2274
timestamp 1710899220
transform 1 0 604 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_2275
timestamp 1710899220
transform 1 0 540 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2276
timestamp 1710899220
transform 1 0 452 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2277
timestamp 1710899220
transform 1 0 436 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_2278
timestamp 1710899220
transform 1 0 420 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2279
timestamp 1710899220
transform 1 0 644 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2280
timestamp 1710899220
transform 1 0 556 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2281
timestamp 1710899220
transform 1 0 492 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2282
timestamp 1710899220
transform 1 0 476 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2283
timestamp 1710899220
transform 1 0 476 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2284
timestamp 1710899220
transform 1 0 476 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2285
timestamp 1710899220
transform 1 0 436 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2286
timestamp 1710899220
transform 1 0 628 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2287
timestamp 1710899220
transform 1 0 596 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2288
timestamp 1710899220
transform 1 0 532 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2289
timestamp 1710899220
transform 1 0 292 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2290
timestamp 1710899220
transform 1 0 364 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2291
timestamp 1710899220
transform 1 0 300 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2292
timestamp 1710899220
transform 1 0 428 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_2293
timestamp 1710899220
transform 1 0 340 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_2294
timestamp 1710899220
transform 1 0 548 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_2295
timestamp 1710899220
transform 1 0 492 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_2296
timestamp 1710899220
transform 1 0 564 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2297
timestamp 1710899220
transform 1 0 508 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2298
timestamp 1710899220
transform 1 0 524 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2299
timestamp 1710899220
transform 1 0 276 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2300
timestamp 1710899220
transform 1 0 332 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_2301
timestamp 1710899220
transform 1 0 292 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_2302
timestamp 1710899220
transform 1 0 428 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2303
timestamp 1710899220
transform 1 0 300 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2304
timestamp 1710899220
transform 1 0 372 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2305
timestamp 1710899220
transform 1 0 308 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2306
timestamp 1710899220
transform 1 0 500 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2307
timestamp 1710899220
transform 1 0 492 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2308
timestamp 1710899220
transform 1 0 468 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2309
timestamp 1710899220
transform 1 0 468 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2310
timestamp 1710899220
transform 1 0 516 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2311
timestamp 1710899220
transform 1 0 476 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2312
timestamp 1710899220
transform 1 0 164 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2313
timestamp 1710899220
transform 1 0 148 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2314
timestamp 1710899220
transform 1 0 252 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_2315
timestamp 1710899220
transform 1 0 188 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2316
timestamp 1710899220
transform 1 0 276 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_2317
timestamp 1710899220
transform 1 0 196 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_2318
timestamp 1710899220
transform 1 0 308 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2319
timestamp 1710899220
transform 1 0 252 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2320
timestamp 1710899220
transform 1 0 468 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_2321
timestamp 1710899220
transform 1 0 284 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_2322
timestamp 1710899220
transform 1 0 364 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2323
timestamp 1710899220
transform 1 0 292 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2324
timestamp 1710899220
transform 1 0 380 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2325
timestamp 1710899220
transform 1 0 340 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2326
timestamp 1710899220
transform 1 0 420 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2327
timestamp 1710899220
transform 1 0 388 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2328
timestamp 1710899220
transform 1 0 380 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2329
timestamp 1710899220
transform 1 0 356 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2330
timestamp 1710899220
transform 1 0 340 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2331
timestamp 1710899220
transform 1 0 444 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2332
timestamp 1710899220
transform 1 0 412 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2333
timestamp 1710899220
transform 1 0 468 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2334
timestamp 1710899220
transform 1 0 428 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2335
timestamp 1710899220
transform 1 0 468 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2336
timestamp 1710899220
transform 1 0 284 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2337
timestamp 1710899220
transform 1 0 380 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2338
timestamp 1710899220
transform 1 0 292 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2339
timestamp 1710899220
transform 1 0 300 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2340
timestamp 1710899220
transform 1 0 228 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2341
timestamp 1710899220
transform 1 0 420 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2342
timestamp 1710899220
transform 1 0 236 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2343
timestamp 1710899220
transform 1 0 348 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2344
timestamp 1710899220
transform 1 0 252 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2345
timestamp 1710899220
transform 1 0 468 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2346
timestamp 1710899220
transform 1 0 284 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2347
timestamp 1710899220
transform 1 0 412 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2348
timestamp 1710899220
transform 1 0 292 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2349
timestamp 1710899220
transform 1 0 300 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2350
timestamp 1710899220
transform 1 0 188 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2351
timestamp 1710899220
transform 1 0 324 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2352
timestamp 1710899220
transform 1 0 220 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2353
timestamp 1710899220
transform 1 0 460 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2354
timestamp 1710899220
transform 1 0 276 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2355
timestamp 1710899220
transform 1 0 372 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2356
timestamp 1710899220
transform 1 0 284 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2357
timestamp 1710899220
transform 1 0 252 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_2358
timestamp 1710899220
transform 1 0 204 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_2359
timestamp 1710899220
transform 1 0 268 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2360
timestamp 1710899220
transform 1 0 212 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2361
timestamp 1710899220
transform 1 0 508 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_2362
timestamp 1710899220
transform 1 0 252 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_2363
timestamp 1710899220
transform 1 0 308 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2364
timestamp 1710899220
transform 1 0 260 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2365
timestamp 1710899220
transform 1 0 484 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_2366
timestamp 1710899220
transform 1 0 284 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_2367
timestamp 1710899220
transform 1 0 404 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2368
timestamp 1710899220
transform 1 0 292 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2369
timestamp 1710899220
transform 1 0 636 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2370
timestamp 1710899220
transform 1 0 580 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2371
timestamp 1710899220
transform 1 0 380 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2372
timestamp 1710899220
transform 1 0 372 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2373
timestamp 1710899220
transform 1 0 364 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2374
timestamp 1710899220
transform 1 0 676 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2375
timestamp 1710899220
transform 1 0 652 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2376
timestamp 1710899220
transform 1 0 652 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2377
timestamp 1710899220
transform 1 0 612 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2378
timestamp 1710899220
transform 1 0 412 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2379
timestamp 1710899220
transform 1 0 388 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2380
timestamp 1710899220
transform 1 0 348 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2381
timestamp 1710899220
transform 1 0 580 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2382
timestamp 1710899220
transform 1 0 548 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2383
timestamp 1710899220
transform 1 0 532 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2384
timestamp 1710899220
transform 1 0 468 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2385
timestamp 1710899220
transform 1 0 444 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2386
timestamp 1710899220
transform 1 0 612 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2387
timestamp 1710899220
transform 1 0 564 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2388
timestamp 1710899220
transform 1 0 564 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2389
timestamp 1710899220
transform 1 0 492 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2390
timestamp 1710899220
transform 1 0 468 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2391
timestamp 1710899220
transform 1 0 460 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2392
timestamp 1710899220
transform 1 0 452 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2393
timestamp 1710899220
transform 1 0 428 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2394
timestamp 1710899220
transform 1 0 564 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2395
timestamp 1710899220
transform 1 0 508 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2396
timestamp 1710899220
transform 1 0 644 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_2397
timestamp 1710899220
transform 1 0 500 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_2398
timestamp 1710899220
transform 1 0 516 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2399
timestamp 1710899220
transform 1 0 220 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2400
timestamp 1710899220
transform 1 0 340 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2401
timestamp 1710899220
transform 1 0 228 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2402
timestamp 1710899220
transform 1 0 444 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2403
timestamp 1710899220
transform 1 0 300 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2404
timestamp 1710899220
transform 1 0 356 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2405
timestamp 1710899220
transform 1 0 324 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2406
timestamp 1710899220
transform 1 0 548 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2407
timestamp 1710899220
transform 1 0 500 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2408
timestamp 1710899220
transform 1 0 612 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2409
timestamp 1710899220
transform 1 0 508 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2410
timestamp 1710899220
transform 1 0 300 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2411
timestamp 1710899220
transform 1 0 228 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2412
timestamp 1710899220
transform 1 0 420 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2413
timestamp 1710899220
transform 1 0 284 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2414
timestamp 1710899220
transform 1 0 340 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2415
timestamp 1710899220
transform 1 0 308 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2416
timestamp 1710899220
transform 1 0 460 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_2417
timestamp 1710899220
transform 1 0 236 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_2418
timestamp 1710899220
transform 1 0 380 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2419
timestamp 1710899220
transform 1 0 244 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2420
timestamp 1710899220
transform 1 0 2292 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2421
timestamp 1710899220
transform 1 0 2212 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2422
timestamp 1710899220
transform 1 0 1916 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2423
timestamp 1710899220
transform 1 0 1836 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2424
timestamp 1710899220
transform 1 0 1868 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2425
timestamp 1710899220
transform 1 0 1804 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2426
timestamp 1710899220
transform 1 0 692 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2427
timestamp 1710899220
transform 1 0 644 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2428
timestamp 1710899220
transform 1 0 356 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_2429
timestamp 1710899220
transform 1 0 292 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2430
timestamp 1710899220
transform 1 0 324 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2431
timestamp 1710899220
transform 1 0 228 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2432
timestamp 1710899220
transform 1 0 292 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2433
timestamp 1710899220
transform 1 0 236 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2434
timestamp 1710899220
transform 1 0 1196 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_2435
timestamp 1710899220
transform 1 0 1140 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_2436
timestamp 1710899220
transform 1 0 1012 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2437
timestamp 1710899220
transform 1 0 972 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2438
timestamp 1710899220
transform 1 0 852 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2439
timestamp 1710899220
transform 1 0 796 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2440
timestamp 1710899220
transform 1 0 324 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2441
timestamp 1710899220
transform 1 0 228 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2442
timestamp 1710899220
transform 1 0 356 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2443
timestamp 1710899220
transform 1 0 292 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2444
timestamp 1710899220
transform 1 0 1748 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2445
timestamp 1710899220
transform 1 0 1676 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2446
timestamp 1710899220
transform 1 0 1700 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_2447
timestamp 1710899220
transform 1 0 1676 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_2448
timestamp 1710899220
transform 1 0 2076 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2449
timestamp 1710899220
transform 1 0 2004 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2450
timestamp 1710899220
transform 1 0 2068 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2451
timestamp 1710899220
transform 1 0 1996 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2452
timestamp 1710899220
transform 1 0 1820 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_2453
timestamp 1710899220
transform 1 0 1724 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_2454
timestamp 1710899220
transform 1 0 1940 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2455
timestamp 1710899220
transform 1 0 1868 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2456
timestamp 1710899220
transform 1 0 2044 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2457
timestamp 1710899220
transform 1 0 1980 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2458
timestamp 1710899220
transform 1 0 2068 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2459
timestamp 1710899220
transform 1 0 1980 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2460
timestamp 1710899220
transform 1 0 2092 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2461
timestamp 1710899220
transform 1 0 2020 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2462
timestamp 1710899220
transform 1 0 1484 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2463
timestamp 1710899220
transform 1 0 1452 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2464
timestamp 1710899220
transform 1 0 1996 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2465
timestamp 1710899220
transform 1 0 1844 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2466
timestamp 1710899220
transform 1 0 1868 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2467
timestamp 1710899220
transform 1 0 1788 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2468
timestamp 1710899220
transform 1 0 1876 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2469
timestamp 1710899220
transform 1 0 1780 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2470
timestamp 1710899220
transform 1 0 1884 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2471
timestamp 1710899220
transform 1 0 1836 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2472
timestamp 1710899220
transform 1 0 1804 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2473
timestamp 1710899220
transform 1 0 1788 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2474
timestamp 1710899220
transform 1 0 1548 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2475
timestamp 1710899220
transform 1 0 1500 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2476
timestamp 1710899220
transform 1 0 1188 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2477
timestamp 1710899220
transform 1 0 1124 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2478
timestamp 1710899220
transform 1 0 852 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2479
timestamp 1710899220
transform 1 0 804 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2480
timestamp 1710899220
transform 1 0 988 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2481
timestamp 1710899220
transform 1 0 900 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2482
timestamp 1710899220
transform 1 0 1188 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2483
timestamp 1710899220
transform 1 0 1116 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2484
timestamp 1710899220
transform 1 0 556 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2485
timestamp 1710899220
transform 1 0 500 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2486
timestamp 1710899220
transform 1 0 532 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_2487
timestamp 1710899220
transform 1 0 460 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_2488
timestamp 1710899220
transform 1 0 628 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2489
timestamp 1710899220
transform 1 0 604 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2490
timestamp 1710899220
transform 1 0 692 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2491
timestamp 1710899220
transform 1 0 628 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2492
timestamp 1710899220
transform 1 0 1348 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2493
timestamp 1710899220
transform 1 0 1276 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2494
timestamp 1710899220
transform 1 0 1476 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2495
timestamp 1710899220
transform 1 0 1412 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2496
timestamp 1710899220
transform 1 0 1324 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2497
timestamp 1710899220
transform 1 0 1260 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2498
timestamp 1710899220
transform 1 0 2468 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2499
timestamp 1710899220
transform 1 0 2436 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2500
timestamp 1710899220
transform 1 0 2356 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_2501
timestamp 1710899220
transform 1 0 2164 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_2502
timestamp 1710899220
transform 1 0 2564 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2503
timestamp 1710899220
transform 1 0 2540 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2504
timestamp 1710899220
transform 1 0 2556 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2505
timestamp 1710899220
transform 1 0 2524 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2506
timestamp 1710899220
transform 1 0 2508 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2507
timestamp 1710899220
transform 1 0 2428 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2508
timestamp 1710899220
transform 1 0 2428 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_2509
timestamp 1710899220
transform 1 0 2380 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_2510
timestamp 1710899220
transform 1 0 2372 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2511
timestamp 1710899220
transform 1 0 2620 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2512
timestamp 1710899220
transform 1 0 2548 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2513
timestamp 1710899220
transform 1 0 2324 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2514
timestamp 1710899220
transform 1 0 2212 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2515
timestamp 1710899220
transform 1 0 2308 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2516
timestamp 1710899220
transform 1 0 2260 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2517
timestamp 1710899220
transform 1 0 2268 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2518
timestamp 1710899220
transform 1 0 2204 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2519
timestamp 1710899220
transform 1 0 2492 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_2520
timestamp 1710899220
transform 1 0 2284 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_2521
timestamp 1710899220
transform 1 0 2292 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2522
timestamp 1710899220
transform 1 0 2268 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2523
timestamp 1710899220
transform 1 0 2372 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2524
timestamp 1710899220
transform 1 0 2260 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2525
timestamp 1710899220
transform 1 0 2380 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2526
timestamp 1710899220
transform 1 0 2332 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2527
timestamp 1710899220
transform 1 0 2444 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2528
timestamp 1710899220
transform 1 0 2364 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2529
timestamp 1710899220
transform 1 0 2244 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2530
timestamp 1710899220
transform 1 0 2364 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_2531
timestamp 1710899220
transform 1 0 2316 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_2532
timestamp 1710899220
transform 1 0 2548 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2533
timestamp 1710899220
transform 1 0 2452 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2534
timestamp 1710899220
transform 1 0 2532 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2535
timestamp 1710899220
transform 1 0 2484 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2536
timestamp 1710899220
transform 1 0 2452 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2537
timestamp 1710899220
transform 1 0 2612 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2538
timestamp 1710899220
transform 1 0 2532 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2539
timestamp 1710899220
transform 1 0 2572 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2540
timestamp 1710899220
transform 1 0 2532 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2541
timestamp 1710899220
transform 1 0 2356 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2542
timestamp 1710899220
transform 1 0 2316 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2543
timestamp 1710899220
transform 1 0 2428 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2544
timestamp 1710899220
transform 1 0 2348 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2545
timestamp 1710899220
transform 1 0 2612 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2546
timestamp 1710899220
transform 1 0 2596 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2547
timestamp 1710899220
transform 1 0 2596 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2548
timestamp 1710899220
transform 1 0 2532 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2549
timestamp 1710899220
transform 1 0 2444 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2550
timestamp 1710899220
transform 1 0 2492 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2551
timestamp 1710899220
transform 1 0 2396 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2552
timestamp 1710899220
transform 1 0 2564 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2553
timestamp 1710899220
transform 1 0 2476 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2554
timestamp 1710899220
transform 1 0 2492 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2555
timestamp 1710899220
transform 1 0 2436 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2556
timestamp 1710899220
transform 1 0 2364 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2557
timestamp 1710899220
transform 1 0 2324 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2558
timestamp 1710899220
transform 1 0 2300 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2559
timestamp 1710899220
transform 1 0 2380 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2560
timestamp 1710899220
transform 1 0 2324 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2561
timestamp 1710899220
transform 1 0 2644 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2562
timestamp 1710899220
transform 1 0 2532 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2563
timestamp 1710899220
transform 1 0 2500 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2564
timestamp 1710899220
transform 1 0 2364 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2565
timestamp 1710899220
transform 1 0 2580 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2566
timestamp 1710899220
transform 1 0 2484 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2567
timestamp 1710899220
transform 1 0 2636 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2568
timestamp 1710899220
transform 1 0 2540 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2569
timestamp 1710899220
transform 1 0 2612 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2570
timestamp 1710899220
transform 1 0 2556 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2571
timestamp 1710899220
transform 1 0 2236 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2572
timestamp 1710899220
transform 1 0 2132 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2573
timestamp 1710899220
transform 1 0 2300 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2574
timestamp 1710899220
transform 1 0 2188 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2575
timestamp 1710899220
transform 1 0 2332 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2576
timestamp 1710899220
transform 1 0 2252 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2577
timestamp 1710899220
transform 1 0 2036 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2578
timestamp 1710899220
transform 1 0 1980 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2579
timestamp 1710899220
transform 1 0 2124 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_2580
timestamp 1710899220
transform 1 0 2044 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_2581
timestamp 1710899220
transform 1 0 2260 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_2582
timestamp 1710899220
transform 1 0 2220 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_2583
timestamp 1710899220
transform 1 0 2116 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_2584
timestamp 1710899220
transform 1 0 2260 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_2585
timestamp 1710899220
transform 1 0 2156 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_2586
timestamp 1710899220
transform 1 0 2172 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2587
timestamp 1710899220
transform 1 0 2116 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2588
timestamp 1710899220
transform 1 0 2028 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2589
timestamp 1710899220
transform 1 0 1492 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2590
timestamp 1710899220
transform 1 0 1380 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2591
timestamp 1710899220
transform 1 0 1684 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2592
timestamp 1710899220
transform 1 0 1524 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2593
timestamp 1710899220
transform 1 0 1764 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_2594
timestamp 1710899220
transform 1 0 1628 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_2595
timestamp 1710899220
transform 1 0 1164 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_2596
timestamp 1710899220
transform 1 0 1324 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2597
timestamp 1710899220
transform 1 0 1012 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2598
timestamp 1710899220
transform 1 0 1284 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_2599
timestamp 1710899220
transform 1 0 1140 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_2600
timestamp 1710899220
transform 1 0 2468 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2601
timestamp 1710899220
transform 1 0 2468 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2602
timestamp 1710899220
transform 1 0 2412 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2603
timestamp 1710899220
transform 1 0 2332 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_2604
timestamp 1710899220
transform 1 0 2220 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_2605
timestamp 1710899220
transform 1 0 2668 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2606
timestamp 1710899220
transform 1 0 2572 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2607
timestamp 1710899220
transform 1 0 2332 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2608
timestamp 1710899220
transform 1 0 2148 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2609
timestamp 1710899220
transform 1 0 2044 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2610
timestamp 1710899220
transform 1 0 2124 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2611
timestamp 1710899220
transform 1 0 2012 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2612
timestamp 1710899220
transform 1 0 2100 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2613
timestamp 1710899220
transform 1 0 1996 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2614
timestamp 1710899220
transform 1 0 1572 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2615
timestamp 1710899220
transform 1 0 1996 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2616
timestamp 1710899220
transform 1 0 1900 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2617
timestamp 1710899220
transform 1 0 1652 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2618
timestamp 1710899220
transform 1 0 1588 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2619
timestamp 1710899220
transform 1 0 1556 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2620
timestamp 1710899220
transform 1 0 2124 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2621
timestamp 1710899220
transform 1 0 2020 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2622
timestamp 1710899220
transform 1 0 2132 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2623
timestamp 1710899220
transform 1 0 2028 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2624
timestamp 1710899220
transform 1 0 1756 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2625
timestamp 1710899220
transform 1 0 1708 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2626
timestamp 1710899220
transform 1 0 1644 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2627
timestamp 1710899220
transform 1 0 1612 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2628
timestamp 1710899220
transform 1 0 1612 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2629
timestamp 1710899220
transform 1 0 1556 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2630
timestamp 1710899220
transform 1 0 1804 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2631
timestamp 1710899220
transform 1 0 1700 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2632
timestamp 1710899220
transform 1 0 1588 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2633
timestamp 1710899220
transform 1 0 1212 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_2634
timestamp 1710899220
transform 1 0 1036 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_2635
timestamp 1710899220
transform 1 0 964 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_2636
timestamp 1710899220
transform 1 0 1140 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2637
timestamp 1710899220
transform 1 0 1068 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_2638
timestamp 1710899220
transform 1 0 1068 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2639
timestamp 1710899220
transform 1 0 892 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_2640
timestamp 1710899220
transform 1 0 1044 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2641
timestamp 1710899220
transform 1 0 1020 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2642
timestamp 1710899220
transform 1 0 1020 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2643
timestamp 1710899220
transform 1 0 956 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2644
timestamp 1710899220
transform 1 0 924 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2645
timestamp 1710899220
transform 1 0 468 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2646
timestamp 1710899220
transform 1 0 340 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2647
timestamp 1710899220
transform 1 0 300 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2648
timestamp 1710899220
transform 1 0 532 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2649
timestamp 1710899220
transform 1 0 492 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2650
timestamp 1710899220
transform 1 0 1004 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2651
timestamp 1710899220
transform 1 0 908 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_2652
timestamp 1710899220
transform 1 0 852 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2653
timestamp 1710899220
transform 1 0 852 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_2654
timestamp 1710899220
transform 1 0 1012 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2655
timestamp 1710899220
transform 1 0 932 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2656
timestamp 1710899220
transform 1 0 1252 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_2657
timestamp 1710899220
transform 1 0 1116 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_2658
timestamp 1710899220
transform 1 0 964 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_2659
timestamp 1710899220
transform 1 0 556 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2660
timestamp 1710899220
transform 1 0 308 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2661
timestamp 1710899220
transform 1 0 388 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2662
timestamp 1710899220
transform 1 0 356 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2663
timestamp 1710899220
transform 1 0 300 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2664
timestamp 1710899220
transform 1 0 508 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2665
timestamp 1710899220
transform 1 0 436 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2666
timestamp 1710899220
transform 1 0 380 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2667
timestamp 1710899220
transform 1 0 332 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2668
timestamp 1710899220
transform 1 0 2052 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2669
timestamp 1710899220
transform 1 0 1948 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2670
timestamp 1710899220
transform 1 0 1916 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2671
timestamp 1710899220
transform 1 0 1820 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2672
timestamp 1710899220
transform 1 0 1596 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2673
timestamp 1710899220
transform 1 0 1524 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2674
timestamp 1710899220
transform 1 0 1484 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2675
timestamp 1710899220
transform 1 0 1484 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2676
timestamp 1710899220
transform 1 0 1452 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2677
timestamp 1710899220
transform 1 0 1396 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2678
timestamp 1710899220
transform 1 0 1516 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2679
timestamp 1710899220
transform 1 0 1372 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2680
timestamp 1710899220
transform 1 0 1932 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2681
timestamp 1710899220
transform 1 0 1836 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2682
timestamp 1710899220
transform 1 0 1940 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_2683
timestamp 1710899220
transform 1 0 1884 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_2684
timestamp 1710899220
transform 1 0 1844 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2685
timestamp 1710899220
transform 1 0 1780 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2686
timestamp 1710899220
transform 1 0 1436 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2687
timestamp 1710899220
transform 1 0 1396 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2688
timestamp 1710899220
transform 1 0 1252 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2689
timestamp 1710899220
transform 1 0 1252 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2690
timestamp 1710899220
transform 1 0 1212 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2691
timestamp 1710899220
transform 1 0 1212 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2692
timestamp 1710899220
transform 1 0 1068 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2693
timestamp 1710899220
transform 1 0 1596 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2694
timestamp 1710899220
transform 1 0 1508 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2695
timestamp 1710899220
transform 1 0 1348 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2696
timestamp 1710899220
transform 1 0 1204 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2697
timestamp 1710899220
transform 1 0 1076 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2698
timestamp 1710899220
transform 1 0 1076 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2699
timestamp 1710899220
transform 1 0 1028 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_2700
timestamp 1710899220
transform 1 0 1028 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2701
timestamp 1710899220
transform 1 0 1140 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2702
timestamp 1710899220
transform 1 0 1132 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2703
timestamp 1710899220
transform 1 0 1052 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2704
timestamp 1710899220
transform 1 0 1044 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2705
timestamp 1710899220
transform 1 0 852 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2706
timestamp 1710899220
transform 1 0 780 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2707
timestamp 1710899220
transform 1 0 708 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2708
timestamp 1710899220
transform 1 0 740 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2709
timestamp 1710899220
transform 1 0 692 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2710
timestamp 1710899220
transform 1 0 644 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2711
timestamp 1710899220
transform 1 0 596 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2712
timestamp 1710899220
transform 1 0 948 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_2713
timestamp 1710899220
transform 1 0 900 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_2714
timestamp 1710899220
transform 1 0 1388 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2715
timestamp 1710899220
transform 1 0 1236 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2716
timestamp 1710899220
transform 1 0 1140 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2717
timestamp 1710899220
transform 1 0 1100 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2718
timestamp 1710899220
transform 1 0 532 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2719
timestamp 1710899220
transform 1 0 468 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2720
timestamp 1710899220
transform 1 0 476 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2721
timestamp 1710899220
transform 1 0 412 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2722
timestamp 1710899220
transform 1 0 636 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2723
timestamp 1710899220
transform 1 0 588 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2724
timestamp 1710899220
transform 1 0 532 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2725
timestamp 1710899220
transform 1 0 492 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2726
timestamp 1710899220
transform 1 0 492 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2727
timestamp 1710899220
transform 1 0 1084 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2728
timestamp 1710899220
transform 1 0 724 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2729
timestamp 1710899220
transform 1 0 716 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2730
timestamp 1710899220
transform 1 0 660 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2731
timestamp 1710899220
transform 1 0 660 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2732
timestamp 1710899220
transform 1 0 580 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2733
timestamp 1710899220
transform 1 0 1964 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2734
timestamp 1710899220
transform 1 0 1836 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2735
timestamp 1710899220
transform 1 0 1924 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2736
timestamp 1710899220
transform 1 0 1820 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2737
timestamp 1710899220
transform 1 0 2300 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2738
timestamp 1710899220
transform 1 0 2244 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2739
timestamp 1710899220
transform 1 0 2428 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2740
timestamp 1710899220
transform 1 0 2308 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2741
timestamp 1710899220
transform 1 0 2172 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2742
timestamp 1710899220
transform 1 0 2116 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2743
timestamp 1710899220
transform 1 0 2332 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_2744
timestamp 1710899220
transform 1 0 2204 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_2745
timestamp 1710899220
transform 1 0 2140 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_2746
timestamp 1710899220
transform 1 0 2076 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_2747
timestamp 1710899220
transform 1 0 1964 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2748
timestamp 1710899220
transform 1 0 1908 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2749
timestamp 1710899220
transform 1 0 1924 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2750
timestamp 1710899220
transform 1 0 1852 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2751
timestamp 1710899220
transform 1 0 1964 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2752
timestamp 1710899220
transform 1 0 1908 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2753
timestamp 1710899220
transform 1 0 1964 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_2754
timestamp 1710899220
transform 1 0 1908 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_2755
timestamp 1710899220
transform 1 0 1988 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_2756
timestamp 1710899220
transform 1 0 1924 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_2757
timestamp 1710899220
transform 1 0 2292 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_2758
timestamp 1710899220
transform 1 0 2180 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_2759
timestamp 1710899220
transform 1 0 2068 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_2760
timestamp 1710899220
transform 1 0 2148 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_2761
timestamp 1710899220
transform 1 0 2060 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_2762
timestamp 1710899220
transform 1 0 2412 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_2763
timestamp 1710899220
transform 1 0 2284 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_2764
timestamp 1710899220
transform 1 0 2156 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_2765
timestamp 1710899220
transform 1 0 2388 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2766
timestamp 1710899220
transform 1 0 2308 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2767
timestamp 1710899220
transform 1 0 2204 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2768
timestamp 1710899220
transform 1 0 2516 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_2769
timestamp 1710899220
transform 1 0 2404 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_2770
timestamp 1710899220
transform 1 0 2644 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_2771
timestamp 1710899220
transform 1 0 2596 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_2772
timestamp 1710899220
transform 1 0 2484 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_2773
timestamp 1710899220
transform 1 0 2668 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_2774
timestamp 1710899220
transform 1 0 2556 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_2775
timestamp 1710899220
transform 1 0 2444 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_2776
timestamp 1710899220
transform 1 0 2500 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_2777
timestamp 1710899220
transform 1 0 2364 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_2778
timestamp 1710899220
transform 1 0 2652 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2779
timestamp 1710899220
transform 1 0 2556 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2780
timestamp 1710899220
transform 1 0 2452 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2781
timestamp 1710899220
transform 1 0 2660 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_2782
timestamp 1710899220
transform 1 0 2548 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_2783
timestamp 1710899220
transform 1 0 2444 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_2784
timestamp 1710899220
transform 1 0 2644 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2785
timestamp 1710899220
transform 1 0 2532 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2786
timestamp 1710899220
transform 1 0 2428 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2787
timestamp 1710899220
transform 1 0 2668 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_2788
timestamp 1710899220
transform 1 0 2572 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_2789
timestamp 1710899220
transform 1 0 2468 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_2790
timestamp 1710899220
transform 1 0 2372 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2791
timestamp 1710899220
transform 1 0 2316 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2792
timestamp 1710899220
transform 1 0 2372 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2793
timestamp 1710899220
transform 1 0 2316 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2794
timestamp 1710899220
transform 1 0 2668 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2795
timestamp 1710899220
transform 1 0 2572 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2796
timestamp 1710899220
transform 1 0 2460 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2797
timestamp 1710899220
transform 1 0 2660 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2798
timestamp 1710899220
transform 1 0 2620 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2799
timestamp 1710899220
transform 1 0 2548 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2800
timestamp 1710899220
transform 1 0 2540 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2801
timestamp 1710899220
transform 1 0 2500 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2802
timestamp 1710899220
transform 1 0 2436 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2803
timestamp 1710899220
transform 1 0 2340 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2804
timestamp 1710899220
transform 1 0 2324 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2805
timestamp 1710899220
transform 1 0 2556 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2806
timestamp 1710899220
transform 1 0 2492 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2807
timestamp 1710899220
transform 1 0 2380 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2808
timestamp 1710899220
transform 1 0 2668 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2809
timestamp 1710899220
transform 1 0 2540 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2810
timestamp 1710899220
transform 1 0 2052 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2811
timestamp 1710899220
transform 1 0 1996 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2812
timestamp 1710899220
transform 1 0 2284 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2813
timestamp 1710899220
transform 1 0 2148 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2814
timestamp 1710899220
transform 1 0 2148 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2815
timestamp 1710899220
transform 1 0 2020 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2816
timestamp 1710899220
transform 1 0 2180 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2817
timestamp 1710899220
transform 1 0 2108 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2818
timestamp 1710899220
transform 1 0 1196 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_2819
timestamp 1710899220
transform 1 0 1092 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2820
timestamp 1710899220
transform 1 0 1092 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_2821
timestamp 1710899220
transform 1 0 940 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2822
timestamp 1710899220
transform 1 0 820 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2823
timestamp 1710899220
transform 1 0 812 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2824
timestamp 1710899220
transform 1 0 780 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2825
timestamp 1710899220
transform 1 0 764 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2826
timestamp 1710899220
transform 1 0 740 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2827
timestamp 1710899220
transform 1 0 740 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2828
timestamp 1710899220
transform 1 0 660 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2829
timestamp 1710899220
transform 1 0 620 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2830
timestamp 1710899220
transform 1 0 620 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2831
timestamp 1710899220
transform 1 0 604 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2832
timestamp 1710899220
transform 1 0 604 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2833
timestamp 1710899220
transform 1 0 580 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2834
timestamp 1710899220
transform 1 0 580 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2835
timestamp 1710899220
transform 1 0 572 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2836
timestamp 1710899220
transform 1 0 564 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2837
timestamp 1710899220
transform 1 0 516 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2838
timestamp 1710899220
transform 1 0 468 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2839
timestamp 1710899220
transform 1 0 356 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2840
timestamp 1710899220
transform 1 0 348 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2841
timestamp 1710899220
transform 1 0 324 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2842
timestamp 1710899220
transform 1 0 1188 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2843
timestamp 1710899220
transform 1 0 1164 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2844
timestamp 1710899220
transform 1 0 1164 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2845
timestamp 1710899220
transform 1 0 1124 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2846
timestamp 1710899220
transform 1 0 1092 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2847
timestamp 1710899220
transform 1 0 1084 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2848
timestamp 1710899220
transform 1 0 1060 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2849
timestamp 1710899220
transform 1 0 844 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2850
timestamp 1710899220
transform 1 0 828 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2851
timestamp 1710899220
transform 1 0 756 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2852
timestamp 1710899220
transform 1 0 668 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2853
timestamp 1710899220
transform 1 0 668 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2854
timestamp 1710899220
transform 1 0 636 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2855
timestamp 1710899220
transform 1 0 636 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2856
timestamp 1710899220
transform 1 0 620 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2857
timestamp 1710899220
transform 1 0 620 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2858
timestamp 1710899220
transform 1 0 604 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2859
timestamp 1710899220
transform 1 0 596 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2860
timestamp 1710899220
transform 1 0 556 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2861
timestamp 1710899220
transform 1 0 548 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2862
timestamp 1710899220
transform 1 0 484 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2863
timestamp 1710899220
transform 1 0 396 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2864
timestamp 1710899220
transform 1 0 300 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2865
timestamp 1710899220
transform 1 0 132 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2866
timestamp 1710899220
transform 1 0 132 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2867
timestamp 1710899220
transform 1 0 100 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2868
timestamp 1710899220
transform 1 0 1308 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_2869
timestamp 1710899220
transform 1 0 1252 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_2870
timestamp 1710899220
transform 1 0 1140 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_2871
timestamp 1710899220
transform 1 0 1124 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2872
timestamp 1710899220
transform 1 0 1092 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2873
timestamp 1710899220
transform 1 0 1036 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2874
timestamp 1710899220
transform 1 0 1028 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2875
timestamp 1710899220
transform 1 0 916 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2876
timestamp 1710899220
transform 1 0 916 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2877
timestamp 1710899220
transform 1 0 900 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2878
timestamp 1710899220
transform 1 0 860 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2879
timestamp 1710899220
transform 1 0 364 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2880
timestamp 1710899220
transform 1 0 324 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2881
timestamp 1710899220
transform 1 0 324 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2882
timestamp 1710899220
transform 1 0 308 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2883
timestamp 1710899220
transform 1 0 300 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2884
timestamp 1710899220
transform 1 0 300 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2885
timestamp 1710899220
transform 1 0 220 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2886
timestamp 1710899220
transform 1 0 188 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2887
timestamp 1710899220
transform 1 0 132 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2888
timestamp 1710899220
transform 1 0 108 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2889
timestamp 1710899220
transform 1 0 108 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2890
timestamp 1710899220
transform 1 0 92 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2891
timestamp 1710899220
transform 1 0 1444 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_2892
timestamp 1710899220
transform 1 0 1308 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_2893
timestamp 1710899220
transform 1 0 1308 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2894
timestamp 1710899220
transform 1 0 1220 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2895
timestamp 1710899220
transform 1 0 1180 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2896
timestamp 1710899220
transform 1 0 1180 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_2897
timestamp 1710899220
transform 1 0 1148 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2898
timestamp 1710899220
transform 1 0 1148 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2899
timestamp 1710899220
transform 1 0 1116 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2900
timestamp 1710899220
transform 1 0 1108 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_2901
timestamp 1710899220
transform 1 0 1076 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2902
timestamp 1710899220
transform 1 0 1076 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2903
timestamp 1710899220
transform 1 0 980 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2904
timestamp 1710899220
transform 1 0 956 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2905
timestamp 1710899220
transform 1 0 804 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2906
timestamp 1710899220
transform 1 0 804 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2907
timestamp 1710899220
transform 1 0 716 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2908
timestamp 1710899220
transform 1 0 668 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2909
timestamp 1710899220
transform 1 0 660 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2910
timestamp 1710899220
transform 1 0 212 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2911
timestamp 1710899220
transform 1 0 188 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2912
timestamp 1710899220
transform 1 0 132 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2913
timestamp 1710899220
transform 1 0 132 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2914
timestamp 1710899220
transform 1 0 84 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2915
timestamp 1710899220
transform 1 0 84 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2916
timestamp 1710899220
transform 1 0 84 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2917
timestamp 1710899220
transform 1 0 1292 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2918
timestamp 1710899220
transform 1 0 1188 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2919
timestamp 1710899220
transform 1 0 1076 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2920
timestamp 1710899220
transform 1 0 1044 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2921
timestamp 1710899220
transform 1 0 1012 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2922
timestamp 1710899220
transform 1 0 1012 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2923
timestamp 1710899220
transform 1 0 748 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_2924
timestamp 1710899220
transform 1 0 748 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2925
timestamp 1710899220
transform 1 0 716 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2926
timestamp 1710899220
transform 1 0 76 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_2927
timestamp 1710899220
transform 1 0 2180 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2928
timestamp 1710899220
transform 1 0 2124 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2929
timestamp 1710899220
transform 1 0 1876 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2930
timestamp 1710899220
transform 1 0 1836 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2931
timestamp 1710899220
transform 1 0 1828 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2932
timestamp 1710899220
transform 1 0 1828 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2933
timestamp 1710899220
transform 1 0 1828 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2934
timestamp 1710899220
transform 1 0 1812 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2935
timestamp 1710899220
transform 1 0 1740 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2936
timestamp 1710899220
transform 1 0 1740 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2937
timestamp 1710899220
transform 1 0 556 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_2938
timestamp 1710899220
transform 1 0 548 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2939
timestamp 1710899220
transform 1 0 508 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_2940
timestamp 1710899220
transform 1 0 500 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2941
timestamp 1710899220
transform 1 0 1852 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2942
timestamp 1710899220
transform 1 0 1788 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_2943
timestamp 1710899220
transform 1 0 1700 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2944
timestamp 1710899220
transform 1 0 1132 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2945
timestamp 1710899220
transform 1 0 1132 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_2946
timestamp 1710899220
transform 1 0 1084 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2947
timestamp 1710899220
transform 1 0 1084 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2948
timestamp 1710899220
transform 1 0 932 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2949
timestamp 1710899220
transform 1 0 916 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2950
timestamp 1710899220
transform 1 0 492 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2951
timestamp 1710899220
transform 1 0 492 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2952
timestamp 1710899220
transform 1 0 484 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2953
timestamp 1710899220
transform 1 0 452 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2954
timestamp 1710899220
transform 1 0 452 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2955
timestamp 1710899220
transform 1 0 1988 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2956
timestamp 1710899220
transform 1 0 1988 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2957
timestamp 1710899220
transform 1 0 1964 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2958
timestamp 1710899220
transform 1 0 1964 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_2959
timestamp 1710899220
transform 1 0 1940 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2960
timestamp 1710899220
transform 1 0 1908 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2961
timestamp 1710899220
transform 1 0 1900 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_2962
timestamp 1710899220
transform 1 0 1892 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_2963
timestamp 1710899220
transform 1 0 1892 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2964
timestamp 1710899220
transform 1 0 1812 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2965
timestamp 1710899220
transform 1 0 1788 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_2966
timestamp 1710899220
transform 1 0 1580 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2967
timestamp 1710899220
transform 1 0 1068 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2968
timestamp 1710899220
transform 1 0 1060 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2969
timestamp 1710899220
transform 1 0 892 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2970
timestamp 1710899220
transform 1 0 668 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2971
timestamp 1710899220
transform 1 0 428 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2972
timestamp 1710899220
transform 1 0 396 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2973
timestamp 1710899220
transform 1 0 396 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2974
timestamp 1710899220
transform 1 0 156 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2975
timestamp 1710899220
transform 1 0 156 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2976
timestamp 1710899220
transform 1 0 92 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2977
timestamp 1710899220
transform 1 0 92 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2978
timestamp 1710899220
transform 1 0 1708 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2979
timestamp 1710899220
transform 1 0 1700 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2980
timestamp 1710899220
transform 1 0 1676 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2981
timestamp 1710899220
transform 1 0 1668 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2982
timestamp 1710899220
transform 1 0 1588 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2983
timestamp 1710899220
transform 1 0 1580 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2984
timestamp 1710899220
transform 1 0 1052 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2985
timestamp 1710899220
transform 1 0 804 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2986
timestamp 1710899220
transform 1 0 804 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2987
timestamp 1710899220
transform 1 0 636 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2988
timestamp 1710899220
transform 1 0 388 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2989
timestamp 1710899220
transform 1 0 388 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2990
timestamp 1710899220
transform 1 0 348 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2991
timestamp 1710899220
transform 1 0 300 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_2992
timestamp 1710899220
transform 1 0 300 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2993
timestamp 1710899220
transform 1 0 260 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2994
timestamp 1710899220
transform 1 0 260 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2995
timestamp 1710899220
transform 1 0 68 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2996
timestamp 1710899220
transform 1 0 68 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2997
timestamp 1710899220
transform 1 0 1724 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2998
timestamp 1710899220
transform 1 0 1692 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2999
timestamp 1710899220
transform 1 0 1676 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_3000
timestamp 1710899220
transform 1 0 1596 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_3001
timestamp 1710899220
transform 1 0 1564 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3002
timestamp 1710899220
transform 1 0 1540 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_3003
timestamp 1710899220
transform 1 0 1396 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3004
timestamp 1710899220
transform 1 0 1396 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_3005
timestamp 1710899220
transform 1 0 1012 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3006
timestamp 1710899220
transform 1 0 668 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3007
timestamp 1710899220
transform 1 0 660 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3008
timestamp 1710899220
transform 1 0 660 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_3009
timestamp 1710899220
transform 1 0 628 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_3010
timestamp 1710899220
transform 1 0 612 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3011
timestamp 1710899220
transform 1 0 612 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_3012
timestamp 1710899220
transform 1 0 588 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_3013
timestamp 1710899220
transform 1 0 484 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3014
timestamp 1710899220
transform 1 0 1524 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3015
timestamp 1710899220
transform 1 0 1524 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_3016
timestamp 1710899220
transform 1 0 1492 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3017
timestamp 1710899220
transform 1 0 1468 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_3018
timestamp 1710899220
transform 1 0 700 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_3019
timestamp 1710899220
transform 1 0 636 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3020
timestamp 1710899220
transform 1 0 620 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_3021
timestamp 1710899220
transform 1 0 612 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_3022
timestamp 1710899220
transform 1 0 604 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_3023
timestamp 1710899220
transform 1 0 540 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_3024
timestamp 1710899220
transform 1 0 444 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3025
timestamp 1710899220
transform 1 0 2140 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_3026
timestamp 1710899220
transform 1 0 2140 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_3027
timestamp 1710899220
transform 1 0 1892 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_3028
timestamp 1710899220
transform 1 0 1884 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_3029
timestamp 1710899220
transform 1 0 1884 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_3030
timestamp 1710899220
transform 1 0 1860 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_3031
timestamp 1710899220
transform 1 0 1844 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_3032
timestamp 1710899220
transform 1 0 1700 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_3033
timestamp 1710899220
transform 1 0 1692 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_3034
timestamp 1710899220
transform 1 0 708 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_3035
timestamp 1710899220
transform 1 0 700 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3036
timestamp 1710899220
transform 1 0 636 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3037
timestamp 1710899220
transform 1 0 388 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_3038
timestamp 1710899220
transform 1 0 2100 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_3039
timestamp 1710899220
transform 1 0 2100 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_3040
timestamp 1710899220
transform 1 0 2100 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3041
timestamp 1710899220
transform 1 0 2092 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3042
timestamp 1710899220
transform 1 0 1932 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_3043
timestamp 1710899220
transform 1 0 1932 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3044
timestamp 1710899220
transform 1 0 1924 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_3045
timestamp 1710899220
transform 1 0 1924 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_3046
timestamp 1710899220
transform 1 0 1884 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_3047
timestamp 1710899220
transform 1 0 1876 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_3048
timestamp 1710899220
transform 1 0 684 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_3049
timestamp 1710899220
transform 1 0 684 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_3050
timestamp 1710899220
transform 1 0 660 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_3051
timestamp 1710899220
transform 1 0 628 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3052
timestamp 1710899220
transform 1 0 628 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_3053
timestamp 1710899220
transform 1 0 604 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3054
timestamp 1710899220
transform 1 0 596 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3055
timestamp 1710899220
transform 1 0 364 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_3056
timestamp 1710899220
transform 1 0 1604 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_3057
timestamp 1710899220
transform 1 0 1524 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3058
timestamp 1710899220
transform 1 0 1404 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3059
timestamp 1710899220
transform 1 0 1388 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_3060
timestamp 1710899220
transform 1 0 1388 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_3061
timestamp 1710899220
transform 1 0 996 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_3062
timestamp 1710899220
transform 1 0 996 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3063
timestamp 1710899220
transform 1 0 692 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_3064
timestamp 1710899220
transform 1 0 692 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_3065
timestamp 1710899220
transform 1 0 604 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_3066
timestamp 1710899220
transform 1 0 460 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_3067
timestamp 1710899220
transform 1 0 444 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_3068
timestamp 1710899220
transform 1 0 436 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_3069
timestamp 1710899220
transform 1 0 884 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3070
timestamp 1710899220
transform 1 0 844 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3071
timestamp 1710899220
transform 1 0 836 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3072
timestamp 1710899220
transform 1 0 716 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3073
timestamp 1710899220
transform 1 0 700 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3074
timestamp 1710899220
transform 1 0 596 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3075
timestamp 1710899220
transform 1 0 596 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_3076
timestamp 1710899220
transform 1 0 556 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_3077
timestamp 1710899220
transform 1 0 436 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_3078
timestamp 1710899220
transform 1 0 436 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_3079
timestamp 1710899220
transform 1 0 428 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3080
timestamp 1710899220
transform 1 0 404 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_3081
timestamp 1710899220
transform 1 0 404 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_3082
timestamp 1710899220
transform 1 0 1564 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_3083
timestamp 1710899220
transform 1 0 1540 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_3084
timestamp 1710899220
transform 1 0 1516 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_3085
timestamp 1710899220
transform 1 0 1476 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3086
timestamp 1710899220
transform 1 0 1364 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3087
timestamp 1710899220
transform 1 0 1204 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3088
timestamp 1710899220
transform 1 0 1188 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_3089
timestamp 1710899220
transform 1 0 900 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3090
timestamp 1710899220
transform 1 0 868 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_3091
timestamp 1710899220
transform 1 0 868 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_3092
timestamp 1710899220
transform 1 0 812 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_3093
timestamp 1710899220
transform 1 0 796 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_3094
timestamp 1710899220
transform 1 0 772 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3095
timestamp 1710899220
transform 1 0 764 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_3096
timestamp 1710899220
transform 1 0 764 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3097
timestamp 1710899220
transform 1 0 756 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_3098
timestamp 1710899220
transform 1 0 692 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3099
timestamp 1710899220
transform 1 0 692 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3100
timestamp 1710899220
transform 1 0 380 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3101
timestamp 1710899220
transform 1 0 380 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3102
timestamp 1710899220
transform 1 0 1580 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_3103
timestamp 1710899220
transform 1 0 1532 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_3104
timestamp 1710899220
transform 1 0 1356 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_3105
timestamp 1710899220
transform 1 0 1308 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_3106
timestamp 1710899220
transform 1 0 1188 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_3107
timestamp 1710899220
transform 1 0 1020 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3108
timestamp 1710899220
transform 1 0 1020 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_3109
timestamp 1710899220
transform 1 0 868 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_3110
timestamp 1710899220
transform 1 0 868 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_3111
timestamp 1710899220
transform 1 0 660 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3112
timestamp 1710899220
transform 1 0 348 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_3113
timestamp 1710899220
transform 1 0 348 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3114
timestamp 1710899220
transform 1 0 332 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3115
timestamp 1710899220
transform 1 0 332 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_3116
timestamp 1710899220
transform 1 0 68 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3117
timestamp 1710899220
transform 1 0 68 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_3118
timestamp 1710899220
transform 1 0 1092 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3119
timestamp 1710899220
transform 1 0 1060 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3120
timestamp 1710899220
transform 1 0 1020 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_3121
timestamp 1710899220
transform 1 0 1020 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_3122
timestamp 1710899220
transform 1 0 956 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_3123
timestamp 1710899220
transform 1 0 660 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_3124
timestamp 1710899220
transform 1 0 652 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_3125
timestamp 1710899220
transform 1 0 628 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_3126
timestamp 1710899220
transform 1 0 628 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_3127
timestamp 1710899220
transform 1 0 604 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_3128
timestamp 1710899220
transform 1 0 596 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_3129
timestamp 1710899220
transform 1 0 588 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3130
timestamp 1710899220
transform 1 0 588 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_3131
timestamp 1710899220
transform 1 0 564 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3132
timestamp 1710899220
transform 1 0 564 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3133
timestamp 1710899220
transform 1 0 564 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_3134
timestamp 1710899220
transform 1 0 564 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_3135
timestamp 1710899220
transform 1 0 548 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_3136
timestamp 1710899220
transform 1 0 548 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3137
timestamp 1710899220
transform 1 0 484 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_3138
timestamp 1710899220
transform 1 0 140 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_3139
timestamp 1710899220
transform 1 0 140 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3140
timestamp 1710899220
transform 1 0 140 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3141
timestamp 1710899220
transform 1 0 140 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_3142
timestamp 1710899220
transform 1 0 1228 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_3143
timestamp 1710899220
transform 1 0 1052 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_3144
timestamp 1710899220
transform 1 0 980 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_3145
timestamp 1710899220
transform 1 0 980 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_3146
timestamp 1710899220
transform 1 0 900 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_3147
timestamp 1710899220
transform 1 0 892 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_3148
timestamp 1710899220
transform 1 0 884 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3149
timestamp 1710899220
transform 1 0 868 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3150
timestamp 1710899220
transform 1 0 868 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_3151
timestamp 1710899220
transform 1 0 868 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_3152
timestamp 1710899220
transform 1 0 860 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_3153
timestamp 1710899220
transform 1 0 844 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_3154
timestamp 1710899220
transform 1 0 844 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_3155
timestamp 1710899220
transform 1 0 788 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3156
timestamp 1710899220
transform 1 0 780 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_3157
timestamp 1710899220
transform 1 0 724 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_3158
timestamp 1710899220
transform 1 0 676 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_3159
timestamp 1710899220
transform 1 0 676 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_3160
timestamp 1710899220
transform 1 0 564 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_3161
timestamp 1710899220
transform 1 0 556 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3162
timestamp 1710899220
transform 1 0 532 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3163
timestamp 1710899220
transform 1 0 516 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_3164
timestamp 1710899220
transform 1 0 492 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3165
timestamp 1710899220
transform 1 0 492 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_3166
timestamp 1710899220
transform 1 0 452 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3167
timestamp 1710899220
transform 1 0 1068 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_3168
timestamp 1710899220
transform 1 0 900 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3169
timestamp 1710899220
transform 1 0 748 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_3170
timestamp 1710899220
transform 1 0 748 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_3171
timestamp 1710899220
transform 1 0 724 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_3172
timestamp 1710899220
transform 1 0 716 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_3173
timestamp 1710899220
transform 1 0 716 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3174
timestamp 1710899220
transform 1 0 700 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3175
timestamp 1710899220
transform 1 0 620 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3176
timestamp 1710899220
transform 1 0 604 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_3177
timestamp 1710899220
transform 1 0 572 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_3178
timestamp 1710899220
transform 1 0 428 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_3179
timestamp 1710899220
transform 1 0 420 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_3180
timestamp 1710899220
transform 1 0 412 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_3181
timestamp 1710899220
transform 1 0 404 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_3182
timestamp 1710899220
transform 1 0 276 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_3183
timestamp 1710899220
transform 1 0 276 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_3184
timestamp 1710899220
transform 1 0 252 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3185
timestamp 1710899220
transform 1 0 236 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_3186
timestamp 1710899220
transform 1 0 1116 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_3187
timestamp 1710899220
transform 1 0 716 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_3188
timestamp 1710899220
transform 1 0 700 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_3189
timestamp 1710899220
transform 1 0 588 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_3190
timestamp 1710899220
transform 1 0 588 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_3191
timestamp 1710899220
transform 1 0 580 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3192
timestamp 1710899220
transform 1 0 572 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_3193
timestamp 1710899220
transform 1 0 564 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_3194
timestamp 1710899220
transform 1 0 548 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_3195
timestamp 1710899220
transform 1 0 540 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_3196
timestamp 1710899220
transform 1 0 532 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_3197
timestamp 1710899220
transform 1 0 532 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_3198
timestamp 1710899220
transform 1 0 452 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_3199
timestamp 1710899220
transform 1 0 396 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_3200
timestamp 1710899220
transform 1 0 268 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_3201
timestamp 1710899220
transform 1 0 268 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_3202
timestamp 1710899220
transform 1 0 796 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3203
timestamp 1710899220
transform 1 0 732 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_3204
timestamp 1710899220
transform 1 0 708 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_3205
timestamp 1710899220
transform 1 0 668 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3206
timestamp 1710899220
transform 1 0 484 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3207
timestamp 1710899220
transform 1 0 484 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_3208
timestamp 1710899220
transform 1 0 460 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_3209
timestamp 1710899220
transform 1 0 452 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_3210
timestamp 1710899220
transform 1 0 444 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3211
timestamp 1710899220
transform 1 0 436 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3212
timestamp 1710899220
transform 1 0 436 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_3213
timestamp 1710899220
transform 1 0 436 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3214
timestamp 1710899220
transform 1 0 436 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_3215
timestamp 1710899220
transform 1 0 396 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_3216
timestamp 1710899220
transform 1 0 396 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_3217
timestamp 1710899220
transform 1 0 316 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_3218
timestamp 1710899220
transform 1 0 316 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_3219
timestamp 1710899220
transform 1 0 316 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3220
timestamp 1710899220
transform 1 0 316 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_3221
timestamp 1710899220
transform 1 0 900 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_3222
timestamp 1710899220
transform 1 0 860 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_3223
timestamp 1710899220
transform 1 0 732 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_3224
timestamp 1710899220
transform 1 0 732 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_3225
timestamp 1710899220
transform 1 0 636 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_3226
timestamp 1710899220
transform 1 0 532 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_3227
timestamp 1710899220
transform 1 0 500 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_3228
timestamp 1710899220
transform 1 0 484 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_3229
timestamp 1710899220
transform 1 0 412 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_3230
timestamp 1710899220
transform 1 0 404 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_3231
timestamp 1710899220
transform 1 0 404 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_3232
timestamp 1710899220
transform 1 0 268 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3233
timestamp 1710899220
transform 1 0 268 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_3234
timestamp 1710899220
transform 1 0 196 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_3235
timestamp 1710899220
transform 1 0 196 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_3236
timestamp 1710899220
transform 1 0 164 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_3237
timestamp 1710899220
transform 1 0 164 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3238
timestamp 1710899220
transform 1 0 124 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_3239
timestamp 1710899220
transform 1 0 124 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_3240
timestamp 1710899220
transform 1 0 996 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_3241
timestamp 1710899220
transform 1 0 980 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_3242
timestamp 1710899220
transform 1 0 980 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3243
timestamp 1710899220
transform 1 0 924 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_3244
timestamp 1710899220
transform 1 0 924 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_3245
timestamp 1710899220
transform 1 0 916 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3246
timestamp 1710899220
transform 1 0 868 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_3247
timestamp 1710899220
transform 1 0 868 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_3248
timestamp 1710899220
transform 1 0 868 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_3249
timestamp 1710899220
transform 1 0 820 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_3250
timestamp 1710899220
transform 1 0 724 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_3251
timestamp 1710899220
transform 1 0 404 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_3252
timestamp 1710899220
transform 1 0 356 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_3253
timestamp 1710899220
transform 1 0 348 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_3254
timestamp 1710899220
transform 1 0 1012 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3255
timestamp 1710899220
transform 1 0 964 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3256
timestamp 1710899220
transform 1 0 924 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_3257
timestamp 1710899220
transform 1 0 924 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3258
timestamp 1710899220
transform 1 0 916 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3259
timestamp 1710899220
transform 1 0 892 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3260
timestamp 1710899220
transform 1 0 828 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3261
timestamp 1710899220
transform 1 0 676 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3262
timestamp 1710899220
transform 1 0 676 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_3263
timestamp 1710899220
transform 1 0 668 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_3264
timestamp 1710899220
transform 1 0 340 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_3265
timestamp 1710899220
transform 1 0 324 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3266
timestamp 1710899220
transform 1 0 316 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3267
timestamp 1710899220
transform 1 0 1068 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3268
timestamp 1710899220
transform 1 0 1036 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3269
timestamp 1710899220
transform 1 0 1036 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_3270
timestamp 1710899220
transform 1 0 972 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_3271
timestamp 1710899220
transform 1 0 956 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3272
timestamp 1710899220
transform 1 0 948 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_3273
timestamp 1710899220
transform 1 0 692 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3274
timestamp 1710899220
transform 1 0 692 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_3275
timestamp 1710899220
transform 1 0 548 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_3276
timestamp 1710899220
transform 1 0 540 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_3277
timestamp 1710899220
transform 1 0 540 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3278
timestamp 1710899220
transform 1 0 524 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_3279
timestamp 1710899220
transform 1 0 484 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_3280
timestamp 1710899220
transform 1 0 476 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3281
timestamp 1710899220
transform 1 0 556 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_3282
timestamp 1710899220
transform 1 0 548 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3283
timestamp 1710899220
transform 1 0 508 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_3284
timestamp 1710899220
transform 1 0 484 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_3285
timestamp 1710899220
transform 1 0 484 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_3286
timestamp 1710899220
transform 1 0 476 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3287
timestamp 1710899220
transform 1 0 460 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_3288
timestamp 1710899220
transform 1 0 452 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_3289
timestamp 1710899220
transform 1 0 444 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3290
timestamp 1710899220
transform 1 0 428 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_3291
timestamp 1710899220
transform 1 0 428 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3292
timestamp 1710899220
transform 1 0 900 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_3293
timestamp 1710899220
transform 1 0 676 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_3294
timestamp 1710899220
transform 1 0 580 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_3295
timestamp 1710899220
transform 1 0 492 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3296
timestamp 1710899220
transform 1 0 460 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_3297
timestamp 1710899220
transform 1 0 436 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_3298
timestamp 1710899220
transform 1 0 436 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3299
timestamp 1710899220
transform 1 0 428 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3300
timestamp 1710899220
transform 1 0 428 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_3301
timestamp 1710899220
transform 1 0 420 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_3302
timestamp 1710899220
transform 1 0 412 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_3303
timestamp 1710899220
transform 1 0 412 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_3304
timestamp 1710899220
transform 1 0 404 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_3305
timestamp 1710899220
transform 1 0 404 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3306
timestamp 1710899220
transform 1 0 388 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3307
timestamp 1710899220
transform 1 0 388 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3308
timestamp 1710899220
transform 1 0 380 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_3309
timestamp 1710899220
transform 1 0 380 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_3310
timestamp 1710899220
transform 1 0 364 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3311
timestamp 1710899220
transform 1 0 620 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_3312
timestamp 1710899220
transform 1 0 556 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3313
timestamp 1710899220
transform 1 0 556 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_3314
timestamp 1710899220
transform 1 0 548 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_3315
timestamp 1710899220
transform 1 0 548 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_3316
timestamp 1710899220
transform 1 0 492 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3317
timestamp 1710899220
transform 1 0 492 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_3318
timestamp 1710899220
transform 1 0 484 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_3319
timestamp 1710899220
transform 1 0 452 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_3320
timestamp 1710899220
transform 1 0 412 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3321
timestamp 1710899220
transform 1 0 364 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3322
timestamp 1710899220
transform 1 0 364 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3323
timestamp 1710899220
transform 1 0 276 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_3324
timestamp 1710899220
transform 1 0 276 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3325
timestamp 1710899220
transform 1 0 156 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_3326
timestamp 1710899220
transform 1 0 140 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3327
timestamp 1710899220
transform 1 0 108 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_3328
timestamp 1710899220
transform 1 0 108 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_3329
timestamp 1710899220
transform 1 0 940 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_3330
timestamp 1710899220
transform 1 0 932 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3331
timestamp 1710899220
transform 1 0 924 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_3332
timestamp 1710899220
transform 1 0 924 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_3333
timestamp 1710899220
transform 1 0 916 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3334
timestamp 1710899220
transform 1 0 916 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_3335
timestamp 1710899220
transform 1 0 892 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_3336
timestamp 1710899220
transform 1 0 884 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_3337
timestamp 1710899220
transform 1 0 852 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3338
timestamp 1710899220
transform 1 0 820 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_3339
timestamp 1710899220
transform 1 0 764 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_3340
timestamp 1710899220
transform 1 0 588 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_3341
timestamp 1710899220
transform 1 0 2420 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3342
timestamp 1710899220
transform 1 0 2268 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3343
timestamp 1710899220
transform 1 0 2252 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_3344
timestamp 1710899220
transform 1 0 2244 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3345
timestamp 1710899220
transform 1 0 2228 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_3346
timestamp 1710899220
transform 1 0 2164 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_3347
timestamp 1710899220
transform 1 0 2108 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3348
timestamp 1710899220
transform 1 0 2460 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3349
timestamp 1710899220
transform 1 0 2420 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3350
timestamp 1710899220
transform 1 0 2660 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3351
timestamp 1710899220
transform 1 0 2620 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3352
timestamp 1710899220
transform 1 0 2668 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_3353
timestamp 1710899220
transform 1 0 2652 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3354
timestamp 1710899220
transform 1 0 2644 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_3355
timestamp 1710899220
transform 1 0 2620 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3356
timestamp 1710899220
transform 1 0 2612 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_3357
timestamp 1710899220
transform 1 0 2596 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3358
timestamp 1710899220
transform 1 0 2596 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_3359
timestamp 1710899220
transform 1 0 2564 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3360
timestamp 1710899220
transform 1 0 2564 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3361
timestamp 1710899220
transform 1 0 2636 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3362
timestamp 1710899220
transform 1 0 2596 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3363
timestamp 1710899220
transform 1 0 2564 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3364
timestamp 1710899220
transform 1 0 2500 0 1 795
box -3 -3 3 3
use MUX2X1  MUX2X1_0
timestamp 1710899220
transform 1 0 168 0 -1 2570
box -5 -3 53 105
use MUX2X1  MUX2X1_1
timestamp 1710899220
transform 1 0 184 0 1 2370
box -5 -3 53 105
use MUX2X1  MUX2X1_2
timestamp 1710899220
transform 1 0 232 0 -1 2370
box -5 -3 53 105
use MUX2X1  MUX2X1_3
timestamp 1710899220
transform 1 0 320 0 1 2370
box -5 -3 53 105
use MUX2X1  MUX2X1_4
timestamp 1710899220
transform 1 0 376 0 -1 2370
box -5 -3 53 105
use MUX2X1  MUX2X1_5
timestamp 1710899220
transform 1 0 344 0 -1 2570
box -5 -3 53 105
use MUX2X1  MUX2X1_6
timestamp 1710899220
transform 1 0 472 0 -1 2570
box -5 -3 53 105
use MUX2X1  MUX2X1_7
timestamp 1710899220
transform 1 0 528 0 1 2370
box -5 -3 53 105
use MUX2X1  MUX2X1_8
timestamp 1710899220
transform 1 0 592 0 1 2370
box -5 -3 53 105
use MUX2X1  MUX2X1_9
timestamp 1710899220
transform 1 0 648 0 -1 2370
box -5 -3 53 105
use MUX2X1  MUX2X1_10
timestamp 1710899220
transform 1 0 648 0 -1 2570
box -5 -3 53 105
use MUX2X1  MUX2X1_11
timestamp 1710899220
transform 1 0 776 0 -1 2570
box -5 -3 53 105
use MUX2X1  MUX2X1_12
timestamp 1710899220
transform 1 0 784 0 1 2370
box -5 -3 53 105
use MUX2X1  MUX2X1_13
timestamp 1710899220
transform 1 0 896 0 1 2370
box -5 -3 53 105
use MUX2X1  MUX2X1_14
timestamp 1710899220
transform 1 0 944 0 1 2370
box -5 -3 53 105
use MUX2X1  MUX2X1_15
timestamp 1710899220
transform 1 0 968 0 -1 2570
box -5 -3 53 105
use MUX2X1  MUX2X1_16
timestamp 1710899220
transform 1 0 1096 0 -1 2570
box -5 -3 53 105
use MUX2X1  MUX2X1_17
timestamp 1710899220
transform 1 0 1240 0 -1 2570
box -5 -3 53 105
use MUX2X1  MUX2X1_18
timestamp 1710899220
transform 1 0 1152 0 1 2370
box -5 -3 53 105
use MUX2X1  MUX2X1_19
timestamp 1710899220
transform 1 0 1208 0 1 2370
box -5 -3 53 105
use MUX2X1  MUX2X1_20
timestamp 1710899220
transform 1 0 1448 0 -1 2570
box -5 -3 53 105
use MUX2X1  MUX2X1_21
timestamp 1710899220
transform 1 0 1576 0 -1 2570
box -5 -3 53 105
use MUX2X1  MUX2X1_22
timestamp 1710899220
transform 1 0 1488 0 1 2370
box -5 -3 53 105
use MUX2X1  MUX2X1_23
timestamp 1710899220
transform 1 0 1336 0 -1 2370
box -5 -3 53 105
use MUX2X1  MUX2X1_24
timestamp 1710899220
transform 1 0 1392 0 -1 2370
box -5 -3 53 105
use MUX2X1  MUX2X1_25
timestamp 1710899220
transform 1 0 1768 0 -1 2570
box -5 -3 53 105
use MUX2X1  MUX2X1_26
timestamp 1710899220
transform 1 0 1680 0 1 2370
box -5 -3 53 105
use MUX2X1  MUX2X1_27
timestamp 1710899220
transform 1 0 1592 0 -1 2370
box -5 -3 53 105
use MUX2X1  MUX2X1_28
timestamp 1710899220
transform 1 0 1568 0 1 2170
box -5 -3 53 105
use MUX2X1  MUX2X1_29
timestamp 1710899220
transform 1 0 1464 0 1 2170
box -5 -3 53 105
use MUX2X1  MUX2X1_30
timestamp 1710899220
transform 1 0 1656 0 -1 2370
box -5 -3 53 105
use MUX2X1  MUX2X1_31
timestamp 1710899220
transform 1 0 1648 0 1 2170
box -5 -3 53 105
use MUX2X1  MUX2X1_32
timestamp 1710899220
transform 1 0 1600 0 -1 2170
box -5 -3 53 105
use MUX2X1  MUX2X1_33
timestamp 1710899220
transform 1 0 1520 0 -1 2170
box -5 -3 53 105
use MUX2X1  MUX2X1_34
timestamp 1710899220
transform 1 0 1384 0 -1 2170
box -5 -3 53 105
use NAND2X1  NAND2X1_0
timestamp 1710899220
transform 1 0 1728 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_1
timestamp 1710899220
transform 1 0 1544 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_2
timestamp 1710899220
transform 1 0 1424 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_3
timestamp 1710899220
transform 1 0 1144 0 -1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_4
timestamp 1710899220
transform 1 0 680 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_5
timestamp 1710899220
transform 1 0 400 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_6
timestamp 1710899220
transform 1 0 120 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_7
timestamp 1710899220
transform 1 0 128 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_8
timestamp 1710899220
transform 1 0 624 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_9
timestamp 1710899220
transform 1 0 712 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_10
timestamp 1710899220
transform 1 0 664 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_11
timestamp 1710899220
transform 1 0 1072 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_12
timestamp 1710899220
transform 1 0 1080 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_13
timestamp 1710899220
transform 1 0 128 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_14
timestamp 1710899220
transform 1 0 2280 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_15
timestamp 1710899220
transform 1 0 928 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_16
timestamp 1710899220
transform 1 0 640 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_17
timestamp 1710899220
transform 1 0 904 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_18
timestamp 1710899220
transform 1 0 600 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_19
timestamp 1710899220
transform 1 0 1064 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_20
timestamp 1710899220
transform 1 0 1008 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_21
timestamp 1710899220
transform 1 0 1280 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_22
timestamp 1710899220
transform 1 0 968 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_23
timestamp 1710899220
transform 1 0 1304 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_24
timestamp 1710899220
transform 1 0 896 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_25
timestamp 1710899220
transform 1 0 792 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_26
timestamp 1710899220
transform 1 0 1128 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_27
timestamp 1710899220
transform 1 0 1080 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_28
timestamp 1710899220
transform 1 0 1232 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_29
timestamp 1710899220
transform 1 0 1104 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_30
timestamp 1710899220
transform 1 0 1352 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_31
timestamp 1710899220
transform 1 0 1296 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_32
timestamp 1710899220
transform 1 0 1360 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_33
timestamp 1710899220
transform 1 0 1320 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_34
timestamp 1710899220
transform 1 0 872 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_35
timestamp 1710899220
transform 1 0 1400 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_36
timestamp 1710899220
transform 1 0 1880 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_37
timestamp 1710899220
transform 1 0 1696 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_38
timestamp 1710899220
transform 1 0 1616 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_39
timestamp 1710899220
transform 1 0 1488 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_40
timestamp 1710899220
transform 1 0 1560 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_41
timestamp 1710899220
transform 1 0 1568 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_42
timestamp 1710899220
transform 1 0 1624 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_43
timestamp 1710899220
transform 1 0 1480 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_44
timestamp 1710899220
transform 1 0 1808 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_45
timestamp 1710899220
transform 1 0 1504 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_46
timestamp 1710899220
transform 1 0 1696 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_47
timestamp 1710899220
transform 1 0 1728 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_48
timestamp 1710899220
transform 1 0 1312 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_49
timestamp 1710899220
transform 1 0 1320 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_50
timestamp 1710899220
transform 1 0 1520 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_51
timestamp 1710899220
transform 1 0 1400 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_52
timestamp 1710899220
transform 1 0 2096 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_53
timestamp 1710899220
transform 1 0 2152 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_54
timestamp 1710899220
transform 1 0 2192 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_55
timestamp 1710899220
transform 1 0 2216 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_56
timestamp 1710899220
transform 1 0 2144 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_57
timestamp 1710899220
transform 1 0 1832 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_58
timestamp 1710899220
transform 1 0 1752 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_59
timestamp 1710899220
transform 1 0 1808 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_60
timestamp 1710899220
transform 1 0 1800 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_61
timestamp 1710899220
transform 1 0 1488 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_62
timestamp 1710899220
transform 1 0 1992 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_63
timestamp 1710899220
transform 1 0 584 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_64
timestamp 1710899220
transform 1 0 1952 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_65
timestamp 1710899220
transform 1 0 1928 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_66
timestamp 1710899220
transform 1 0 376 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_67
timestamp 1710899220
transform 1 0 352 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_68
timestamp 1710899220
transform 1 0 1784 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_69
timestamp 1710899220
transform 1 0 1304 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_70
timestamp 1710899220
transform 1 0 1376 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_71
timestamp 1710899220
transform 1 0 1400 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_72
timestamp 1710899220
transform 1 0 1368 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_73
timestamp 1710899220
transform 1 0 1344 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_74
timestamp 1710899220
transform 1 0 1344 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_75
timestamp 1710899220
transform 1 0 1408 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_76
timestamp 1710899220
transform 1 0 1432 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_77
timestamp 1710899220
transform 1 0 1456 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_78
timestamp 1710899220
transform 1 0 1384 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_79
timestamp 1710899220
transform 1 0 1432 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_80
timestamp 1710899220
transform 1 0 1408 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_81
timestamp 1710899220
transform 1 0 1264 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_82
timestamp 1710899220
transform 1 0 1192 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_83
timestamp 1710899220
transform 1 0 808 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_84
timestamp 1710899220
transform 1 0 736 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_85
timestamp 1710899220
transform 1 0 664 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_86
timestamp 1710899220
transform 1 0 640 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_87
timestamp 1710899220
transform 1 0 856 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_88
timestamp 1710899220
transform 1 0 984 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_89
timestamp 1710899220
transform 1 0 1104 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_90
timestamp 1710899220
transform 1 0 680 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_91
timestamp 1710899220
transform 1 0 656 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_92
timestamp 1710899220
transform 1 0 704 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_93
timestamp 1710899220
transform 1 0 696 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_94
timestamp 1710899220
transform 1 0 1728 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_95
timestamp 1710899220
transform 1 0 2104 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_96
timestamp 1710899220
transform 1 0 1176 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_97
timestamp 1710899220
transform 1 0 1176 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_98
timestamp 1710899220
transform 1 0 1352 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_99
timestamp 1710899220
transform 1 0 1480 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_100
timestamp 1710899220
transform 1 0 1328 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_101
timestamp 1710899220
transform 1 0 1536 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_102
timestamp 1710899220
transform 1 0 784 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_103
timestamp 1710899220
transform 1 0 760 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_104
timestamp 1710899220
transform 1 0 1000 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_105
timestamp 1710899220
transform 1 0 968 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_106
timestamp 1710899220
transform 1 0 1096 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_107
timestamp 1710899220
transform 1 0 1120 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_108
timestamp 1710899220
transform 1 0 1072 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_109
timestamp 1710899220
transform 1 0 760 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_110
timestamp 1710899220
transform 1 0 600 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_111
timestamp 1710899220
transform 1 0 576 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_112
timestamp 1710899220
transform 1 0 528 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_113
timestamp 1710899220
transform 1 0 504 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_114
timestamp 1710899220
transform 1 0 272 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_115
timestamp 1710899220
transform 1 0 576 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_116
timestamp 1710899220
transform 1 0 552 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_117
timestamp 1710899220
transform 1 0 640 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_118
timestamp 1710899220
transform 1 0 616 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_119
timestamp 1710899220
transform 1 0 184 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_120
timestamp 1710899220
transform 1 0 336 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_121
timestamp 1710899220
transform 1 0 416 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_122
timestamp 1710899220
transform 1 0 464 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_123
timestamp 1710899220
transform 1 0 440 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_124
timestamp 1710899220
transform 1 0 200 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_125
timestamp 1710899220
transform 1 0 664 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_126
timestamp 1710899220
transform 1 0 624 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_127
timestamp 1710899220
transform 1 0 600 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_128
timestamp 1710899220
transform 1 0 576 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_129
timestamp 1710899220
transform 1 0 2184 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_130
timestamp 1710899220
transform 1 0 2312 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_131
timestamp 1710899220
transform 1 0 2512 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_132
timestamp 1710899220
transform 1 0 2376 0 1 170
box -8 -3 32 105
use NAND3X1  NAND3X1_0
timestamp 1710899220
transform 1 0 1256 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_1
timestamp 1710899220
transform 1 0 1032 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_2
timestamp 1710899220
transform 1 0 1000 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_3
timestamp 1710899220
transform 1 0 1216 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_4
timestamp 1710899220
transform 1 0 1288 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_5
timestamp 1710899220
transform 1 0 1320 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_6
timestamp 1710899220
transform 1 0 2248 0 -1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_7
timestamp 1710899220
transform 1 0 1640 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_8
timestamp 1710899220
transform 1 0 1528 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_9
timestamp 1710899220
transform 1 0 1536 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_10
timestamp 1710899220
transform 1 0 2136 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_11
timestamp 1710899220
transform 1 0 2208 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_12
timestamp 1710899220
transform 1 0 2048 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_13
timestamp 1710899220
transform 1 0 2256 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_14
timestamp 1710899220
transform 1 0 2224 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_15
timestamp 1710899220
transform 1 0 1512 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_16
timestamp 1710899220
transform 1 0 1504 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_17
timestamp 1710899220
transform 1 0 1376 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_18
timestamp 1710899220
transform 1 0 1416 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_19
timestamp 1710899220
transform 1 0 1032 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_20
timestamp 1710899220
transform 1 0 1760 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_21
timestamp 1710899220
transform 1 0 544 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_22
timestamp 1710899220
transform 1 0 1784 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_23
timestamp 1710899220
transform 1 0 1264 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_24
timestamp 1710899220
transform 1 0 832 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_25
timestamp 1710899220
transform 1 0 1672 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_26
timestamp 1710899220
transform 1 0 1608 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_27
timestamp 1710899220
transform 1 0 1656 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_28
timestamp 1710899220
transform 1 0 1760 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_29
timestamp 1710899220
transform 1 0 1704 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_30
timestamp 1710899220
transform 1 0 1640 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_31
timestamp 1710899220
transform 1 0 1952 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_32
timestamp 1710899220
transform 1 0 2000 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_33
timestamp 1710899220
transform 1 0 1712 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_34
timestamp 1710899220
transform 1 0 1680 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_35
timestamp 1710899220
transform 1 0 1624 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_36
timestamp 1710899220
transform 1 0 1648 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_37
timestamp 1710899220
transform 1 0 1848 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_38
timestamp 1710899220
transform 1 0 1920 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_39
timestamp 1710899220
transform 1 0 856 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_40
timestamp 1710899220
transform 1 0 328 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_41
timestamp 1710899220
transform 1 0 496 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_42
timestamp 1710899220
transform 1 0 544 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_43
timestamp 1710899220
transform 1 0 384 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_44
timestamp 1710899220
transform 1 0 1024 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_45
timestamp 1710899220
transform 1 0 1712 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_46
timestamp 1710899220
transform 1 0 608 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_47
timestamp 1710899220
transform 1 0 744 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_48
timestamp 1710899220
transform 1 0 2128 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_49
timestamp 1710899220
transform 1 0 2496 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_50
timestamp 1710899220
transform 1 0 2240 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_51
timestamp 1710899220
transform 1 0 2464 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_52
timestamp 1710899220
transform 1 0 2352 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_53
timestamp 1710899220
transform 1 0 2408 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_54
timestamp 1710899220
transform 1 0 2408 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_55
timestamp 1710899220
transform 1 0 2504 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_56
timestamp 1710899220
transform 1 0 2264 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_57
timestamp 1710899220
transform 1 0 2440 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_58
timestamp 1710899220
transform 1 0 2608 0 1 770
box -8 -3 40 105
use NOR2X1  NOR2X1_0
timestamp 1710899220
transform 1 0 1568 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_1
timestamp 1710899220
transform 1 0 1440 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_2
timestamp 1710899220
transform 1 0 1328 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_3
timestamp 1710899220
transform 1 0 1056 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_4
timestamp 1710899220
transform 1 0 856 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_5
timestamp 1710899220
transform 1 0 480 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_6
timestamp 1710899220
transform 1 0 288 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_7
timestamp 1710899220
transform 1 0 144 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_8
timestamp 1710899220
transform 1 0 1248 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_9
timestamp 1710899220
transform 1 0 1160 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_10
timestamp 1710899220
transform 1 0 1032 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_11
timestamp 1710899220
transform 1 0 960 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_12
timestamp 1710899220
transform 1 0 904 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_13
timestamp 1710899220
transform 1 0 1208 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_14
timestamp 1710899220
transform 1 0 1136 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_15
timestamp 1710899220
transform 1 0 984 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_16
timestamp 1710899220
transform 1 0 856 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_17
timestamp 1710899220
transform 1 0 880 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_18
timestamp 1710899220
transform 1 0 1072 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_19
timestamp 1710899220
transform 1 0 680 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_20
timestamp 1710899220
transform 1 0 832 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_21
timestamp 1710899220
transform 1 0 648 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_22
timestamp 1710899220
transform 1 0 480 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_23
timestamp 1710899220
transform 1 0 704 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_24
timestamp 1710899220
transform 1 0 696 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_25
timestamp 1710899220
transform 1 0 504 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_26
timestamp 1710899220
transform 1 0 424 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_27
timestamp 1710899220
transform 1 0 272 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_28
timestamp 1710899220
transform 1 0 720 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_29
timestamp 1710899220
transform 1 0 672 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_30
timestamp 1710899220
transform 1 0 456 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_31
timestamp 1710899220
transform 1 0 248 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_32
timestamp 1710899220
transform 1 0 232 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_33
timestamp 1710899220
transform 1 0 712 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_34
timestamp 1710899220
transform 1 0 544 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_35
timestamp 1710899220
transform 1 0 1336 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_36
timestamp 1710899220
transform 1 0 1288 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_37
timestamp 1710899220
transform 1 0 1320 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_38
timestamp 1710899220
transform 1 0 1344 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_39
timestamp 1710899220
transform 1 0 1320 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_40
timestamp 1710899220
transform 1 0 1272 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_41
timestamp 1710899220
transform 1 0 1320 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_42
timestamp 1710899220
transform 1 0 1352 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_43
timestamp 1710899220
transform 1 0 688 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_44
timestamp 1710899220
transform 1 0 760 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_45
timestamp 1710899220
transform 1 0 784 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_46
timestamp 1710899220
transform 1 0 736 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_47
timestamp 1710899220
transform 1 0 1080 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_48
timestamp 1710899220
transform 1 0 1328 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_49
timestamp 1710899220
transform 1 0 960 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_50
timestamp 1710899220
transform 1 0 880 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_51
timestamp 1710899220
transform 1 0 712 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_52
timestamp 1710899220
transform 1 0 688 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_53
timestamp 1710899220
transform 1 0 760 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_54
timestamp 1710899220
transform 1 0 784 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_55
timestamp 1710899220
transform 1 0 1216 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_56
timestamp 1710899220
transform 1 0 1240 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_57
timestamp 1710899220
transform 1 0 1312 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_58
timestamp 1710899220
transform 1 0 1360 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_59
timestamp 1710899220
transform 1 0 1280 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_60
timestamp 1710899220
transform 1 0 736 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_61
timestamp 1710899220
transform 1 0 1392 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_62
timestamp 1710899220
transform 1 0 1416 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_63
timestamp 1710899220
transform 1 0 1496 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_64
timestamp 1710899220
transform 1 0 1472 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_65
timestamp 1710899220
transform 1 0 1512 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_66
timestamp 1710899220
transform 1 0 1576 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_67
timestamp 1710899220
transform 1 0 1912 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_68
timestamp 1710899220
transform 1 0 2232 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_69
timestamp 1710899220
transform 1 0 2240 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_70
timestamp 1710899220
transform 1 0 2264 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_71
timestamp 1710899220
transform 1 0 1464 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_72
timestamp 1710899220
transform 1 0 1712 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_73
timestamp 1710899220
transform 1 0 1368 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_74
timestamp 1710899220
transform 1 0 1368 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_75
timestamp 1710899220
transform 1 0 1392 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_76
timestamp 1710899220
transform 1 0 1064 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_77
timestamp 1710899220
transform 1 0 1232 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_78
timestamp 1710899220
transform 1 0 1240 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_79
timestamp 1710899220
transform 1 0 1704 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_80
timestamp 1710899220
transform 1 0 1648 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_81
timestamp 1710899220
transform 1 0 1608 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_82
timestamp 1710899220
transform 1 0 1688 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_83
timestamp 1710899220
transform 1 0 1736 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_84
timestamp 1710899220
transform 1 0 1568 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_85
timestamp 1710899220
transform 1 0 1904 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_86
timestamp 1710899220
transform 1 0 1792 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_87
timestamp 1710899220
transform 1 0 1712 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_88
timestamp 1710899220
transform 1 0 1592 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_89
timestamp 1710899220
transform 1 0 1712 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_90
timestamp 1710899220
transform 1 0 1880 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_91
timestamp 1710899220
transform 1 0 832 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_92
timestamp 1710899220
transform 1 0 488 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_93
timestamp 1710899220
transform 1 0 936 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_94
timestamp 1710899220
transform 1 0 424 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_95
timestamp 1710899220
transform 1 0 1048 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_96
timestamp 1710899220
transform 1 0 1024 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_97
timestamp 1710899220
transform 1 0 1056 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_98
timestamp 1710899220
transform 1 0 1568 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_99
timestamp 1710899220
transform 1 0 1096 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_100
timestamp 1710899220
transform 1 0 904 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_101
timestamp 1710899220
transform 1 0 640 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_102
timestamp 1710899220
transform 1 0 1848 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_103
timestamp 1710899220
transform 1 0 1824 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_104
timestamp 1710899220
transform 1 0 1256 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_105
timestamp 1710899220
transform 1 0 2112 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_106
timestamp 1710899220
transform 1 0 1952 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_107
timestamp 1710899220
transform 1 0 2152 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_108
timestamp 1710899220
transform 1 0 1008 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_109
timestamp 1710899220
transform 1 0 808 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_110
timestamp 1710899220
transform 1 0 1048 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_111
timestamp 1710899220
transform 1 0 824 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_112
timestamp 1710899220
transform 1 0 808 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_113
timestamp 1710899220
transform 1 0 904 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_114
timestamp 1710899220
transform 1 0 800 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_115
timestamp 1710899220
transform 1 0 2368 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_116
timestamp 1710899220
transform 1 0 2432 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_117
timestamp 1710899220
transform 1 0 2560 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_118
timestamp 1710899220
transform 1 0 2400 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_119
timestamp 1710899220
transform 1 0 2360 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_120
timestamp 1710899220
transform 1 0 2640 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_121
timestamp 1710899220
transform 1 0 2600 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_122
timestamp 1710899220
transform 1 0 2584 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_123
timestamp 1710899220
transform 1 0 2264 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_124
timestamp 1710899220
transform 1 0 2352 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_125
timestamp 1710899220
transform 1 0 2496 0 -1 370
box -8 -3 32 105
use OAI21X1  OAI21X1_0
timestamp 1710899220
transform 1 0 592 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_1
timestamp 1710899220
transform 1 0 1120 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_2
timestamp 1710899220
transform 1 0 1088 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_3
timestamp 1710899220
transform 1 0 952 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_4
timestamp 1710899220
transform 1 0 1328 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_5
timestamp 1710899220
transform 1 0 664 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_6
timestamp 1710899220
transform 1 0 1064 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_7
timestamp 1710899220
transform 1 0 928 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_8
timestamp 1710899220
transform 1 0 1120 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_9
timestamp 1710899220
transform 1 0 624 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_10
timestamp 1710899220
transform 1 0 1096 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_11
timestamp 1710899220
transform 1 0 1032 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_12
timestamp 1710899220
transform 1 0 1128 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_13
timestamp 1710899220
transform 1 0 976 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_14
timestamp 1710899220
transform 1 0 1160 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_15
timestamp 1710899220
transform 1 0 992 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_16
timestamp 1710899220
transform 1 0 1152 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_17
timestamp 1710899220
transform 1 0 864 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_18
timestamp 1710899220
transform 1 0 1200 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_19
timestamp 1710899220
transform 1 0 816 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_20
timestamp 1710899220
transform 1 0 1232 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_21
timestamp 1710899220
transform 1 0 1152 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_22
timestamp 1710899220
transform 1 0 1224 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_23
timestamp 1710899220
transform 1 0 1104 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_24
timestamp 1710899220
transform 1 0 1192 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_25
timestamp 1710899220
transform 1 0 1256 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_26
timestamp 1710899220
transform 1 0 1256 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_27
timestamp 1710899220
transform 1 0 1128 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_28
timestamp 1710899220
transform 1 0 1216 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_29
timestamp 1710899220
transform 1 0 1320 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_30
timestamp 1710899220
transform 1 0 1288 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_31
timestamp 1710899220
transform 1 0 1328 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_32
timestamp 1710899220
transform 1 0 1320 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_33
timestamp 1710899220
transform 1 0 840 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_34
timestamp 1710899220
transform 1 0 1256 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_35
timestamp 1710899220
transform 1 0 1368 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_36
timestamp 1710899220
transform 1 0 1376 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_37
timestamp 1710899220
transform 1 0 1848 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_38
timestamp 1710899220
transform 1 0 1656 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_39
timestamp 1710899220
transform 1 0 1720 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_40
timestamp 1710899220
transform 1 0 1688 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_41
timestamp 1710899220
transform 1 0 1512 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_42
timestamp 1710899220
transform 1 0 1528 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_43
timestamp 1710899220
transform 1 0 1584 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_44
timestamp 1710899220
transform 1 0 1560 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_45
timestamp 1710899220
transform 1 0 1592 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_46
timestamp 1710899220
transform 1 0 1640 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_47
timestamp 1710899220
transform 1 0 1832 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_48
timestamp 1710899220
transform 1 0 1720 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_49
timestamp 1710899220
transform 1 0 1720 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_50
timestamp 1710899220
transform 1 0 1584 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_51
timestamp 1710899220
transform 1 0 1752 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_52
timestamp 1710899220
transform 1 0 1552 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_53
timestamp 1710899220
transform 1 0 1336 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_54
timestamp 1710899220
transform 1 0 1344 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_55
timestamp 1710899220
transform 1 0 1544 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_56
timestamp 1710899220
transform 1 0 1424 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_57
timestamp 1710899220
transform 1 0 2120 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_58
timestamp 1710899220
transform 1 0 2160 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_59
timestamp 1710899220
transform 1 0 2184 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_60
timestamp 1710899220
transform 1 0 1800 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_61
timestamp 1710899220
transform 1 0 1680 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_62
timestamp 1710899220
transform 1 0 1776 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_63
timestamp 1710899220
transform 1 0 1736 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_64
timestamp 1710899220
transform 1 0 1928 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_65
timestamp 1710899220
transform 1 0 1960 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_66
timestamp 1710899220
transform 1 0 1840 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_67
timestamp 1710899220
transform 1 0 1472 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_68
timestamp 1710899220
transform 1 0 1008 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_69
timestamp 1710899220
transform 1 0 744 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_70
timestamp 1710899220
transform 1 0 1632 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_71
timestamp 1710899220
transform 1 0 1968 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_72
timestamp 1710899220
transform 1 0 1928 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_73
timestamp 1710899220
transform 1 0 1040 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_74
timestamp 1710899220
transform 1 0 1616 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_75
timestamp 1710899220
transform 1 0 1680 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_76
timestamp 1710899220
transform 1 0 1904 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_77
timestamp 1710899220
transform 1 0 360 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_78
timestamp 1710899220
transform 1 0 416 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_79
timestamp 1710899220
transform 1 0 392 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_80
timestamp 1710899220
transform 1 0 1680 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_81
timestamp 1710899220
transform 1 0 736 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_82
timestamp 1710899220
transform 1 0 1424 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_83
timestamp 1710899220
transform 1 0 1792 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_84
timestamp 1710899220
transform 1 0 1752 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_85
timestamp 1710899220
transform 1 0 1520 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_86
timestamp 1710899220
transform 1 0 1392 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_87
timestamp 1710899220
transform 1 0 1392 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_88
timestamp 1710899220
transform 1 0 1752 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_89
timestamp 1710899220
transform 1 0 1808 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_90
timestamp 1710899220
transform 1 0 1760 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_91
timestamp 1710899220
transform 1 0 1360 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_92
timestamp 1710899220
transform 1 0 1480 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_93
timestamp 1710899220
transform 1 0 1424 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_94
timestamp 1710899220
transform 1 0 1304 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_95
timestamp 1710899220
transform 1 0 1160 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_96
timestamp 1710899220
transform 1 0 888 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_97
timestamp 1710899220
transform 1 0 800 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_98
timestamp 1710899220
transform 1 0 648 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_99
timestamp 1710899220
transform 1 0 608 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_100
timestamp 1710899220
transform 1 0 824 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_101
timestamp 1710899220
transform 1 0 960 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_102
timestamp 1710899220
transform 1 0 1088 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_103
timestamp 1710899220
transform 1 0 536 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_104
timestamp 1710899220
transform 1 0 512 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_105
timestamp 1710899220
transform 1 0 600 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_106
timestamp 1710899220
transform 1 0 664 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_107
timestamp 1710899220
transform 1 0 1144 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_108
timestamp 1710899220
transform 1 0 1144 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_109
timestamp 1710899220
transform 1 0 1320 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_110
timestamp 1710899220
transform 1 0 1448 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_111
timestamp 1710899220
transform 1 0 1296 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_112
timestamp 1710899220
transform 1 0 808 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_113
timestamp 1710899220
transform 1 0 960 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_114
timestamp 1710899220
transform 1 0 976 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_115
timestamp 1710899220
transform 1 0 856 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_116
timestamp 1710899220
transform 1 0 872 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_117
timestamp 1710899220
transform 1 0 1104 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_118
timestamp 1710899220
transform 1 0 1072 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_119
timestamp 1710899220
transform 1 0 728 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_120
timestamp 1710899220
transform 1 0 736 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_121
timestamp 1710899220
transform 1 0 736 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_122
timestamp 1710899220
transform 1 0 728 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_123
timestamp 1710899220
transform 1 0 880 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_124
timestamp 1710899220
transform 1 0 824 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_125
timestamp 1710899220
transform 1 0 680 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_126
timestamp 1710899220
transform 1 0 728 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_127
timestamp 1710899220
transform 1 0 696 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_128
timestamp 1710899220
transform 1 0 608 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_129
timestamp 1710899220
transform 1 0 728 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_130
timestamp 1710899220
transform 1 0 592 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_131
timestamp 1710899220
transform 1 0 208 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_132
timestamp 1710899220
transform 1 0 176 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_133
timestamp 1710899220
transform 1 0 368 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_134
timestamp 1710899220
transform 1 0 584 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_135
timestamp 1710899220
transform 1 0 336 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_136
timestamp 1710899220
transform 1 0 496 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_137
timestamp 1710899220
transform 1 0 296 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_138
timestamp 1710899220
transform 1 0 496 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_139
timestamp 1710899220
transform 1 0 144 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_140
timestamp 1710899220
transform 1 0 184 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_141
timestamp 1710899220
transform 1 0 280 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_142
timestamp 1710899220
transform 1 0 280 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_143
timestamp 1710899220
transform 1 0 232 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_144
timestamp 1710899220
transform 1 0 280 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_145
timestamp 1710899220
transform 1 0 208 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_146
timestamp 1710899220
transform 1 0 272 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_147
timestamp 1710899220
transform 1 0 168 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_148
timestamp 1710899220
transform 1 0 200 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_149
timestamp 1710899220
transform 1 0 280 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_150
timestamp 1710899220
transform 1 0 504 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_151
timestamp 1710899220
transform 1 0 312 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_152
timestamp 1710899220
transform 1 0 496 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_153
timestamp 1710899220
transform 1 0 280 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_154
timestamp 1710899220
transform 1 0 232 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_155
timestamp 1710899220
transform 1 0 2528 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_156
timestamp 1710899220
transform 1 0 2536 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_157
timestamp 1710899220
transform 1 0 2208 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_158
timestamp 1710899220
transform 1 0 2272 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_159
timestamp 1710899220
transform 1 0 2304 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_160
timestamp 1710899220
transform 1 0 2336 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_161
timestamp 1710899220
transform 1 0 2464 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_162
timestamp 1710899220
transform 1 0 2552 0 1 970
box -8 -3 34 105
use OAI22X1  OAI22X1_0
timestamp 1710899220
transform 1 0 1784 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_1
timestamp 1710899220
transform 1 0 1880 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_2
timestamp 1710899220
transform 1 0 1744 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_3
timestamp 1710899220
transform 1 0 1880 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_4
timestamp 1710899220
transform 1 0 680 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_5
timestamp 1710899220
transform 1 0 336 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_6
timestamp 1710899220
transform 1 0 304 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_7
timestamp 1710899220
transform 1 0 272 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_8
timestamp 1710899220
transform 1 0 1120 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_9
timestamp 1710899220
transform 1 0 992 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_10
timestamp 1710899220
transform 1 0 776 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_11
timestamp 1710899220
transform 1 0 504 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_12
timestamp 1710899220
transform 1 0 296 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_13
timestamp 1710899220
transform 1 0 344 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_14
timestamp 1710899220
transform 1 0 968 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_15
timestamp 1710899220
transform 1 0 1088 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_16
timestamp 1710899220
transform 1 0 1144 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_17
timestamp 1710899220
transform 1 0 1656 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_18
timestamp 1710899220
transform 1 0 1576 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_19
timestamp 1710899220
transform 1 0 1656 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_20
timestamp 1710899220
transform 1 0 1984 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_21
timestamp 1710899220
transform 1 0 1976 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_22
timestamp 1710899220
transform 1 0 1952 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_23
timestamp 1710899220
transform 1 0 1624 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_24
timestamp 1710899220
transform 1 0 1808 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_25
timestamp 1710899220
transform 1 0 1848 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_26
timestamp 1710899220
transform 1 0 1952 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_27
timestamp 1710899220
transform 1 0 1960 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_28
timestamp 1710899220
transform 1 0 2000 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_29
timestamp 1710899220
transform 1 0 1256 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_30
timestamp 1710899220
transform 1 0 1256 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_31
timestamp 1710899220
transform 1 0 1688 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_32
timestamp 1710899220
transform 1 0 1256 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_33
timestamp 1710899220
transform 1 0 1352 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_34
timestamp 1710899220
transform 1 0 1056 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_35
timestamp 1710899220
transform 1 0 936 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_36
timestamp 1710899220
transform 1 0 1136 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_37
timestamp 1710899220
transform 1 0 1096 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_38
timestamp 1710899220
transform 1 0 768 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_39
timestamp 1710899220
transform 1 0 1032 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_40
timestamp 1710899220
transform 1 0 904 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_41
timestamp 1710899220
transform 1 0 632 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_42
timestamp 1710899220
transform 1 0 512 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_43
timestamp 1710899220
transform 1 0 680 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_44
timestamp 1710899220
transform 1 0 632 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_45
timestamp 1710899220
transform 1 0 656 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_46
timestamp 1710899220
transform 1 0 568 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_47
timestamp 1710899220
transform 1 0 568 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_48
timestamp 1710899220
transform 1 0 512 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_49
timestamp 1710899220
transform 1 0 672 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_50
timestamp 1710899220
transform 1 0 632 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_51
timestamp 1710899220
transform 1 0 552 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_52
timestamp 1710899220
transform 1 0 504 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_53
timestamp 1710899220
transform 1 0 392 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_54
timestamp 1710899220
transform 1 0 448 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_55
timestamp 1710899220
transform 1 0 600 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_56
timestamp 1710899220
transform 1 0 616 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_57
timestamp 1710899220
transform 1 0 336 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_58
timestamp 1710899220
transform 1 0 408 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_59
timestamp 1710899220
transform 1 0 544 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_60
timestamp 1710899220
transform 1 0 528 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_61
timestamp 1710899220
transform 1 0 352 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_62
timestamp 1710899220
transform 1 0 408 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_63
timestamp 1710899220
transform 1 0 456 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_64
timestamp 1710899220
transform 1 0 472 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_65
timestamp 1710899220
transform 1 0 344 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_66
timestamp 1710899220
transform 1 0 448 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_67
timestamp 1710899220
transform 1 0 360 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_68
timestamp 1710899220
transform 1 0 448 0 1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_69
timestamp 1710899220
transform 1 0 328 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_70
timestamp 1710899220
transform 1 0 400 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_71
timestamp 1710899220
transform 1 0 392 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_72
timestamp 1710899220
transform 1 0 448 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_73
timestamp 1710899220
transform 1 0 312 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_74
timestamp 1710899220
transform 1 0 400 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_75
timestamp 1710899220
transform 1 0 352 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_76
timestamp 1710899220
transform 1 0 440 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_77
timestamp 1710899220
transform 1 0 384 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_78
timestamp 1710899220
transform 1 0 464 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_79
timestamp 1710899220
transform 1 0 624 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_80
timestamp 1710899220
transform 1 0 536 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_81
timestamp 1710899220
transform 1 0 344 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_82
timestamp 1710899220
transform 1 0 424 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_83
timestamp 1710899220
transform 1 0 584 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_84
timestamp 1710899220
transform 1 0 528 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_85
timestamp 1710899220
transform 1 0 320 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_86
timestamp 1710899220
transform 1 0 400 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_87
timestamp 1710899220
transform 1 0 360 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_88
timestamp 1710899220
transform 1 0 440 0 1 770
box -8 -3 46 105
use OR2X1  OR2X1_0
timestamp 1710899220
transform 1 0 1704 0 -1 2370
box -8 -3 40 105
use OR2X1  OR2X1_1
timestamp 1710899220
transform 1 0 1656 0 -1 2570
box -8 -3 40 105
use OR2X1  OR2X1_2
timestamp 1710899220
transform 1 0 1336 0 -1 2570
box -8 -3 40 105
use OR2X1  OR2X1_3
timestamp 1710899220
transform 1 0 856 0 -1 2570
box -8 -3 40 105
use OR2X1  OR2X1_4
timestamp 1710899220
transform 1 0 536 0 -1 2570
box -8 -3 40 105
use OR2X1  OR2X1_5
timestamp 1710899220
transform 1 0 232 0 -1 2570
box -8 -3 40 105
use OR2X1  OR2X1_6
timestamp 1710899220
transform 1 0 1040 0 1 570
box -8 -3 40 105
use OR2X1  OR2X1_7
timestamp 1710899220
transform 1 0 104 0 -1 1170
box -8 -3 40 105
use OR2X1  OR2X1_8
timestamp 1710899220
transform 1 0 128 0 -1 1370
box -8 -3 40 105
use OR2X1  OR2X1_9
timestamp 1710899220
transform 1 0 312 0 -1 1370
box -8 -3 40 105
use OR2X1  OR2X1_10
timestamp 1710899220
transform 1 0 128 0 -1 970
box -8 -3 40 105
use OR2X1  OR2X1_11
timestamp 1710899220
transform 1 0 2120 0 -1 1370
box -8 -3 40 105
use OR2X1  OR2X1_12
timestamp 1710899220
transform 1 0 1360 0 1 1770
box -8 -3 40 105
use OR2X1  OR2X1_13
timestamp 1710899220
transform 1 0 2176 0 1 1170
box -8 -3 40 105
use OR2X1  OR2X1_14
timestamp 1710899220
transform 1 0 1496 0 1 970
box -8 -3 40 105
use OR2X1  OR2X1_15
timestamp 1710899220
transform 1 0 2280 0 1 170
box -8 -3 40 105
use OR2X1  OR2X1_16
timestamp 1710899220
transform 1 0 2288 0 -1 970
box -8 -3 40 105
use top_module_VIA0  top_module_VIA0_0
timestamp 1710899220
transform 1 0 2720 0 1 2617
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_1
timestamp 1710899220
transform 1 0 2720 0 1 23
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_2
timestamp 1710899220
transform 1 0 24 0 1 2617
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_3
timestamp 1710899220
transform 1 0 24 0 1 23
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_4
timestamp 1710899220
transform 1 0 2696 0 1 2593
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_5
timestamp 1710899220
transform 1 0 2696 0 1 47
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_6
timestamp 1710899220
transform 1 0 48 0 1 2593
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_7
timestamp 1710899220
transform 1 0 48 0 1 47
box -10 -10 10 10
use top_module_VIA1  top_module_VIA1_0
timestamp 1710899220
transform 1 0 2720 0 1 2470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_1
timestamp 1710899220
transform 1 0 2720 0 1 2270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_2
timestamp 1710899220
transform 1 0 2720 0 1 2070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_3
timestamp 1710899220
transform 1 0 2720 0 1 1870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_4
timestamp 1710899220
transform 1 0 2720 0 1 1670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_5
timestamp 1710899220
transform 1 0 2720 0 1 1470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_6
timestamp 1710899220
transform 1 0 2720 0 1 1270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_7
timestamp 1710899220
transform 1 0 2720 0 1 1070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_8
timestamp 1710899220
transform 1 0 2720 0 1 870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_9
timestamp 1710899220
transform 1 0 2720 0 1 670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_10
timestamp 1710899220
transform 1 0 2720 0 1 470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_11
timestamp 1710899220
transform 1 0 2720 0 1 270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_12
timestamp 1710899220
transform 1 0 2720 0 1 70
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_13
timestamp 1710899220
transform 1 0 24 0 1 2470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_14
timestamp 1710899220
transform 1 0 24 0 1 2270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_15
timestamp 1710899220
transform 1 0 24 0 1 2070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_16
timestamp 1710899220
transform 1 0 24 0 1 1870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_17
timestamp 1710899220
transform 1 0 24 0 1 1670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_18
timestamp 1710899220
transform 1 0 24 0 1 1470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_19
timestamp 1710899220
transform 1 0 24 0 1 1270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_20
timestamp 1710899220
transform 1 0 24 0 1 1070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_21
timestamp 1710899220
transform 1 0 24 0 1 870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_22
timestamp 1710899220
transform 1 0 24 0 1 670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_23
timestamp 1710899220
transform 1 0 24 0 1 470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_24
timestamp 1710899220
transform 1 0 24 0 1 270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_25
timestamp 1710899220
transform 1 0 24 0 1 70
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_26
timestamp 1710899220
transform 1 0 48 0 1 170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_27
timestamp 1710899220
transform 1 0 48 0 1 370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_28
timestamp 1710899220
transform 1 0 48 0 1 570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_29
timestamp 1710899220
transform 1 0 48 0 1 770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_30
timestamp 1710899220
transform 1 0 48 0 1 970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_31
timestamp 1710899220
transform 1 0 48 0 1 1170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_32
timestamp 1710899220
transform 1 0 48 0 1 1370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_33
timestamp 1710899220
transform 1 0 48 0 1 1570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_34
timestamp 1710899220
transform 1 0 48 0 1 1770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_35
timestamp 1710899220
transform 1 0 48 0 1 1970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_36
timestamp 1710899220
transform 1 0 48 0 1 2170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_37
timestamp 1710899220
transform 1 0 48 0 1 2370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_38
timestamp 1710899220
transform 1 0 48 0 1 2570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_39
timestamp 1710899220
transform 1 0 2696 0 1 170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_40
timestamp 1710899220
transform 1 0 2696 0 1 370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_41
timestamp 1710899220
transform 1 0 2696 0 1 570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_42
timestamp 1710899220
transform 1 0 2696 0 1 770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_43
timestamp 1710899220
transform 1 0 2696 0 1 970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_44
timestamp 1710899220
transform 1 0 2696 0 1 1170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_45
timestamp 1710899220
transform 1 0 2696 0 1 1370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_46
timestamp 1710899220
transform 1 0 2696 0 1 1570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_47
timestamp 1710899220
transform 1 0 2696 0 1 1770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_48
timestamp 1710899220
transform 1 0 2696 0 1 1970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_49
timestamp 1710899220
transform 1 0 2696 0 1 2170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_50
timestamp 1710899220
transform 1 0 2696 0 1 2370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_51
timestamp 1710899220
transform 1 0 2696 0 1 2570
box -10 -3 10 3
use XNOR2X1  XNOR2X1_0
timestamp 1710899220
transform 1 0 1464 0 -1 2170
box -8 -3 64 105
use XNOR2X1  XNOR2X1_1
timestamp 1710899220
transform 1 0 1672 0 -1 2170
box -8 -3 64 105
use XNOR2X1  XNOR2X1_2
timestamp 1710899220
transform 1 0 1368 0 1 2170
box -8 -3 64 105
use XNOR2X1  XNOR2X1_3
timestamp 1710899220
transform 1 0 1488 0 -1 2370
box -8 -3 64 105
use XNOR2X1  XNOR2X1_4
timestamp 1710899220
transform 1 0 1280 0 -1 2370
box -8 -3 64 105
use XNOR2X1  XNOR2X1_5
timestamp 1710899220
transform 1 0 1368 0 1 2370
box -8 -3 64 105
use XNOR2X1  XNOR2X1_6
timestamp 1710899220
transform 1 0 1088 0 1 2370
box -8 -3 64 105
use XNOR2X1  XNOR2X1_7
timestamp 1710899220
transform 1 0 1168 0 -1 2570
box -8 -3 64 105
use XNOR2X1  XNOR2X1_8
timestamp 1710899220
transform 1 0 912 0 -1 2370
box -8 -3 64 105
use XNOR2X1  XNOR2X1_9
timestamp 1710899220
transform 1 0 704 0 1 2370
box -8 -3 64 105
use XNOR2X1  XNOR2X1_10
timestamp 1710899220
transform 1 0 584 0 -1 2370
box -8 -3 64 105
use XNOR2X1  XNOR2X1_11
timestamp 1710899220
transform 1 0 432 0 1 2370
box -8 -3 64 105
use XNOR2X1  XNOR2X1_12
timestamp 1710899220
transform 1 0 312 0 -1 2370
box -8 -3 64 105
use XNOR2X1  XNOR2X1_13
timestamp 1710899220
transform 1 0 144 0 -1 2370
box -8 -3 64 105
use XNOR2X1  XNOR2X1_14
timestamp 1710899220
transform 1 0 72 0 -1 2570
box -8 -3 64 105
use XNOR2X1  XNOR2X1_15
timestamp 1710899220
transform 1 0 656 0 -1 1370
box -8 -3 64 105
use XNOR2X1  XNOR2X1_16
timestamp 1710899220
transform 1 0 136 0 -1 1170
box -8 -3 64 105
use XNOR2X1  XNOR2X1_17
timestamp 1710899220
transform 1 0 160 0 -1 1370
box -8 -3 64 105
use XNOR2X1  XNOR2X1_18
timestamp 1710899220
transform 1 0 344 0 -1 1370
box -8 -3 64 105
use XNOR2X1  XNOR2X1_19
timestamp 1710899220
transform 1 0 72 0 -1 970
box -8 -3 64 105
use XNOR2X1  XNOR2X1_20
timestamp 1710899220
transform 1 0 1624 0 -1 1170
box -8 -3 64 105
use XNOR2X1  XNOR2X1_21
timestamp 1710899220
transform 1 0 752 0 -1 1370
box -8 -3 64 105
use XNOR2X1  XNOR2X1_22
timestamp 1710899220
transform 1 0 2000 0 1 1570
box -8 -3 64 105
use XNOR2X1  XNOR2X1_23
timestamp 1710899220
transform 1 0 2080 0 1 1570
box -8 -3 64 105
use XNOR2X1  XNOR2X1_24
timestamp 1710899220
transform 1 0 2176 0 -1 1370
box -8 -3 64 105
use XNOR2X1  XNOR2X1_25
timestamp 1710899220
transform 1 0 1464 0 -1 1170
box -8 -3 64 105
use XNOR2X1  XNOR2X1_26
timestamp 1710899220
transform 1 0 1728 0 -1 1370
box -8 -3 64 105
use XNOR2X1  XNOR2X1_27
timestamp 1710899220
transform 1 0 1456 0 1 1170
box -8 -3 64 105
use XNOR2X1  XNOR2X1_28
timestamp 1710899220
transform 1 0 1480 0 -1 1370
box -8 -3 64 105
use XNOR2X1  XNOR2X1_29
timestamp 1710899220
transform 1 0 1592 0 1 1170
box -8 -3 64 105
use XNOR2X1  XNOR2X1_30
timestamp 1710899220
transform 1 0 2584 0 -1 370
box -8 -3 64 105
use XOR2X1  XOR2X1_0
timestamp 1710899220
transform 1 0 72 0 1 2370
box -8 -3 64 105
use XOR2X1  XOR2X1_1
timestamp 1710899220
transform 1 0 2064 0 -1 1570
box -8 -3 64 105
use XOR2X1  XOR2X1_2
timestamp 1710899220
transform 1 0 2616 0 1 1170
box -8 -3 64 105
use XOR2X1  XOR2X1_3
timestamp 1710899220
transform 1 0 248 0 -1 1370
box -8 -3 64 105
use XOR2X1  XOR2X1_4
timestamp 1710899220
transform 1 0 136 0 1 770
box -8 -3 64 105
use XOR2X1  XOR2X1_5
timestamp 1710899220
transform 1 0 72 0 1 2170
box -8 -3 64 105
use XOR2X1  XOR2X1_6
timestamp 1710899220
transform 1 0 200 0 1 2170
box -8 -3 64 105
use XOR2X1  XOR2X1_7
timestamp 1710899220
transform 1 0 312 0 1 2170
box -8 -3 64 105
use XOR2X1  XOR2X1_8
timestamp 1710899220
transform 1 0 424 0 1 2170
box -8 -3 64 105
use XOR2X1  XOR2X1_9
timestamp 1710899220
transform 1 0 504 0 -1 2370
box -8 -3 64 105
use XOR2X1  XOR2X1_10
timestamp 1710899220
transform 1 0 1320 0 -1 2170
box -8 -3 64 105
use XOR2X1  XOR2X1_11
timestamp 1710899220
transform 1 0 72 0 -1 1370
box -8 -3 64 105
use XOR2X1  XOR2X1_12
timestamp 1710899220
transform 1 0 88 0 1 970
box -8 -3 64 105
use XOR2X1  XOR2X1_13
timestamp 1710899220
transform 1 0 88 0 1 1170
box -8 -3 64 105
use XOR2X1  XOR2X1_14
timestamp 1710899220
transform 1 0 2272 0 1 1570
box -8 -3 64 105
use XOR2X1  XOR2X1_15
timestamp 1710899220
transform 1 0 2176 0 1 1570
box -8 -3 64 105
use XOR2X1  XOR2X1_16
timestamp 1710899220
transform 1 0 1408 0 1 970
box -8 -3 64 105
use XOR2X1  XOR2X1_17
timestamp 1710899220
transform 1 0 1360 0 -1 1170
box -8 -3 64 105
use XOR2X1  XOR2X1_18
timestamp 1710899220
transform 1 0 1304 0 -1 1170
box -8 -3 64 105
use XOR2X1  XOR2X1_19
timestamp 1710899220
transform 1 0 1200 0 -1 1170
box -8 -3 64 105
use XOR2X1  XOR2X1_20
timestamp 1710899220
transform 1 0 1632 0 -1 1370
box -8 -3 64 105
use XOR2X1  XOR2X1_21
timestamp 1710899220
transform 1 0 1192 0 -1 1370
box -8 -3 64 105
use XOR2X1  XOR2X1_22
timestamp 1710899220
transform 1 0 1112 0 -1 1370
box -8 -3 64 105
use XOR2X1  XOR2X1_23
timestamp 1710899220
transform 1 0 1520 0 1 1170
box -8 -3 64 105
use XOR2X1  XOR2X1_24
timestamp 1710899220
transform 1 0 1560 0 -1 1370
box -8 -3 64 105
use XOR2X1  XOR2X1_25
timestamp 1710899220
transform 1 0 1408 0 -1 1370
box -8 -3 64 105
use XOR2X1  XOR2X1_26
timestamp 1710899220
transform 1 0 1296 0 -1 1370
box -8 -3 64 105
use XOR2X1  XOR2X1_27
timestamp 1710899220
transform 1 0 1360 0 1 1170
box -8 -3 64 105
use XOR2X1  XOR2X1_28
timestamp 1710899220
transform 1 0 1296 0 1 1170
box -8 -3 64 105
use XOR2X1  XOR2X1_29
timestamp 1710899220
transform 1 0 1176 0 1 1170
box -8 -3 64 105
<< labels >>
rlabel metal1 2012 1325 2012 1325 4 in_clka
rlabel electrodecontact s 2268 995 2268 995 4 in_clkb
rlabel electrodecontact s 2308 1015 2308 1015 4 in_restart
rlabel electrodecontact s 260 2005 260 2005 4 in_mult[4]
rlabel electrodecontact s 276 2005 276 2005 4 in_mult[3]
rlabel electrodecontact s 932 2005 932 2005 4 in_mult[2]
rlabel electrodecontact s 1188 2005 1188 2005 4 in_mult[1]
rlabel electrodecontact s 1236 2135 1236 2135 4 in_mult[0]
rlabel electrodecontact s 796 2325 796 2325 4 in_incr[4]
rlabel electrodecontact s 1004 2325 1004 2325 4 in_incr[3]
rlabel electrodecontact s 1156 2325 1156 2325 4 in_incr[2]
rlabel electrodecontact s 1244 2215 1244 2215 4 in_incr[1]
rlabel electrodecontact s 1324 2135 1324 2135 4 in_incr[0]
rlabel electrodecontact s 2228 1605 2228 1605 4 in_n_mines[4]
rlabel electrodecontact s 2228 1335 2228 1335 4 in_n_mines[3]
rlabel electrodecontact s 2324 1605 2324 1605 4 in_n_mines[2]
rlabel electrodecontact s 2132 1605 2132 1605 4 in_n_mines[1]
rlabel electrodecontact s 2052 1605 2052 1605 4 in_n_mines[0]
rlabel metal1 2500 935 2500 935 4 out_state_main[3]
rlabel electrodecontact s 2668 615 2668 615 4 out_state_main[2]
rlabel electrodecontact s 2628 735 2628 735 4 out_state_main[1]
rlabel electrodecontact s 2556 805 2556 805 4 out_state_main[0]
rlabel electrodecontact s 2556 1005 2556 1005 4 in_place
rlabel electrodecontact s 2460 815 2460 815 4 in_data_in
rlabel electrodecontact s 1332 935 1332 935 4 in_data[4]
rlabel electrodecontact s 1484 935 1484 935 4 in_data[3]
rlabel electrodecontact s 1356 1005 1356 1005 4 in_data[2]
rlabel electrodecontact s 1180 1005 1180 1005 4 in_data[1]
rlabel electrodecontact s 1180 935 1180 935 4 in_data[0]
rlabel electrodecontact s 2252 1005 2252 1005 4 out_start
rlabel electrodecontact s 2420 1125 2420 1125 4 out_place_done
rlabel electrodecontact s 764 1205 764 1205 4 out_mines[24]
rlabel metal1 564 735 564 735 4 out_mines[23]
rlabel electrodecontact s 676 1205 676 1205 4 out_mines[22]
rlabel metal1 468 735 468 735 4 out_mines[21]
rlabel electrodecontact s 972 805 972 805 4 out_mines[20]
rlabel electrodecontact s 828 735 828 735 4 out_mines[19]
rlabel electrodecontact s 812 735 812 735 4 out_mines[18]
rlabel electrodecontact s 532 335 532 335 4 out_mines[17]
rlabel metal1 780 1815 780 1815 4 out_mines[16]
rlabel electrodecontact s 452 205 452 205 4 out_mines[15]
rlabel metal1 948 405 948 405 4 out_mines[14]
rlabel electrodecontact s 972 335 972 335 4 out_mines[13]
rlabel electrodecontact s 988 805 988 805 4 out_mines[12]
rlabel electrodecontact s 1188 405 1188 405 4 out_mines[11]
rlabel electrodecontact s 1556 535 1556 535 4 out_mines[10]
rlabel electrodecontact s 844 805 844 805 4 out_mines[9]
rlabel electrodecontact s 1604 805 1604 805 4 out_mines[8]
rlabel electrodecontact s 1924 535 1924 535 4 out_mines[7]
rlabel electrodecontact s 1892 405 1892 405 4 out_mines[6]
rlabel electrodecontact s 1532 1005 1532 1005 4 out_mines[5]
rlabel electrodecontact s 1540 935 1540 935 4 out_mines[4]
rlabel electrodecontact s 1668 935 1668 935 4 out_mines[3]
rlabel electrodecontact s 1964 1615 1964 1615 4 out_mines[2]
rlabel electrodecontact s 1788 1005 1788 1005 4 out_mines[1]
rlabel electrodecontact s 1828 805 1828 805 4 out_mines[0]
rlabel electrodecontact s 2132 805 2132 805 4 out_load
rlabel electrodecontact s 716 805 716 805 4 out_temp_data_in[4]
rlabel electrodecontact s 716 1345 716 1345 4 out_temp_data_in[3]
rlabel metal1 1276 835 1276 835 4 out_temp_data_in[2]
rlabel metal1 524 1335 524 1335 4 out_temp_data_in[1]
rlabel electrodecontact s 516 1325 516 1325 4 out_temp_data_in[0]
rlabel electrodecontact s 2180 605 2180 605 4 out_decode
rlabel electrodecontact s 2164 605 2164 605 4 out_alu
rlabel metal1 2252 935 2252 935 4 out_alu_done
rlabel electrodecontact s 2148 1015 2148 1015 4 out_gameover
rlabel metal1 2044 1415 2044 1415 4 out_win
rlabel electrodecontact s 2668 1205 2668 1205 4 out_global_score[31]
rlabel electrodecontact s 2500 1205 2500 1205 4 out_global_score[30]
rlabel electrodecontact s 2380 1205 2380 1205 4 out_global_score[29]
rlabel electrodecontact s 2372 1335 2372 1335 4 out_global_score[28]
rlabel electrodecontact s 2348 1535 2348 1535 4 out_global_score[27]
rlabel electrodecontact s 2428 1535 2428 1535 4 out_global_score[26]
rlabel electrodecontact s 2548 1535 2548 1535 4 out_global_score[25]
rlabel electrodecontact s 2460 1735 2460 1735 4 out_global_score[24]
rlabel electrodecontact s 2380 1735 2380 1735 4 out_global_score[23]
rlabel electrodecontact s 2380 1805 2380 1805 4 out_global_score[22]
rlabel electrodecontact s 2460 1805 2460 1805 4 out_global_score[21]
rlabel electrodecontact s 2428 1935 2428 1935 4 out_global_score[20]
rlabel electrodecontact s 2444 2005 2444 2005 4 out_global_score[19]
rlabel electrodecontact s 2444 2205 2444 2205 4 out_global_score[18]
rlabel metal1 2364 2205 2364 2205 4 out_global_score[17]
rlabel electrodecontact s 2444 2335 2444 2335 4 out_global_score[16]
rlabel electrodecontact s 2484 2405 2484 2405 4 out_global_score[15]
rlabel electrodecontact s 2404 2405 2404 2405 4 out_global_score[14]
rlabel electrodecontact s 2204 2405 2204 2405 4 out_global_score[13]
rlabel electrodecontact s 2156 2335 2156 2335 4 out_global_score[12]
rlabel metal1 2068 2335 2068 2335 4 out_global_score[11]
rlabel electrodecontact s 2068 2535 2068 2535 4 out_global_score[10]
rlabel electrodecontact s 1988 2535 1988 2535 4 out_global_score[9]
rlabel electrodecontact s 1972 2405 1972 2405 4 out_global_score[8]
rlabel electrodecontact s 1972 2205 1972 2205 4 out_global_score[7]
rlabel electrodecontact s 1940 2135 1940 2135 4 out_global_score[6]
rlabel electrodecontact s 1972 2005 1972 2005 4 out_global_score[5]
rlabel metal1 2084 2005 2084 2005 4 out_global_score[4]
rlabel electrodecontact s 2172 2005 2172 2005 4 out_global_score[3]
rlabel electrodecontact s 2180 2135 2180 2135 4 out_global_score[2]
rlabel electrodecontact s 2276 2135 2276 2135 4 out_global_score[1]
rlabel electrodecontact s 2308 2205 2308 2205 4 out_global_score[0]
rlabel electrodecontact s 1924 1215 1924 1215 4 out_n_nearby[1]
rlabel electrodecontact s 1972 1125 1972 1125 4 out_n_nearby[0]
rlabel metal1 724 535 724 535 4 out_temp_decoded[24]
rlabel electrodecontact s 588 405 588 405 4 out_temp_decoded[23]
rlabel metal1 420 535 420 535 4 out_temp_decoded[22]
rlabel metal1 476 605 476 605 4 out_temp_decoded[21]
rlabel electrodecontact s 1140 535 1140 535 4 out_temp_decoded[20]
rlabel metal1 948 535 948 535 4 out_temp_decoded[19]
rlabel metal1 836 535 836 535 4 out_temp_decoded[18]
rlabel electrodecontact s 596 205 596 205 4 out_temp_decoded[17]
rlabel electrodecontact s 684 205 684 205 4 out_temp_decoded[16]
rlabel electrodecontact s 780 205 780 205 4 out_temp_decoded[15]
rlabel electrodecontact s 924 205 924 205 4 out_temp_decoded[14]
rlabel electrodecontact s 1132 205 1132 205 4 out_temp_decoded[13]
rlabel metal1 1228 205 1228 205 4 out_temp_decoded[12]
rlabel metal1 1556 205 1556 205 4 out_temp_decoded[11]
rlabel metal1 1612 335 1612 335 4 out_temp_decoded[10]
rlabel electrodecontact s 1396 205 1396 205 4 out_temp_decoded[9]
rlabel metal1 1796 205 1796 205 4 out_temp_decoded[8]
rlabel electrodecontact s 1940 335 1940 335 4 out_temp_decoded[7]
rlabel electrodecontact s 1836 405 1836 405 4 out_temp_decoded[6]
rlabel electrodecontact s 1548 805 1548 805 4 out_temp_decoded[5]
rlabel electrodecontact s 1452 805 1452 805 4 out_temp_decoded[4]
rlabel electrodecontact s 1620 805 1620 805 4 out_temp_decoded[3]
rlabel electrodecontact s 1820 605 1820 605 4 out_temp_decoded[2]
rlabel electrodecontact s 1948 735 1948 735 4 out_temp_decoded[1]
rlabel metal1 1556 605 1556 605 4 out_temp_decoded[0]
rlabel electrodecontact s 692 735 692 735 4 out_temp_cleared[24]
rlabel electrodecontact s 380 405 380 405 4 out_temp_cleared[23]
rlabel electrodecontact s 348 535 348 535 4 out_temp_cleared[22]
rlabel metal1 316 605 316 605 4 out_temp_cleared[21]
rlabel electrodecontact s 1124 535 1124 535 4 out_temp_cleared[20]
rlabel electrodecontact s 1012 735 1012 735 4 out_temp_cleared[19]
rlabel electrodecontact s 844 735 844 735 4 out_temp_cleared[18]
rlabel electrodecontact s 492 205 492 205 4 out_temp_cleared[17]
rlabel electrodecontact s 340 335 340 335 4 out_temp_cleared[16]
rlabel metal1 332 205 332 205 4 out_temp_cleared[15]
rlabel electrodecontact s 1012 205 1012 205 4 out_temp_cleared[14]
rlabel metal1 1076 205 1076 205 4 out_temp_cleared[13]
rlabel electrodecontact s 1188 205 1188 205 4 out_temp_cleared[12]
rlabel electrodecontact s 1700 335 1700 335 4 out_temp_cleared[11]
rlabel electrodecontact s 1620 205 1620 205 4 out_temp_cleared[10]
rlabel electrodecontact s 1700 205 1700 205 4 out_temp_cleared[9]
rlabel electrodecontact s 2028 535 2028 535 4 out_temp_cleared[8]
rlabel electrodecontact s 2020 335 2020 335 4 out_temp_cleared[7]
rlabel electrodecontact s 1996 205 1996 205 4 out_temp_cleared[6]
rlabel electrodecontact s 1556 935 1556 935 4 out_temp_cleared[5]
rlabel metal1 1764 1005 1764 1005 4 out_temp_cleared[4]
rlabel electrodecontact s 1892 935 1892 935 4 out_temp_cleared[3]
rlabel electrodecontact s 1996 605 1996 605 4 out_temp_cleared[2]
rlabel electrodecontact s 2004 805 2004 805 4 out_temp_cleared[1]
rlabel electrodecontact s 2044 935 2044 935 4 out_temp_cleared[0]
rlabel metal1 2284 525 2284 525 4 out_display
rlabel electrodecontact s 2332 725 2332 725 4 out_display_done
rlabel electrodecontact s 1140 1935 1140 1935 4 out_temp_index[4]
rlabel electrodecontact s 1012 2005 1012 2005 4 out_temp_index[3]
rlabel electrodecontact s 1156 1935 1156 1935 4 out_temp_index[2]
rlabel electrodecontact s 1508 2005 1508 2005 4 out_temp_index[1]
rlabel electrodecontact s 1380 2005 1380 2005 4 out_temp_index[0]
rlabel electrodecontact s 2116 1535 2116 1535 4 out_temp_mine_cnt[4]
rlabel electrodecontact s 2124 1535 2124 1535 4 out_temp_mine_cnt[3]
rlabel electrodecontact s 2116 1735 2116 1735 4 out_temp_mine_cnt[2]
rlabel electrodecontact s 2036 1735 2036 1735 4 out_temp_mine_cnt[1]
rlabel electrodecontact s 2020 1735 2020 1735 4 out_temp_mine_cnt[0]
rlabel metal2 38 37 38 37 4 gnd
rlabel metal2 14 13 14 13 4 vdd
<< properties >>
string path 20700.000 18945.000 20700.000 19035.000 
<< end >>
